netcdf CGMR_SRA1B_1_uas-change_2070-2099 {
dimensions:
	time = 12 ;
	latitude = 48 ;
	longitude = 96 ;
	bounds = 2 ;
Data:
 eastward_wind_anomaly =
  -0.02101934, -0.009349227, 0.0007255077, 0.008635581, 0.01405549, 
    0.01796177, 0.0207938, 0.02352816, 0.02598587, 0.02805299, 0.03010368, 
    0.03236604, 0.03438413, 0.03742802, 0.03863251, 0.03902304, 0.03920221, 
    0.0378511, 0.03591466, 0.03534484, 0.03184557, 0.02968097, 0.02543187, 
    0.0195725, 0.01262236, 0.00676322, 0.001245737, -0.001635313, 
    -0.002921104, -0.002285242, 0.00123024, 0.007659435, 0.01763654, 
    0.03116179, 0.04934204, 0.07137978, 0.09693307, 0.125937, 0.1578869, 
    0.1920177, 0.2267183, 0.2617931, 0.2966563, 0.3300548, 0.3644463, 
    0.398512, 0.4331801, 0.4495702, 0.471787, 0.4708431, 0.509531, 0.506048, 
    0.4611752, 0.5615656, 0.5717056, 0.5818455, 0.6013281, 0.6095312, 
    0.5980728, 0.576263, 0.554925, 0.556162, 0.5415624, 0.5121027, 0.4771416, 
    0.4400972, 0.4066826, 0.369736, 0.3347751, 0.2993746, 0.259596, 
    0.2219007, 0.1830498, 0.1551524, 0.09161103, 0.06317675, 0.0355401, 
    0.02769494, -0.01817083, -0.04922557, -0.07302094, -0.09299159, 
    -0.1075749, -0.1210353, -0.1297917, -0.1337795, -0.1329005, -0.1280665, 
    -0.1212795, -0.1106837, -0.09863949, -0.08522797, -0.07217455, 
    -0.05905628, -0.04603553, -0.03351927,
  -0.06901741, -0.05549202, -0.04180387, -0.03042692, -0.02544641, 
    -0.02655321, -0.03317755, -0.04535204, -0.06159556, -0.07918996, 
    -0.09466845, -0.1064686, -0.1164132, -0.1252837, -0.130492, -0.1311268, 
    -0.1327218, -0.1324614, -0.131908, -0.1307199, -0.1300037, -0.1272368, 
    -0.1223377, -0.1197987, -0.1161366, -0.1107816, -0.1107165, -0.1163156, 
    -0.1211979, -0.1320379, -0.1443262, -0.1533921, -0.1540756, -0.1449773, 
    -0.1275294, -0.1061265, -0.08223343, -0.05707061, -0.03083384, 
    -0.005443156, 0.01941033, 0.04411735, 0.05572221, 0.09069926, 0.1144136, 
    0.09696567, 0.1694756, 0.1896091, 0.1992933, 0.1904228, 0.2272391, 
    0.2746353, 0.2425224, 0.3003514, 0.2048272, 0.3798926, 0.3890233, 
    0.3774347, 0.3785416, 0.3744234, 0.3812432, 0.3872161, 0.3804293, 
    0.3791434, 0.393336, 0.434368, 0.4614676, 0.4782157, 0.508359, 0.5216565, 
    0.5252535, 0.495452, 0.4490652, 0.4108492, 0.3395926, 0.2916922, 
    0.2330334, 0.1845145, 0.119687, 0.08404249, 0.06096303, 0.0382905, 
    -0.01333708, -0.01302797, -0.05760789, -0.07948297, -0.1043364, 
    -0.1137928, -0.11905, -0.12058, -0.1202382, -0.1161691, -0.1110095, 
    -0.1044991, -0.09585661, -0.08290088,
  -0.04307342, 0.02188429, 0.08609326, 0.1319266, 0.1617444, 0.178818, 
    0.1774018, 0.1478771, 0.1048758, 0.05432236, 0.007268369, -0.03530985, 
    -0.0781157, -0.1210031, -0.1722075, -0.2280994, -0.2828195, -0.3384672, 
    -0.3928456, -0.4305734, -0.4353423, -0.4164621, -0.3752673, -0.3177153, 
    -0.2585031, -0.2078032, -0.1778716, -0.1670317, -0.1721098, -0.1948963, 
    -0.2316475, -0.2767159, -0.324388, -0.3652248, -0.3980865, -0.4133861, 
    -0.4171946, -0.4167063, -0.4074614, -0.385505, -0.3503973, -0.2782784, 
    -0.1994697, -0.1252348, -0.0591867, -0.01522508, 0.009400554, 0.0205985, 
    0.02865511, 0.04864198, 0.05819613, 0.05342722, 0.05406207, 0.06610626, 
    0.0935477, 0.1115816, 0.1284598, 0.1317638, 0.1202893, 0.09078074, 
    0.0491792, 0.01395783, 0.001522958, 0.001327634, 0.0127697, 0.02813429, 
    0.05845656, 0.09553337, 0.1225516, 0.1396903, 0.1405855, 0.1442801, 
    0.1507417, 0.1495861, 0.1360444, 0.141562, 0.06524366, 0.08334264, 
    0.09177363, 0.0619396, 0.04384065, 0.03086865, 0.02108675, -0.00252974, 
    -0.0312407, -0.0786202, -0.1033273, -0.1399485, -0.1677316, -0.1746001, 
    -0.1860259, -0.1740141, -0.165339, -0.1554757, -0.1317617, -0.09300828,
  -0.3100166, -0.3438872, -0.3659248, -0.3592353, -0.3363347, -0.3051662, 
    -0.2554755, -0.1894438, -0.1324939, -0.08978558, -0.05117881, 
    0.0008066893, 0.03410757, 0.03776968, 0.04081333, 0.05145785, 0.05922152, 
    0.05552685, 0.0512951, 0.04322219, 0.01493454, -0.041641, -0.1144762, 
    -0.1849028, -0.2375558, -0.2682362, -0.2607818, -0.2292387, -0.2205637, 
    -0.2348052, -0.2714588, -0.3123767, -0.3509673, -0.3727771, -0.3729886, 
    -0.3876694, -0.4279363, -0.4971588, -0.5724518, -0.6289296, -0.6453359, 
    -0.5928943, -0.4471099, -0.2483301, -0.1244534, -0.1021553, -0.09611702, 
    -0.1009673, -0.08055711, -0.07632535, -0.09823291, -0.1023507, 
    -0.06504604, -0.001488119, 0.04006463, 0.06224883, 0.1108329, 0.2017183, 
    0.2263439, 0.2288829, 0.1974703, 0.1694268, 0.1566175, 0.1933525, 
    0.2516532, 0.3253353, 0.3734636, 0.4112401, 0.4067316, 0.3836846, 
    0.3669205, 0.3466079, 0.3263931, 0.2878675, 0.288307, 0.28554, 0.2957287, 
    0.3006929, 0.2818452, 0.2543224, 0.2392508, 0.2057222, 0.1769624, 
    0.1433687, 0.1101167, 0.06543893, -0.01035857, -0.07564175, -0.1262928, 
    -0.1902413, -0.2039783, -0.209675, -0.2253488, -0.2332426, -0.2582753, 
    -0.2745512,
  -0.1849841, -0.2066637, -0.245189, -0.230948, -0.259073, -0.1875563, 
    -0.1249914, -0.06136823, 0.02450418, 0.1179123, 0.2218673, 0.3082447, 
    0.3510344, 0.3338301, 0.2635834, 0.2030367, 0.1676364, 0.1461519, 
    0.1436616, 0.1329846, 0.1110609, 0.02867079, -0.134871, -0.2913649, 
    -0.3835356, -0.4280181, -0.4336984, -0.4171293, -0.3792386, -0.3517158, 
    -0.3420316, -0.3380276, -0.3267322, -0.3056221, -0.2833076, -0.2816639, 
    -0.3123443, -0.3746164, -0.4490305, -0.5161041, -0.5378813, -0.5205636, 
    -0.4659901, -0.3724517, -0.3102609, -0.2972076, -0.3739653, -0.3511952, 
    -0.3413807, -0.3415272, -0.3191964, -0.3350168, -0.3383045, -0.3491932, 
    -0.3204008, -0.2640857, -0.1801503, -0.08003628, 0.06101173, 0.1592702, 
    0.2257416, 0.2761484, 0.3538991, 0.4445405, 0.5419365, 0.595322, 
    0.6489027, 0.7484798, 0.8920175, 0.9259369, 0.8104258, 0.6621842, 
    0.6092052, 0.499277, 0.4707936, 0.5127534, 0.5260346, 0.5706962, 
    0.5725842, 0.5731376, 0.4694916, 0.4948661, 0.4615164, 0.470631, 
    0.4803478, 0.4501232, 0.367864, 0.2492443, 0.1320405, 0.02247024, 
    -0.04543352, -0.1105701, -0.1385323, -0.1562569, -0.1627185, -0.1662341,
  -0.2273669, -0.145238, 0.03851855, 0.1273695, 0.126165, 0.1540294, 
    0.1419363, 0.05559206, 0.01405549, 0.002841473, -0.02785516, -0.04170609, 
    0.05666661, 0.2109303, 0.3376882, 0.3295343, 0.3209896, 0.2882417, 
    0.2958264, 0.2923433, 0.2991793, 0.2683039, 0.2411058, 0.09309149, 
    -0.06561565, -0.1326895, -0.1303945, -0.07744884, -0.01966858, 
    0.01005173, 0.02898073, 0.0655365, 0.1313081, 0.1681733, 0.2301519, 
    0.2725184, 0.3163013, 0.2993093, 0.3089938, 0.2890558, 0.3085058, 
    0.3186784, 0.3220801, 0.2378349, 0.1165619, -0.110733, -0.2798573, 
    -0.3371326, -0.5352933, -0.6382232, -0.631729, -0.6393461, -0.6690662, 
    -0.6912341, -0.6912504, -0.6927153, -0.6471099, -0.5376046, -0.3592681, 
    -0.1904367, -0.02505582, 0.09720981, 0.2316987, 0.3720796, 0.5451102, 
    0.7488211, 0.8775808, 1.000205, 1.095599, 1.032024, 0.9991302, 0.7239025, 
    0.6296479, 0.5807222, 0.5236908, 0.4745208, 0.4803639, 0.5247489, 
    0.5585542, 0.6256603, 0.5490978, 0.5263602, 0.5096934, 0.5015229, 
    0.52623, 0.4972423, 0.5101492, 0.5074148, 0.5089447, 0.5034435, 0.471982, 
    0.4207449, 0.3542737, 0.2527275, 0.09649384, -0.1056546,
  0.3508067, 0.3265231, 0.2574964, 0.2275977, 0.1473405, 0.03713536, 
    -0.0436914, -0.05466151, -0.04865575, -0.01608753, 0.01752257, 
    -0.005475283, 0.004810572, 0.1159592, 0.2183354, 0.3685145, 0.4116786, 
    0.4846766, 0.5493746, 0.5989511, 0.7181735, 0.8088958, 0.853704, 
    0.709075, 0.5106049, 0.3153417, 0.2348239, 0.1881933, 0.1499772, 
    0.1205499, 0.1561935, 0.1881764, 0.2091889, 0.1333745, 0.1640234, 
    0.2478769, 0.326246, 0.3433034, 0.6472585, 0.8518159, 0.875237, 
    0.8963146, 0.9627044, 0.9833913, 0.8694432, 0.6642345, 0.4295014, 
    0.1725353, -0.01579475, -0.1230538, -0.1793852, -0.2252512, -0.2301014, 
    -0.150186, -0.0548898, -0.03358448, -0.1205962, -0.2138742, -0.2010487, 
    -0.08848356, 0.1167085, 0.336077, 0.5260185, 0.7283622, 1.004616, 
    1.300302, 1.584108, 1.795143, 1.896005, 1.866204, 1.797324, 1.756943, 
    1.756422, 1.718922, 1.553232, 1.313762, 1.203102, 1.141578, 1.048919, 
    0.7761323, 0.6511649, 0.5375417, 0.4332124, 0.3698173, 0.2926524, 
    0.1705171, 0.07175404, 0.05105096, 0.06742465, 0.1751558, 0.3453218, 
    0.4992118, 0.5362723, 0.4994395, 0.4619396, 0.4213472,
  1.753948, 1.799391, 1.821478, 1.912168, 1.984205, 2.033505, 2.038242, 
    2.069915, 2.153525, 2.215699, 2.305494, 2.387314, 2.383277, 2.314332, 
    2.235637, 2.19996, 2.177988, 2.141301, 2.04773, 1.984677, 2.003818, 
    2.077271, 2.102223, 2.098072, 1.945778, 1.655804, 1.347258, 1.146787, 
    0.998382, 0.8384863, 0.6971126, 0.6046159, 0.6244559, 0.7319429, 
    0.7847748, 0.7636328, 0.8094174, 1.037493, 1.247942, 1.318727, 1.249961, 
    1.213795, 1.323675, 1.522552, 1.68012, 1.692945, 1.584921, 1.46277, 
    1.364234, 1.282268, 1.120745, 0.951816, 0.8039644, 0.7797456, 0.853232, 
    0.9540619, 0.9841565, 0.9425875, 0.9061943, 0.9901625, 1.145517, 
    1.335556, 1.440146, 1.458017, 1.518027, 1.670615, 1.904941, 2.136256, 
    2.291758, 2.39166, 2.431813, 2.478916, 2.483294, 2.386533, 2.244411, 
    2.074554, 1.947633, 1.962184, 1.999163, 1.947194, 1.851165, 1.818499, 
    1.842148, 1.871477, 1.705787, 1.427304, 1.183831, 0.9273205, 0.7203543, 
    0.6106212, 0.73956, 1.027076, 1.293776, 1.449635, 1.526588, 1.646917,
  2.233994, 2.315325, 2.408587, 2.558261, 2.748984, 2.97859, 3.189056, 
    3.272731, 3.230853, 3.211093, 3.300563, 3.408213, 3.451979, 3.462102, 
    3.454973, 3.436858, 3.368792, 3.254339, 3.132936, 3.079762, 3.045029, 
    3.013844, 2.973089, 2.989267, 2.956357, 2.788665, 2.543385, 2.384954, 
    2.340813, 2.277646, 2.169671, 2.075416, 2.061484, 2.093027, 2.07234, 
    1.971738, 1.821673, 1.73235, 1.778427, 1.898658, 2.08331, 2.304729, 
    2.60263, 2.913632, 3.16806, 3.225237, 3.177158, 3.052598, 2.911761, 
    2.812282, 2.631732, 2.354486, 2.029046, 1.713714, 1.570322, 1.600351, 
    1.662884, 1.735996, 1.806211, 1.843385, 1.919491, 2.040015, 2.193824, 
    2.296965, 2.272795, 2.191773, 2.147567, 2.200774, 2.202662, 2.12566, 
    2.076214, 2.088323, 2.112053, 2.155803, 2.260784, 2.37081, 2.281162, 
    2.113258, 2.123577, 2.193775, 2.153476, 2.090586, 2.24472, 2.506715, 
    2.670077, 2.660882, 2.617067, 2.494329, 2.21417, 1.920859, 1.78012, 
    1.827191, 1.931243, 1.956243, 2.019638, 2.154485,
  2.405755, 2.462672, 2.576344, 2.623658, 2.676848, 2.872389, 3.119117, 
    3.288437, 3.311224, 3.335019, 3.357203, 3.287916, 3.194394, 3.130966, 
    3.1212, 3.234237, 3.407561, 3.482691, 3.41067, 3.328248, 3.395175, 
    3.465227, 3.458424, 3.508537, 3.639088, 3.773219, 3.859709, 3.887151, 
    3.863144, 3.84, 3.775938, 3.633652, 3.390422, 3.127532, 2.91456, 
    2.740553, 2.574488, 2.456047, 2.460328, 2.542587, 2.608668, 2.674212, 
    2.899797, 3.329273, 3.794035, 4.035491, 4.032333, 3.952158, 3.917636, 
    3.863177, 3.71347, 3.46902, 3.122308, 2.716627, 2.380576, 2.180852, 
    2.033359, 1.931975, 1.924195, 1.950514, 1.924896, 1.897861, 1.969964, 
    2.070224, 2.092228, 2.027255, 2.068189, 2.223203, 2.264657, 2.161565, 
    2.086761, 2.107903, 2.010067, 1.928833, 1.989608, 1.976359, 1.751701, 
    1.57164, 1.638339, 1.897535, 2.145957, 2.15372, 2.237656, 2.627109, 
    3.060296, 3.310719, 3.453182, 3.472682, 3.283749, 2.9969, 2.678476, 
    2.401132, 2.263047, 2.271038, 2.358798, 2.39135,
  2.107186, 2.153865, 2.169181, 2.14633, 2.075008, 2.120028, 2.313029, 
    2.515682, 2.595809, 2.537199, 2.42867, 2.325154, 2.314478, 2.320727, 
    2.216414, 2.157641, 2.284985, 2.465096, 2.437687, 2.290894, 2.350903, 
    2.599341, 2.846281, 3.085261, 3.34335, 3.568807, 3.707771, 3.696898, 
    3.637963, 3.670988, 3.725562, 3.673625, 3.513859, 3.29449, 3.081453, 
    2.955445, 2.840031, 2.695354, 2.589152, 2.629485, 2.661402, 2.607707, 
    2.613013, 2.875578, 3.28925, 3.597649, 3.746053, 3.788713, 3.925205, 
    3.987265, 3.914918, 3.757399, 3.472112, 3.050466, 2.718955, 2.505185, 
    2.282171, 2.0643, 1.944818, 1.864804, 1.796673, 1.699065, 1.52081, 
    1.413062, 1.375367, 1.356275, 1.385653, 1.519263, 1.640535, 1.645712, 
    1.648999, 1.634888, 1.532251, 1.454988, 1.379988, 1.185133, 1.00512, 
    1.170826, 1.442831, 1.661093, 1.726555, 1.671249, 1.684546, 1.993401, 
    2.425611, 2.804631, 3.065308, 3.099407, 2.9726, 2.875529, 2.747535, 
    2.508585, 2.253622, 2.126262, 2.058586, 2.062687,
  0.972095, 1.011645, 1.004175, 0.9300375, 0.8538494, 0.7900476, 0.7703371, 
    0.8130779, 0.9117918, 0.946867, 0.8779702, 0.7960205, 0.7343993, 
    0.6728268, 0.5923424, 0.5578213, 0.5789795, 0.7433186, 0.9539633, 
    1.112784, 1.280982, 1.418204, 1.520499, 1.695028, 1.936989, 2.146966, 
    2.328183, 2.434465, 2.485898, 2.542897, 2.537558, 2.450626, 2.416317, 
    2.412313, 2.270451, 2.117407, 2.064119, 1.923983, 1.772062, 1.791707, 
    1.927465, 2.046248, 2.035392, 1.950627, 2.033716, 2.288305, 2.417977, 
    2.610279, 2.821541, 3.024211, 3.04524, 3.010556, 2.983163, 2.810833, 
    2.561695, 2.305071, 2.041595, 1.742099, 1.52439, 1.327467, 1.210638, 
    1.137232, 1.000057, 0.9015551, 0.8657475, 0.8557057, 0.820159, 0.8104258, 
    0.8264575, 0.8157964, 0.7692471, 0.7162685, 0.621314, 0.6329679, 
    0.7065034, 0.4748783, 0.238925, 0.3705816, 0.4836841, 0.4142666, 
    0.5504804, 0.7753992, 0.8135991, 0.8364673, 0.9815025, 1.201197, 
    1.454843, 1.635164, 1.728199, 1.803165, 1.805688, 1.712524, 1.51049, 
    1.276196, 1.090014, 0.9890051,
  -0.09216309, -0.1758709, -0.2540445, -0.303442, -0.3276129, -0.3466558, 
    -0.3935461, -0.5585527, -0.6792231, -0.6485758, -0.6352124, -0.6906815, 
    -0.7438226, -0.6886144, -0.5571194, -0.4311275, -0.3041916, -0.141902, 
    0.003881454, 0.1029053, 0.1677818, 0.1365805, 0.108798, 0.2120209, 
    0.3859787, 0.6104918, 0.8191013, 0.9894295, 1.037444, 1.024747, 1.127092, 
    1.149324, 1.03933, 0.9641199, 0.9160728, 0.893384, 0.8131447, 0.6196384, 
    0.630558, 0.587688, 0.2878661, 0.2287025, 0.4140706, 0.4650965, 
    0.5509686, 0.8157964, 1.069508, 1.084904, 1.227255, 1.552661, 1.720175, 
    1.651506, 1.632512, 1.608472, 1.550041, 1.386776, 1.108407, 0.8315196, 
    0.6201262, 0.404469, 0.2542734, 0.1627693, 0.1173759, 0.1073327, 
    0.03291893, -0.07337999, -0.1225009, -0.1774487, -0.1642485, -0.1957917, 
    -0.2291412, -0.08726311, -0.0125556, -0.1354074, -0.1472077, -0.1523027, 
    -0.120564, -0.1379795, -0.5290923, -0.8656976, -0.5675371, -0.2125239, 
    -0.224731, -0.2578201, -0.2126374, -0.1281161, -0.002155781, 0.1342373, 
    0.3640385, 0.5179124, 0.4910736, 0.4248462, 0.3232837, 0.1915126, 
    0.1333418, 0.04327011,
  -0.7123771, -0.8190336, -0.950983, -1.138012, -1.42906, -1.706224, 
    -1.811921, -1.883519, -2.078084, -2.109251, -1.873997, -1.649453, 
    -1.589753, -1.53264, -1.400805, -1.323103, -1.292374, -1.189541, 
    -1.13448, -1.14934, -1.146361, -1.125707, -1.043969, -1.011206, 
    -1.004874, -0.8901606, -0.8852453, -0.8657141, -0.7078848, -0.6972728, 
    -0.6909251, -0.672533, -0.6548738, -0.490356, -0.4283934, -0.4307203, 
    -0.498282, -0.7440014, -0.7835193, -0.9905181, -1.728995, -1.741088, 
    -1.324845, -1.203328, -1.044571, -0.7116609, -0.3225818, -0.1419511, 
    -0.2457108, -0.0350008, 0.276392, 0.4603281, 0.4769135, 0.3829193, 
    0.422307, 0.4374275, 0.3191824, 0.1687427, -0.04562902, -0.2850337, 
    -0.4512444, -0.5866451, -0.6298575, -0.5804601, -0.647696, -0.6970935, 
    -0.7133698, -0.8358469, -0.7864165, -0.579174, -0.5405836, -0.5427809, 
    -0.4817295, -0.4764881, -0.5494218, -0.5710361, -0.2895741, -0.1454341, 
    -0.5890857, -1.10375, -0.9083567, -0.9118559, -1.096084, -1.174601, 
    -1.240698, -1.177449, -0.9815669, -0.8561759, -0.7279215, -0.5516677, 
    -0.4718499, -0.4525623, -0.432478, -0.4800854, -0.533308, -0.5960684,
  -1.196801, -1.263288, -1.418757, -1.762702, -2.223428, -2.702823, 
    -3.073282, -3.046361, -2.638435, -2.469701, -2.419929, -2.317569, 
    -2.318822, -2.327628, -2.153881, -1.925772, -1.955558, -2.090877, 
    -2.122663, -2.103669, -2.156762, -2.201342, -2.138679, -2.142163, 
    -2.240388, -2.122046, -2.158927, -2.30852, -2.190665, -2.282006, 
    -2.506729, -2.460977, -2.163435, -1.580134, -1.414899, -1.561286, 
    -1.356648, -1.01944, -0.7217841, -1.050381, -1.745092, -1.748152, 
    -1.722273, -2.145564, -2.274909, -2.20821, -1.993578, -1.722827, 
    -1.562833, -1.315161, -1.056013, -0.8550038, -0.7479563, -0.7032297, 
    -0.5830636, -0.5182853, -0.4617584, -0.4937727, -0.6437082, -0.7613026, 
    -0.8945378, -0.9817452, -0.9851959, -0.9691966, -0.9868886, -1.015258, 
    -0.9527416, -0.9087148, -0.9162018, -0.8516185, -0.6384513, -0.5204172, 
    -0.5729725, -0.5290272, -0.4571682, -0.4261137, -0.08880901, 0.3227146, 
    -0.2111398, -0.5666082, -0.4284085, -0.6953031, -1.014883, -1.183617, 
    -1.183292, -1.017536, -0.8959218, -0.7761297, -0.8532617, -0.8824773, 
    -0.8114011, -0.8674717, -0.8880448, -0.9101143, -1.001635, -1.08404,
  -1.127725, -1.23448, -1.272387, -1.26319, -0.9375395, -0.6858957, 
    -0.9353096, -1.179939, -0.8270576, -1.036628, -1.725121, -2.257917, 
    -2.434528, -2.282233, -2.035635, -1.865062, -1.795922, -1.873152, 
    -2.009415, -2.212263, -2.326065, -2.492601, -2.659365, -2.676944, 
    -2.802904, -2.831436, -2.756631, -2.849177, -2.867976, -2.837018, 
    -2.437018, -1.980215, -1.644701, -1.182852, -0.8675524, -0.812214, 
    -0.8660551, -0.8618559, -0.7440662, -1.089249, -1.683991, -1.63723, 
    -1.903929, -2.540974, -2.872094, -3.065144, -3.074828, -2.921459, 
    -2.615176, -2.228653, -2.029645, -1.764867, -1.43404, -1.267032, 
    -1.147712, -1.075772, -0.9932524, -0.9465889, -0.9820219, -0.9248442, 
    -1.01472, -1.112751, -1.116462, -1.120043, -1.100332, -1.120255, 
    -1.089037, -0.9456125, -0.8447662, -0.9116281, -0.7930245, -0.5891346, 
    -0.4878813, -0.4435453, -0.3690825, -0.1216704, 0.1383229, 0.459873, 
    -0.01861051, -0.4712636, -0.1594632, -0.1298733, -0.2944238, -0.408975, 
    -0.5343819, -0.4486072, -0.691348, -0.8340402, -1.022712, -1.155866, 
    -1.035195, -1.039443, -1.006452, -0.9835678, -0.9820546, -0.9715403,
  -0.7260814, -0.6746166, -0.4973214, -0.021492, 0.3755467, 0.2990002, 
    0.02491158, -0.2197498, -0.2180897, -0.381485, -0.7196529, -1.151635, 
    -1.660262, -1.843432, -1.41529, -1.024747, -1.056078, -1.273835, 
    -1.480834, -1.664574, -1.765746, -1.877839, -2.120059, -2.181338, 
    -2.28308, -2.461742, -2.411466, -2.387589, -2.201602, -1.676716, 
    -1.112295, -1.066608, -1.143253, -0.9509189, -0.8685942, -0.663044, 
    -0.4172597, -0.5724028, -0.849893, -1.173102, -1.653897, -1.892976, 
    -2.387849, -2.902464, -3.169685, -3.181208, -3.021589, -2.833292, 
    -2.618024, -2.295482, -2.119701, -1.853099, -1.472192, -1.290779, 
    -1.113646, -1.072956, -1.148965, -1.141641, -1.171638, -1.081843, 
    -0.969799, -0.9608303, -1.070808, -1.188875, -1.233634, -1.19335, 
    -1.132787, -1.179646, -0.9710686, -0.8783109, -0.8880768, -0.7771881, 
    -0.4680741, -0.2836502, -0.2220454, 0.01024699, -0.1726144, 0.3754165, 
    0.1698985, -0.5585847, -0.125479, 0.1908298, 0.1183689, 0.03344035, 
    -0.3868394, -0.4276114, -0.2872138, -0.3933011, -0.5692779, -0.6815337, 
    -0.7186592, -0.7503977, -0.7523017, -0.7855375, -0.7822335, -0.7125558,
  -0.008291245, 0.2597423, 0.4117932, 0.7585547, 0.6773693, 0.001734734, 
    -0.3052967, -0.1787829, 0.04379153, 0.002109289, 0.1690514, 0.2040782, 
    -0.3790598, -1.024878, -1.029271, -0.6068268, -0.5734124, -0.7565341, 
    -0.9490476, -1.016772, -1.167455, -1.238273, -1.270011, -1.391186, 
    -1.42242, -1.45673, -1.40367, -1.284626, -0.894392, -0.07702541, 
    0.2901297, -0.2430571, -0.5638092, -0.4617915, -0.6310129, -0.561645, 
    -0.1905341, -0.2569567, -0.6478096, -1.032689, -1.534382, -1.756681, 
    -1.917374, -2.174861, -2.335229, -2.286905, -2.215763, -2.095581, 
    -1.903913, -1.608064, -1.25113, -1.213158, -1.144408, -1.001276, 
    -0.9237208, -0.8516183, -0.9567454, -1.011401, -1.137475, -1.308878, 
    -1.312329, -1.313305, -1.419359, -1.428311, -1.448119, -1.404353, 
    -1.200642, -1.191999, -1.02115, -0.9602447, -0.8002191, -0.6276608, 
    -0.442276, -0.1784415, -0.04914522, 0.1031022, -0.4794993, 0.1074641, 
    0.3480887, -0.7434146, -0.2515044, 0.1218843, 0.01410425, 0.111614, 
    -0.3588122, -0.6012442, -0.3253984, -0.3404367, -0.4633529, -0.4072175, 
    -0.4959869, -0.4363515, -0.4378815, -0.4179106, -0.3193274, -0.203474,
  0.4335055, 0.5490975, 0.3778744, 0.2195244, 0.04405236, 0.02727187, 
    0.03137338, -0.1761138, -0.1940668, -0.06880546, 0.1783452, 0.2031506, 
    -0.0381743, -0.349323, -0.7281322, -0.4167881, -0.1328855, -0.1620674, 
    -0.4553461, -0.5484776, -0.514185, -0.5218339, -0.5813718, -0.565063, 
    -0.4469967, -0.3812251, -0.2407465, -0.06141663, 0.09102416, 0.3404877, 
    0.6443941, 0.7358654, 0.6024507, 0.2497325, -0.1018794, -0.1058824, 
    0.02095664, 0.0207938, -0.3856189, -0.8549552, -1.211873, -1.203897, 
    -0.7982011, -0.792325, -1.00279, -1.162149, -1.300529, -1.158667, 
    -0.8580647, -0.8175044, -0.5316806, -0.4893146, -0.6019278, -0.5526767, 
    -0.6540275, -0.6452389, -0.6995034, -0.9272699, -1.164835, -1.423721, 
    -1.530053, -1.485164, -1.445532, -1.388859, -1.249633, -1.154923, 
    -1.040974, -0.9438882, -0.7532463, -0.6701736, -0.4888582, -0.3754306, 
    -0.3041086, -0.06052208, -0.09473372, 0.01491833, -0.07694387, 0.2718511, 
    0.306715, -0.4214424, -0.5093331, -0.2278877, -0.08815801, -0.08978564, 
    -0.1495675, -0.7041245, -0.4578364, -0.2702062, -0.3065176, -0.163744, 
    -0.1949782, -0.06047297, -0.03319454, 0.05227137, 0.1955328, 0.3491945,
  0.514641, 0.5337498, 0.2324637, -0.08573282, -0.4806381, -0.392634, 
    0.01587844, 0.01573205, -0.204385, -0.2647206, -0.0976305, -0.06633186, 
    -0.3672271, -0.6591052, -1.196898, -0.888582, -0.2030835, 0.2101321, 
    0.371624, 0.3200288, 0.3284917, 0.4457121, 0.3680425, 0.3350029, 
    0.3791752, 0.4261804, 0.4118581, 0.3634043, 0.4372818, 0.4617605, 
    0.3449963, 0.69568, 1.192685, 1.047308, 0.7559175, 0.3252697, 0.08716762, 
    0.2072847, -0.1216378, -0.1486893, 0.1439538, 0.4798751, 0.6341074, 
    0.5485771, 0.3249273, 0.1831145, 0.007219791, -0.1212478, 0.10953, 
    0.1486416, 0.07118416, 0.04665613, -0.1625881, -0.2915435, -0.4232821, 
    -0.6808996, -0.8133702, -0.9603758, -1.108211, -1.346101, -1.375236, 
    -1.26726, -1.088354, -0.933341, -0.821053, -0.670125, -0.5186758, 
    -0.4114656, -0.4304762, -0.3288813, -0.3241286, -0.2367587, -0.1154208, 
    -0.01652718, -0.006337881, 0.1717703, 0.4222423, 0.4452567, 0.2178316, 
    0.05957961, -0.3935454, -0.5177315, -0.2013579, -0.1551502, -0.1211333, 
    -0.5994208, -0.3518953, 0.03451443, -0.00288868, 0.1427169, 0.1563892, 
    0.2228928, 0.3347578, 0.4101648, 0.4064708, 0.4951429,
  0.2572851, 0.2007092, 0.07500929, 0.1536391, -0.10445, -0.2623118, 
    -0.06880581, 0.02997348, 0.06389278, -0.06115615, -0.2633858, -0.2787828, 
    -0.5208892, -0.9077055, -1.301992, -1.21267, -0.5184155, 0.2113531, 
    0.670191, 0.8317306, 0.8230553, 1.092994, 1.168645, 1.041203, 0.9410899, 
    0.9469817, 0.8414648, 0.7934663, 0.7673109, 0.8225353, 0.5340912, 
    0.06963754, 0.1517177, 0.5321538, 0.8323498, 0.5237558, 0.3911226, 
    0.6758558, 0.2878348, 0.2144296, 0.6253673, 1.046412, 1.227809, 1.250286, 
    0.8928641, 0.8947846, 0.9152762, 0.3396418, -0.1822982, -0.2773178, 
    -0.5081782, -0.5141354, -0.4900632, -0.7633371, -0.6729407, -0.6725335, 
    -0.5812092, -0.6033278, -0.6654863, -0.7843013, -0.7962971, -0.8102942, 
    -0.7447019, -0.3707099, -0.1725655, -0.1066475, -0.1011629, -0.007673264, 
    -0.03457785, -0.005313396, -0.06919718, -0.00217247, -0.08488703, 
    -0.1381414, 0.0974865, 0.1108003, 0.1202729, 0.02100538, 0.0004650056, 
    0.05396436, -0.117341, -0.3209542, -0.3393462, -0.2253813, -0.02380258, 
    -0.31516, -0.1588449, 0.0950613, 0.2174411, 0.37675, 0.3870201, 
    0.4469161, 0.4350514, 0.4156671, 0.3985114, 0.3671966,
  0.1399507, 0.05064398, 0.006780148, 0.02019191, 0.03378248, 0.008359432, 
    -0.09427774, -0.136921, 0.02637655, -0.002057761, -0.0959053, 
    -0.06667352, -0.365339, -0.6110747, -0.4185454, -0.5124745, -0.330964, 
    0.2072521, 0.5938732, 0.9362723, 1.056845, 1.083424, 1.135703, 1.236679, 
    1.180153, 1.277776, 1.119947, 1.055283, 0.6877863, 0.1938729, 
    0.001799583, -0.2076077, -0.3359771, -0.2362056, 0.2371182, 0.5990167, 
    0.92942, 0.8432703, 0.2956961, 0.190846, 0.336484, 0.6921154, 0.9244885, 
    1.263128, 1.099049, 0.8072359, 0.6070405, 0.1946056, -0.5179105, 
    -0.8327541, -1.024942, -1.152757, -1.06337, -1.244116, -1.016967, 
    -0.8598866, -0.5367751, -0.4671459, -0.4100337, -0.1968985, -0.1361732, 
    -0.1674228, -0.261075, -0.2018957, -0.1312742, 0.09344959, 0.1156497, 
    0.05970955, 0.04816961, -0.02920675, -0.03757262, -0.07269597, 
    -0.1242256, -0.151016, -0.1319894, -0.1586494, -0.02868538, -0.05778694, 
    -0.05161832, -0.1231841, -0.1628813, -0.2485584, -0.3006905, -0.5209217, 
    -0.4223213, -0.08947623, -0.06573033, -0.1578522, -0.0925045, 0.06464148, 
    0.1937747, 0.2254643, 0.2046316, 0.2729583, 0.1802177, 0.1795828,
  0.06648064, 0.006584883, 0.08070612, 0.04810524, 0.170012, 0.09043932, 
    0.01136994, 0.006828845, 0.1261323, 0.2385021, 0.4238541, 0.1839609, 
    -0.05171561, -0.03882536, 0.1617931, 0.04358011, -0.1939524, -0.04930699, 
    0.2731538, 0.4982189, 0.5899344, 0.6735933, 0.7589937, 0.8928153, 
    0.8673272, 0.9684339, 0.7680595, 0.3008723, -0.05567098, -0.2696366, 
    -0.4467361, -0.5073478, -0.3797114, -0.2744532, 0.160181, 0.6097584, 
    0.5621514, 0.06469023, -0.00607796, 0.1431733, 0.4496351, 0.3887461, 
    0.2046967, 0.5285575, 0.659075, 0.4147065, 0.002222836, -0.2920155, 
    -0.736921, -0.9509182, -0.8964424, -0.8771555, -0.6432526, -0.6029372, 
    -0.5364823, -0.5159249, -0.2478261, -0.0645256, 0.004468918, 0.2185965, 
    0.361711, 0.4668384, 0.4702563, 0.4416757, 0.4365163, 0.4933686, 
    0.5220957, 0.3699629, 0.3391526, 0.2071373, 0.1317966, -0.09172225, 
    -0.1296945, -0.1948149, -0.2761626, 0.07066357, 0.1274507, -0.05344124, 
    -0.03830452, 0.01327425, 0.01319289, -0.1476633, -0.1021391, -0.3925036, 
    -0.5399971, -0.2002999, -0.119652, -0.09888458, -0.252969, -0.1880603, 
    -0.05700541, 0.004745722, 0.004452705, 0.08869743, -0.0642648, 0.02211215,
  0.02362597, 0.06125617, 0.06888986, 0.09943962, 0.06623673, -0.01662493, 
    -0.03369839, -0.1037993, 0.09213167, 0.4748952, 0.7719817, 0.0005943775, 
    0.05064344, 0.42291, 0.4254162, 0.4766694, 0.2607677, 0.0883068, 
    0.1206148, 0.1550223, 0.1326753, 0.2828055, 0.2163667, 0.2525158, 
    0.3507417, 0.1379325, 0.06713152, -0.01856169, -0.2623442, -0.2396393, 
    -0.01403707, -0.09883513, -0.07505582, -0.1123117, 0.1664155, 0.1430106, 
    0.02043572, -0.01162808, 0.1416597, 0.3331798, 0.06355095, -0.1451893, 
    -0.1313219, 0.04810512, -0.1172104, -0.362165, -0.5634999, -0.826798, 
    -1.118155, -1.229353, -1.168546, -1.050415, -0.8489656, -0.6383047, 
    -0.465209, -0.2203035, -0.06932688, 0.04286385, 0.1448336, 0.2778082, 
    0.4264092, 0.5571542, 0.6971283, 0.7066658, 0.7476649, 0.7760503, 
    0.8296478, 0.6683202, 0.5885184, 0.4505137, 0.3170503, 0.1213146, 
    -0.04844451, -0.2673411, -0.2777251, 0.06374645, 0.257838, 0.1275809, 
    0.03122672, -0.002676278, 0.04847935, -0.2015369, -0.1557038, -0.342227, 
    -0.2788806, -0.2068756, -0.2605708, -0.06096029, -0.2024809, -0.2427151, 
    -0.2473704, -0.06935921, -0.136449, -0.06164438, -0.07406294, 0.009579659,
  0.03112924, 0.09524059, -0.06061959, 0.05983996, 0.05914012, -0.01662484, 
    0.001848474, 0.03093376, 0.4689871, 0.4724706, 0.6647549, 0.2974212, 
    0.1164966, 0.330657, 0.44594, 0.454567, 0.3377538, 0.3543718, 0.1942642, 
    0.1537044, 0.07520509, 0.1441336, 0.08104777, -0.02264708, -0.03906949, 
    -0.3165596, -0.1588449, -0.1155506, -0.6118721, -0.3817289, 0.02313751, 
    0.007626459, -0.01921272, 0.02227497, 0.1141374, 0.3232183, 0.3557053, 
    0.3552337, 0.2949967, 0.3508229, 0.2089448, 0.04952049, -0.004059792, 
    0.03368378, -0.05886173, -0.2627025, -0.4642811, -0.6025462, -0.6259189, 
    -0.6798739, -0.7502842, -0.7328033, -0.7910876, -0.7612538, -0.8397369, 
    -0.7977448, -0.6709871, -0.4847732, -0.2693758, -0.1985912, -0.111661, 
    -0.03244591, 0.1607838, 0.2022879, 0.3204188, 0.4773686, 0.6533782, 
    0.7282643, 0.7936457, 0.7596447, 0.6096445, 0.4688894, 0.2628837, 
    0.01299787, -0.01439452, 0.200937, 0.4286388, 0.1259533, 0.1154227, 
    0.03241485, -0.1415108, -0.1357329, -0.466527, -0.4806547, -0.4287186, 
    -0.2995195, -0.2338285, -0.06063604, -0.1031978, -0.03718138, -0.044994, 
    -0.04805386, -0.08674201, 0.1979262, 0.09030879, -0.004238605,
  0.02247022, -0.01013067, 0.118336, 0.01516227, 0.1573497, 0.1626557, 
    0.1405854, 0.2333752, 0.3404715, 0.01618767, 0.1329844, 0.5501883, 
    0.2604585, 0.2054772, 0.4477949, 0.5421314, 0.4718513, 0.4499111, 
    0.2113214, 0.2561131, 0.343401, 0.1156178, 0.07097244, 0.06571531, 
    -0.07088971, -0.1268135, -0.06296271, -0.2510322, -0.5308995, -0.1679764, 
    0.05456614, 0.03560519, 0.1165782, 0.2668059, 0.3533125, 0.6041594, 
    0.6636643, 0.5427332, 0.5002203, 0.518271, 0.4100184, 0.2119393, 
    -0.03853273, -0.1435943, -0.2238026, -0.3085356, -0.3925695, -0.4654536, 
    -0.467114, -0.4082108, -0.3359609, -0.3070383, -0.3981032, -0.5184321, 
    -0.6717038, -0.8346105, -0.9268632, -1.043107, -1.065535, -1.024503, 
    -0.8515205, -0.7155352, -0.5288806, -0.3723221, -0.1618233, 0.1328869, 
    0.4441981, 0.7701421, 0.9597092, 0.9864349, 0.8753667, 0.8902924, 
    0.7376392, 0.516497, 0.4725354, 0.1731213, 0.8555918, -0.07399774, 
    0.05910754, -0.2065336, -0.4032946, -0.5573969, -0.5692301, -0.3633375, 
    -0.3269448, -0.1289301, -0.1024165, 0.02006149, 0.0757575, 0.2486742, 
    0.3221126, 0.3608003, 0.6192964, 0.6924411, 0.1464123, 0.009563319,
  0.03272414, 0.02313757, 0.05796838, 0.08451486, 0.1409111, 0.09292924, 
    0.1425064, 0.1868587, 0.1566499, 0.3375582, 0.2464122, 0.1937594, 
    0.0166266, 0.005298138, 0.1633229, 0.3851161, 0.4014568, 0.3509531, 
    0.4034104, 0.5445075, 0.6864345, 0.03272367, -0.124486, -0.007071018, 
    -0.2667394, -0.294116, -0.3875403, -0.3459873, -0.2977452, -0.1771398, 
    0.1909428, 0.365211, 0.3399825, 0.2178645, 0.2293868, 0.3787355, 
    0.4404063, 0.4394298, 0.4645596, 0.3388758, 0.2277265, 0.1463308, 
    0.04650974, 0.06350136, -0.0209713, -0.04937363, -0.06171131, 
    -0.06311035, -0.05207539, -0.0665617, -0.04904842, -0.1163979, 
    -0.08337307, -0.1604567, -0.1502028, -0.2371168, -0.4535069, -0.651114, 
    -0.6196527, -0.5755935, -0.676847, -0.6345129, -0.4607177, -0.3785067, 
    -0.2883863, 0.06093025, 0.3161058, 0.7293062, 1.150741, 1.327792, 
    1.356877, 1.612184, 1.123545, 0.243824, 0.1528413, 0.2770275, 0.4849213, 
    -0.1971593, -0.2724843, -0.5979724, -0.5834384, -0.395597, -0.5439849, 
    -0.222827, -0.2774167, -0.2137775, -0.1563554, 0.04800653, 0.1970954, 
    0.4682541, 0.6860926, 1.062232, 1.192945, 0.5565522, 0.09512663, 
    0.06050742,
  -0.09165692, -0.09405065, -0.02839279, -0.1452057, -0.1610098, -0.1041088, 
    0.06203699, 0.1742604, 0.2817312, 0.5745047, 0.2822847, -0.06992865, 
    -0.1301823, -0.07969499, -0.02028751, 0.05788612, 0.2174077, 0.4044032, 
    0.4981213, 0.4917409, 0.3920176, -0.1560457, -0.1815991, -0.1159253, 
    -0.3822989, -0.3422108, -0.3902094, -0.1363188, -0.2425196, -0.002887487, 
    0.2818613, 0.03542519, 0.01602459, -0.06312633, -0.04444122, 0.2147064, 
    0.3031826, 0.3079839, 0.2650642, 0.3058681, 0.2963791, 0.2049074, 
    0.06975174, -0.01553535, 0.002335548, 0.002205849, -0.03068924, 
    0.04590702, 0.1910725, 0.197258, 0.2510986, 0.234107, 0.2797613, 
    0.2341881, 0.1860104, 0.07884979, -0.002155304, -0.07544708, -0.1516848, 
    -0.1324291, -0.1359453, 0.005770206, 0.09493065, 0.05708885, 0.1021085, 
    0.2832122, 0.3498464, 0.7861257, 1.330055, 1.638371, 1.579078, 1.348186, 
    0.7174566, 0.218677, 0.7494559, 0.8705654, 0.6847744, 0.05069351, 
    -0.2665768, -0.3846102, -0.3457108, -0.287703, -0.2584715, -0.2767334, 
    -0.382853, -0.3041091, -0.2051015, -0.08980227, 0.04618359, 0.3791914, 
    0.6550221, 1.031519, 0.5489842, 0.1393642, 0.03296757, 0.07813454,
  -0.09300852, -0.0416255, -0.002855301, -0.1140528, -0.2112536, -0.2018628, 
    -0.01174259, 0.1768317, 0.3036062, 0.4961518, 0.3649506, 0.006177902, 
    -0.1572011, -0.08327508, -0.1496325, -0.2442126, -0.2207913, 0.1458263, 
    0.3399661, 0.4628022, 0.3639579, -0.3345768, -0.3810779, -0.1796457, 
    -0.2806872, -0.3399483, -0.2960194, -0.326504, -0.2819896, 0.1444106, 
    -0.04421329, -0.5247788, -0.3148022, -0.2754798, -0.4427648, -0.3044834, 
    -0.1872311, -0.1403718, -0.2237215, -0.1871982, -0.180346, -0.1463284, 
    -0.124877, -0.2429109, -0.2277741, -0.1671295, 0.07123232, 0.1423268, 
    0.2565198, 0.400188, 0.4369884, 0.5183196, 0.6552987, 0.7438407, 
    0.7259531, 0.6766539, 0.5815682, 0.3992281, 0.2072029, 0.1707926, 
    0.1953545, 0.3303633, 0.3594818, 0.3464613, 0.3425055, 0.3240161, 
    0.4290133, 0.5778742, 0.5665781, 0.4179454, 0.2542249, -0.2073473, 
    -0.02144253, 0.7973723, 1.232073, 1.066171, 0.8205814, 0.3860273, 
    0.03415537, 0.09239149, -0.04808664, -0.3241124, -0.3735595, -0.5429602, 
    -0.5311923, -0.5251379, -0.494441, -0.32587, -0.02575636, 0.3036542, 
    0.6546474, 1.004159, 0.3706791, 0.2078214, 0.1123459, -0.02536559,
  0.1179297, 0.02821493, -0.1109121, -0.1308172, -0.1928945, -0.2665758, 
    -0.1308823, 0.09737301, 0.1906831, 0.2643484, 0.538958, 0.1040294, 
    -0.3676348, -0.1433662, -0.06387418, -0.3978422, -0.544832, -0.0137279, 
    0.1567957, 0.03482318, -0.1418037, -0.3133534, -0.2961823, -0.3499907, 
    -0.6960357, -0.190632, -0.02533251, -0.219115, -0.1304431, 0.1293875, 
    -0.2819085, -0.6680417, -0.7965894, -0.7956457, -0.9615636, -0.8050036, 
    -0.7179279, -0.7634192, -0.7305412, -0.614819, -0.4806385, -0.50948, 
    -0.5461497, -0.4817452, -0.29003, -0.2491932, -0.2064033, -0.1906972, 
    0.129941, 0.4371176, 0.5921803, 0.8859949, 1.060442, 1.151343, 1.143531, 
    1.062217, 0.8559828, 0.7021418, 0.652988, 0.6078053, 0.539495, 0.5190682, 
    0.5159926, 0.5030036, 0.4287362, 0.4176846, 0.5631441, 0.3882582, 
    0.2479748, 0.30595, 0.133945, -0.02171922, 0.4187105, 1.00258, 0.8475184, 
    0.635572, 0.6009855, 0.4509201, 0.152873, -0.01330471, -0.1918688, 
    -0.3692942, -0.4417062, -0.5359774, -0.5509028, -0.6661367, -0.5536537, 
    -0.3363681, -0.1439528, 0.1041589, 0.5002527, 0.8167572, 0.3609135, 
    0.2394781, 0.1516366, 0.1427495,
  -0.003733635, -0.134886, -0.4026599, -0.450837, -0.6112047, -0.5667713, 
    -0.2112701, -0.1509348, 0.03929967, 0.09792596, -0.05565476, -0.3599353, 
    -0.3484933, -0.01585984, -0.1000233, -0.3665435, -0.199356, 0.2644624, 
    0.02079391, -0.1451077, -0.3143136, -0.281957, -0.2825103, -0.7320546, 
    -0.7365468, -0.01218152, -0.08200568, -1.012523, -0.2631581, 0.2261, 
    -0.1221912, -0.1160712, -0.2296131, -0.3300691, -0.5037508, -0.4997308, 
    -0.5621333, -0.7173243, -0.7432035, -0.9208401, -0.9887438, -1.021947, 
    -0.8030666, -0.6240953, -0.544831, -0.4208566, -0.3617094, -0.2065659, 
    0.05601549, 0.2393489, 0.6040134, 0.9635673, 1.083587, 1.286028, 
    1.347275, 1.184938, 0.9854903, 0.8727627, 0.7134686, 0.6673427, 
    0.6934013, 0.6103444, 0.5841393, 0.524863, 0.514267, 0.5537691, 
    0.4472749, 0.1889741, 0.3058035, 0.4584728, 0.168564, 0.3519461, 
    0.9724051, 0.9345469, 0.5937586, 0.5441172, 0.3868251, 0.116122, 
    -0.05103302, -0.1669176, -0.2803292, -0.4082754, -0.5595117, -0.6510494, 
    -0.628181, -0.6091866, -0.439949, -0.2948968, -0.106029, 0.2277761, 
    0.4777107, 0.5865002, 0.3119717, 0.07157493, -0.01804161, -0.004320383,
  -0.2915596, -0.5302316, -0.7337959, -0.6081775, -0.7957428, -0.6518788, 
    -0.3201731, -0.4035714, -0.09907925, 0.02391878, -0.3874744, -0.3850819, 
    -0.04631233, -0.08718146, -0.3536854, -0.2591054, 0.1236747, 0.04439408, 
    0.004289865, 0.1109468, 0.05515251, 0.1339285, 0.1042736, -0.4088938, 
    -0.07516968, 0.7350845, -0.001520634, -0.8075265, 0.1728113, 0.2442153, 
    -0.01817095, 0.1694919, -0.156729, -0.1538801, -0.01745462, -0.02774137, 
    -0.1340728, -0.2347889, -0.3179269, -0.5048085, -0.5742582, -0.7781971, 
    -0.7275784, -0.6107328, -0.5684478, -0.2335193, 0.0584892, 0.3069593, 
    0.4626559, 0.5742282, 0.774277, 0.8003676, 0.9827894, 1.120973, 
    0.8806734, 0.7194917, 0.6485119, 0.5591238, 0.5042572, 0.5850677, 
    0.6259532, 0.6084077, 0.60888, 0.4991955, 0.5723724, 0.5953869, 
    0.3885184, 0.4140556, 0.3279227, 0.03034782, -0.1985748, 0.08776969, 
    0.4665298, 0.4740007, 0.2748465, 0.3461193, 0.2241466, -0.03397509, 
    -0.3251047, -0.5847726, -0.6843007, -0.7717518, -0.9031157, -0.8993235, 
    -0.681078, -0.5066639, -0.4161528, -0.07538104, 0.3816504, 0.6060481, 
    0.5918386, 0.5974207, 0.4967213, 0.04734039, -0.1298735, -0.1719143,
  -0.3656645, -0.5955311, -0.7218495, -0.6990629, -0.9230052, -1.115844, 
    -0.5196031, -0.4176335, -0.4955313, -0.3814686, -0.3133533, -0.0923247, 
    -0.1097075, -0.454076, -0.5333403, 0.04224569, -0.09992561, -0.4219308, 
    0.02842712, 0.1864678, 0.1089776, 0.5213147, 0.6975188, 0.1456795, 
    0.1634369, 0.2972741, -0.5621982, -0.2268624, 0.5108483, 0.1503511, 
    -0.04932344, 0.1002536, 0.07084262, 0.1493257, 0.3402437, 0.3043387, 
    0.1647555, 0.01355124, -0.1200273, -0.2696362, -0.2340083, -0.2061758, 
    -0.05170012, 0.1760182, 0.2779222, 0.3628674, 0.4973888, 0.7702885, 
    0.955689, 1.103378, 1.099212, 0.909596, 0.9541109, 0.8307545, 0.5822194, 
    0.5790622, 0.4014742, 0.2103935, 0.2358655, 0.3321057, 0.4266044, 
    0.5450125, 0.5027925, 0.3109956, 0.3266858, 0.1307222, 0.05402946, 
    0.3320405, 0.1618258, -0.07842505, 0.07290971, 0.1459891, 0.1648856, 
    0.1623628, 0.07826436, -0.03433299, -0.1816963, -0.2841864, -0.3746977, 
    -0.4736569, -0.5703366, -0.755769, -0.8042226, -0.6560776, -0.4512274, 
    -0.3156972, -0.1359766, 0.3266369, 0.6665294, 0.6973563, 0.7094655, 
    0.6253185, 0.2908621, 0.03308201, -0.02904344, -0.1354237,
  -0.2704822, -0.3658106, -0.4756744, -0.2367911, -0.3634355, -0.5018463, 
    -0.1862863, -0.1423084, -0.5127845, -0.3554434, -0.00484097, -0.1317941, 
    -0.4089426, -0.3566149, -0.101179, -0.04178759, -0.2767648, -0.2666411, 
    0.08472609, 0.1036389, 0.04525667, 0.3075943, 0.2038178, 0.2741628, 
    0.1808677, -0.1347082, -0.08301544, 0.2915458, 0.2082124, -0.01227909, 
    0.03002229, 0.2448172, 0.3834893, 0.3865488, 0.1083908, 0.1325936, 
    0.08601201, -0.01587558, 0.147193, 0.316545, 0.3931408, 0.6109467, 
    0.7600346, 0.7256598, 0.7700281, 0.8777919, 1.006747, 1.202287, 1.271493, 
    1.345142, 1.369003, 1.268368, 1.145696, 0.9009209, 0.7449474, 0.561142, 
    0.2587652, 0.2202725, 0.2159591, 0.0918386, 0.1069758, 0.08835602, 
    -0.00962615, -0.03488654, -0.07565805, -0.1490629, -0.1653553, -0.15502, 
    -0.3291087, -0.05301762, 0.2670178, 0.2663668, 0.2103935, 0.1106377, 
    -0.08736038, -0.09953475, -0.2023025, -0.3061762, -0.3447666, -0.3487544, 
    -0.3363523, -0.3976474, -0.3697338, -0.160522, 0.1148686, 0.342001, 
    0.5167732, 0.6896739, 0.7816668, 0.7961519, 0.7672783, 0.6667087, 
    0.6610935, 0.6868747, 0.3812919, -0.1017323,
  0.06270456, 0.1892667, 0.3764248, 0.6344655, 0.6077569, 0.5075614, 
    0.3801851, 0.1040946, -0.1551338, 0.06895459, 0.1962007, -0.02455127, 
    -0.165583, -0.08495176, -0.01418342, -0.2674061, -0.06877327, 0.2814546, 
    0.005315244, 0.03119409, 0.2681413, 0.09139943, -0.1440174, 0.003899276, 
    0.2337658, 0.2871675, 0.5996351, 0.4161065, 0.003899336, 0.04828429, 
    0.172291, 0.1219983, 0.274863, 0.5129814, 0.5711679, 0.3908782, 
    0.4361744, 0.4307709, 0.6086345, 0.9691982, 1.081455, 1.06858, 0.9726162, 
    0.951262, 1.130299, 1.31565, 1.419914, 1.54843, 1.708049, 1.860034, 
    1.791481, 1.592652, 1.417376, 1.155559, 0.8805757, 0.5627041, 0.2394295, 
    0.1041265, -0.1252513, -0.2769928, -0.3111405, -0.5515215, -0.5454985, 
    -0.3354887, -0.3451405, -0.2981515, -0.08547246, -0.155638, -0.4264402, 
    -0.02035213, 0.4673109, 0.3769791, 0.2357515, 0.04388976, -0.09922576, 
    0.003443956, -0.1490142, -0.29213, -0.2497792, -0.259089, -0.2743726, 
    -0.1468825, 0.101213, 0.3931074, 0.6554613, 0.7635508, 0.7540131, 
    0.7827892, 0.9632416, 1.190911, 1.108896, 0.9920497, 1.063111, 0.8295178, 
    0.2303153, 0.0220471,
  0.1420822, 0.2086837, 0.6723075, 0.793206, 0.5725679, 0.4209566, 0.2251721, 
    0.07416296, 0.07058215, 0.2277275, 0.2592542, 0.1964613, -0.007103324, 
    -0.114216, 0.1977959, 0.164023, 0.3080333, 0.3832449, 0.2051525, 
    0.1279228, 0.1149018, 0.0225352, 0.06488568, 0.1968844, 0.01760364, 
    -0.04750049, 0.2933197, 0.2524834, 0.09592438, 0.2605398, 0.2881112, 
    0.1572032, 0.2613204, 0.4353764, 0.2560966, 0.1174893, 0.3934493, 
    0.7652917, 1.197405, 1.179355, 1.452613, 1.480331, 1.385995, 1.514446, 
    1.701604, 1.806356, 1.972682, 2.051783, 2.020012, 2.008912, 1.939234, 
    1.775872, 1.64454, 1.437753, 1.173268, 0.8360281, 0.4657645, 0.2069426, 
    -0.03734493, -0.2134514, -0.5579019, -1.059122, -0.9876211, -0.4280832, 
    -0.3350331, -0.3341866, -0.4782298, -0.6821361, -0.4570875, 0.1351814, 
    0.291008, 0.01551962, -0.05402732, 0.04375863, 0.1725998, 0.2498953, 
    0.150856, 0.06890512, 0.2891202, 0.3396082, 0.2307868, 0.2622809, 
    0.3994064, 0.5201583, 0.6790619, 0.8416591, 1.012037, 1.103785, 1.2622, 
    1.466529, 1.421005, 1.200888, 0.9600353, 0.5572197, 0.1707287, 0.1941173,
  -0.02503943, 0.05764276, 0.4605075, 0.3377373, 0.1504975, 0.3134534, 
    0.396152, 0.1896579, 0.229176, 0.3023366, 0.3930595, 0.5353935, 
    0.5800388, 0.5618745, 0.6994233, 0.5272227, 0.2991629, 0.2647879, 
    0.3821707, 0.2867443, 0.06192334, 0.01692009, 0.03856723, 0.03200798, 
    -0.02352588, 0.05090442, 0.3117123, 0.4638436, 0.3577075, 0.223707, 
    0.1970305, 0.3105068, 0.2883224, 0.3205495, 0.3641851, 0.2763438, 
    0.3083906, 0.7753181, 1.137672, 1.369605, 1.56622, 1.596346, 1.56246, 
    1.763616, 1.953525, 1.901718, 1.764104, 1.662525, 1.592391, 1.658261, 
    1.745565, 1.628166, 1.299862, 0.8978765, 0.5487878, 0.1607509, 
    -0.1699781, -0.3743567, -0.5528235, -0.8627348, -1.222419, -1.311595, 
    -1.000853, -0.4120674, -0.2191476, -0.1544502, -0.2357335, -0.2127676, 
    0.0630784, 0.3285892, 0.2981215, 0.1885999, 0.3924248, 0.4977307, 
    0.2725028, 0.1442964, 0.06942642, 0.07522094, 0.146266, 0.3604259, 
    0.341496, 0.4734297, 0.4830494, 0.6206307, 0.8597913, 0.8703051, 
    0.6572523, 0.4941335, 0.5726323, 0.6688404, 0.5396576, 0.3390875, 
    0.2556734, 0.2173433, 0.2623143, 0.1941819,
  -0.1604557, 0.08550715, 0.3415451, 0.1623621, 0.06783152, 0.3271906, 
    0.3109796, 0.1037204, 0.1868907, 0.3594005, 0.4759696, 0.5479747, 
    0.614853, 0.4547131, 0.1887951, -0.003229648, -0.1992908, -0.2776925, 
    -0.2996489, -0.3340403, -0.1731515, -0.007363766, 0.04393834, 
    -0.04203174, -0.00178051, 0.07430887, 0.2289472, 0.2176199, 0.1658297, 
    0.1200445, 0.225286, 0.08980417, -0.1000724, 0.08088446, 0.331763, 
    0.08034706, 0.07302284, 0.6045339, 1.588892, 1.403296, 0.8906016, 
    0.8773198, 1.01386, 1.194492, 1.313909, 1.240944, 1.090585, 1.060752, 
    1.144687, 1.23318, 1.195452, 1.007285, 0.6739839, 0.283831, -0.1207261, 
    -0.5341055, -0.8612051, -1.08085, -1.231663, -1.39737, -1.427823, 
    -1.085652, -0.5166247, -0.3433014, -0.2309315, -0.1216538, 0.2378187, 
    0.5281177, 0.6292732, 0.5909765, 0.4560966, 0.4400483, 0.4247977, 
    0.3858981, 0.3965915, 0.3155042, 0.1420015, 0.01540637, 0.01892209, 
    0.1386162, 0.3566504, 0.4276298, 0.3078375, 0.4923592, 0.7136157, 
    0.5802827, 0.2879, 0.2310309, 0.2940192, 0.1891365, 0.01138639, 
    -0.03296661, -0.06893659, -0.1953366, -0.2716384, -0.2645586,
  -0.1055734, -0.1200273, -0.04566145, -0.2039945, -0.3783758, -0.450886, 
    -0.4135482, -0.2724029, -0.04359424, 0.2063407, 0.2208263, 0.1206799, 
    0.05489206, -0.005817533, -0.1586171, -0.249535, -0.3188384, -0.3223048, 
    -0.3928614, -0.3538809, -0.1581132, -0.0164783, -0.04541707, 
    -0.005117416, 0.0654068, -0.01236033, -0.09367537, -0.1015694, 
    -0.2000885, -0.2418686, -0.183748, -0.2794347, -0.129158, 0.07274711, 
    0.0737561, -0.03241205, 0.3564708, 1.342066, 1.424276, 0.5356369, 
    -0.4565988, -0.2151925, 0.1475353, 0.1073173, -0.0181222, 0.1876234, 
    0.6106702, 0.9276623, 1.125758, 1.170598, 1.103671, 0.9345796, 0.5768159, 
    0.04187126, -0.6294016, -1.206452, -1.571752, -1.64615, -1.435928, 
    -1.160261, -0.8858467, -0.5840731, -0.1587145, 0.03038038, 0.08731401, 
    0.2760837, 0.694638, 0.8770113, 0.7276624, 0.5617445, 0.5859143, 
    0.6794202, 1.045094, 1.409075, 1.623984, 1.396591, 0.347926, -0.07808334, 
    -0.0584054, 0.07699513, 0.02395105, -0.005801916, -0.1811924, 0.09069872, 
    0.1661546, -0.00646925, -0.123852, -0.1153228, -0.2275462, -0.4149976, 
    -0.4034576, -0.2144444, -0.1756263, -0.2361073, -0.1370674, -0.06395543,
  -0.924356, -1.000625, -0.8594146, -0.8201405, -0.9117908, -1.201667, 
    -1.010505, -0.5588124, -0.199893, -0.1045806, -0.05458057, -0.09520561, 
    -0.05956101, -0.04960009, -0.1523019, -0.3400136, -0.4025135, -0.4250231, 
    -0.2913315, -0.1683986, -0.1143625, -0.2025294, -0.3523347, -0.3138254, 
    -0.1896229, -0.1676339, -0.1413968, -0.2096423, -0.1996, -0.1891832, 
    -0.2551508, -0.4340243, -0.4690669, -0.3382552, -0.2018623, -0.01516056, 
    0.3934169, 0.4693131, -0.2294178, -1.509773, -2.285261, -1.674063, 
    -0.3854396, -0.1637601, -0.1092358, 0.3613205, 0.7384202, 0.9165614, 
    1.026442, 1.091106, 0.8514252, 0.2866142, -0.4610419, -1.198835, 
    -1.700544, -1.902692, -1.90891, -1.580801, -1.038272, -0.5562246, 
    -0.457608, 0.009563446, 0.3437755, 0.424228, 0.4449638, 0.430478, 
    0.5348238, 0.5376884, 0.3682711, 0.3075615, 0.4525156, 0.7507255, 
    0.9246669, 0.9460219, 0.5390394, -0.1572498, -0.8757557, -0.9196848, 
    -0.4782131, -0.2284257, -0.1091549, -0.6714921, -0.7890693, -0.6150135, 
    -0.7837473, -1.050121, -1.094115, -0.9123443, -0.7638087, -0.7074614, 
    -0.6270905, -0.6089588, -0.6994532, -0.7261949, -0.6453357, -0.6524481,
  -1.972419, -1.813679, -1.160098, -0.7935942, -0.771166, -0.9972564, 
    -0.7491118, -0.5395904, -0.3365141, -0.21988, -0.192341, -0.2285063, 
    -0.2481841, -0.2567127, -0.3028065, -0.3617909, -0.4278227, -0.4800202, 
    -0.4622303, -0.3309966, -0.2697011, -0.2654855, -0.3187408, -0.3067941, 
    -0.2567616, -0.2582753, -0.2463775, -0.2535062, -0.2814196, -0.310472, 
    -0.4230051, -0.6210032, -0.5174062, -0.1800851, 0.05712199, 0.1197522, 
    0.008879721, -0.1628, -0.4690824, -0.6628163, -0.5656483, -0.3342357, 
    -0.1698472, -0.1134343, -0.05832362, -0.06232858, -0.2893143, -0.992439, 
    -1.162215, -1.265323, -1.525789, -1.950837, -1.658747, -1.689183, 
    -1.36158, -0.8616279, -0.5220282, -0.274616, -0.03316092, 0.09393847, 
    0.201409, 0.3252534, 0.3972262, 0.3738699, 0.2510835, 0.2237071, 
    0.1704032, 0.1391206, 0.2288668, 0.3077079, 0.4852633, 0.3335054, 
    0.1777924, -0.1902414, -0.600772, -0.9077544, -0.9915596, -0.7982004, 
    -0.5636952, -0.5194732, -0.8406318, -1.32683, -1.511758, -1.351456, 
    -1.33697, -1.669815, -1.60458, -1.280329, -1.00834, -0.930427, 
    -0.9969472, -1.171898, -1.352221, -1.49584, -1.617211, -1.817553,
  -2.088598, -2.100284, -1.889428, -1.324975, -1.008812, -0.8480377, 
    -0.6358957, -0.6663808, -0.5614817, -0.4879791, -0.4307362, -0.4357655, 
    -0.5092844, -0.6175201, -0.7199941, -0.7669667, -0.7249094, -0.7690012, 
    -0.7060781, -0.6224517, -0.5464587, -0.4831288, -0.4621001, -0.455313, 
    -0.4430408, -0.4924061, -0.5411366, -0.5637928, -0.5802151, -0.5452543, 
    -0.4666246, -0.3611723, -0.1579009, -0.006712722, -0.004466623, 
    -0.1817778, -0.4877836, -0.559561, -0.5656483, -0.3287343, -0.121231, 
    -0.1502838, -0.2446848, -0.4067125, -0.4939846, -0.5544989, -0.5949612, 
    -0.6650624, -0.7213776, -0.8418363, -1.085082, -1.619929, -1.372159, 
    -1.055915, -0.6186593, -0.3389229, -0.07028675, -0.01940811, 0.008440256, 
    0.04416618, 0.02040315, 0.03571892, 0.0339611, -0.05324593, -0.1417225, 
    -0.1561105, -0.09767953, -0.04528695, 0.004322469, 0.05246705, 
    0.005282715, -0.1460194, -0.3019764, -0.4543039, -0.5469309, -0.5622954, 
    -0.5547108, -0.4771391, -0.4014231, -0.4932686, -0.8759669, -1.059968, 
    -0.7579821, -0.8503332, -1.085636, -0.84532, -0.7346425, -0.696476, 
    -0.4768143, -0.3986402, -0.5601475, -0.8794346, -1.035147, -1.283552, 
    -1.560131, -1.856957,
  -1.560033, -1.585717, -1.571931, -1.480883, -1.273331, -0.8268462, 
    -0.6601633, -0.4470124, -0.2614816, -0.1601957, -0.1605864, -0.2074612, 
    -0.2584707, -0.4944406, -0.7861887, -0.8618557, -0.8721426, -0.8412992, 
    -0.7675686, -0.7278227, -0.6932036, -0.6845937, -0.7167551, -0.726423, 
    -0.7423897, -0.741869, -0.7064356, -0.6392157, -0.5261624, -0.380687, 
    -0.2378812, -0.1740142, -0.2039783, -0.265339, -0.2363352, -0.3330636, 
    -0.3547922, -0.2482327, -0.1577543, -0.03945994, -0.03487015, -0.1015042, 
    -0.1273833, -0.09618212, -0.05502002, -0.05759162, -0.06211637, 
    -0.007965982, -0.04032266, -0.2165597, -0.4838937, -0.8185128, 
    -0.9176993, -0.941267, -0.7296622, -0.5110257, -0.3472239, -0.2728748, 
    -0.2083403, -0.1337147, -0.09588915, -0.0731352, -0.1329985, -0.2266997, 
    -0.2398019, -0.187507, -0.07219112, 0.04335243, 0.1022066, 0.02689737, 
    -0.1022368, -0.2391834, -0.3014068, -0.2445382, -0.2976307, -0.2410226, 
    -0.2042224, -0.1556873, -0.2062243, -0.3737371, -0.3473703, -0.5032622, 
    -0.5406485, -0.7724688, -0.9826088, -0.9108467, -0.8335356, -0.601895, 
    -0.6068429, -0.5238513, -0.6032947, -0.8319407, -1.272224, -1.381648, 
    -1.456745, -1.536612,
  -1.319766, -1.056029, -0.7513416, -0.4493558, -0.1889719, 0.0402925, 
    0.2334566, 0.3293712, 0.3294689, 0.2442476, 0.1297781, -0.04976296, 
    -0.2285389, -0.4116281, -0.3158435, -0.1875558, -0.279727, -0.237979, 
    -0.1763905, -0.115925, -0.1464913, -0.2202707, -0.3304595, -0.4435943, 
    -0.553718, -0.6384994, -0.621052, -0.5304432, -0.3925853, -0.2074773, 
    -0.09963226, -0.03967154, -0.06820345, -0.1160388, -0.1533597, 
    -0.2549219, -0.1565174, -0.07420933, 0.03523076, 0.04717726, -0.04325247, 
    -0.01810595, 0.002645999, 0.02071241, 0.02006137, -0.03198941, 
    -0.1040272, -0.1772856, -0.2440011, -0.3284901, -0.4328194, -0.5198799, 
    -0.5926175, -0.6111071, -0.5685617, -0.4901599, -0.4300853, -0.4122791, 
    -0.4114328, -0.4233957, -0.4211822, -0.4192128, -0.3281646, -0.3754953, 
    -0.3319406, -0.2692615, -0.2273507, -0.2195057, -0.2329985, -0.3344145, 
    -0.2847401, -0.2990955, -0.4155669, -0.3111724, -0.2493072, -0.2198149, 
    -0.2697824, -0.4917387, -0.4257882, -0.3657296, -0.4554919, -0.340632, 
    -0.3078356, -0.4246492, -0.562865, -0.6253163, -0.6815176, -0.5426021, 
    -0.1745844, 0.01836801, -0.01996112, -0.2107331, -0.5188384, -0.8587798, 
    -1.258112, -1.39029,
  -0.9986559, -0.6984931, -0.2013576, 0.2733166, 0.5065196, 0.4970305, 
    0.08957624, 0.06991434, -0.05047846, -0.08469081, -0.1834054, -0.25113, 
    -0.3150134, -0.332901, -0.2893624, -0.1962961, -0.1261788, -0.07168669, 
    -0.08819059, -0.1226795, -0.2115142, -0.256371, -0.2502511, -0.228897, 
    -0.1568266, -0.06983119, 0.004664242, 0.1075777, 0.1780041, 0.2496838, 
    0.2396903, 0.1321382, 0.1104748, 0.1253348, 0.09312452, 0.09045524, 
    0.09429639, 0.09174105, 0.08422153, 0.05956332, 0.04226188, 0.04455681, 
    0.04483348, 0.05455032, 0.07722279, 0.08374941, 0.08350533, 0.05889595, 
    0.01127231, -0.02585334, -0.06655973, -0.1360421, -0.208487, -0.2942454, 
    -0.3741446, -0.4488839, -0.495759, -0.495824, -0.4811755, -0.4712146, 
    -0.4719633, -0.4538644, -0.425772, -0.4039621, -0.460977, -0.4881906, 
    -0.5325592, -0.5835682, -0.6132557, -0.6058826, -0.5717681, -0.4894113, 
    -0.4418364, -0.3838937, -0.3539296, -0.4147531, -0.3444242, -0.5170479, 
    -0.4663643, -0.4421458, -0.292244, -0.220727, -0.3094635, -0.3811269, 
    -0.4641834, -0.5926341, -0.6879635, -0.6376052, -0.4067621, -0.2485104, 
    -0.1657948, -0.2417549, -0.385977, -0.6094471, -0.7898344, -0.8474028,
  -0.3682036, -0.2349679, -0.007786751, 0.1181084, 0.1972262, 0.2621187, 
    0.2908622, 0.1343192, 0.01727796, -0.1172922, -0.2365629, -0.3080473, 
    -0.3215401, -0.293643, -0.2181385, -0.1305245, -0.05503631, 0.01381135, 
    0.05282503, 0.05116487, 0.03444934, 0.04943961, 0.09491491, 0.1692313, 
    0.222747, 0.3939057, 0.4530366, 0.3677176, 0.3915132, 0.4024995, 
    0.3733166, 0.373463, 0.3608817, 0.3574474, 0.3709565, 0.4022228, 
    0.4265718, 0.4397554, 0.4207124, 0.3878185, 0.3457938, 0.2924572, 
    0.2363537, 0.1682384, 0.09817009, 0.0225516, -0.06183968, -0.1426502, 
    -0.2120675, -0.2629139, -0.3064848, -0.349063, -0.3888416, -0.416283, 
    -0.4378488, -0.4341216, -0.4336333, -0.4117583, -0.3799875, -0.3693917, 
    -0.3637278, -0.3881907, -0.4357167, -0.4857981, -0.5256418, -0.5397206, 
    -0.5419016, -0.5207264, -0.4560129, -0.3697498, -0.2879627, -0.1402739, 
    -0.06141639, -0.00692445, 0.02891552, 0.02510715, 0.008098602, 
    -0.03456092, -0.07572293, -0.1295642, -0.1905668, -0.2982816, -0.4120676, 
    -0.5121163, -0.5874095, -0.5904858, -0.6141353, -0.5900788, -0.5149813, 
    -0.4058995, -0.3164618, -0.3251207, -0.3951732, -0.4787506, -0.4994373, 
    -0.4748279,
  -0.3782297, -0.3109933, -0.2315336, -0.1423897, -0.04800498, 0.03431916, 
    0.1049247, 0.1672944, 0.2261811, 0.2616304, 0.281243, 0.2922293, 
    0.3024994, 0.3136486, 0.3249115, 0.339739, 0.3626231, 0.384905, 
    0.4147066, 0.4583914, 0.5144299, 0.5599377, 0.6052339, 0.6560639, 
    0.7070731, 0.7561452, 0.813616, 0.8472586, 0.8703217, 0.8960053, 
    0.9007254, 0.8872163, 0.8858979, 0.8584728, 0.8321218, 0.7965587, 
    0.7581798, 0.716383, 0.6760184, 0.6379813, 0.5890067, 0.5433686, 
    0.4946382, 0.4372489, 0.3778576, 0.3177828, 0.252288, 0.1781669, 
    0.09909785, 0.02976191, -0.03233123, -0.08254284, -0.1298899, -0.1694406, 
    -0.2015858, -0.2179758, -0.2356679, -0.264981, -0.3017648, -0.3314686, 
    -0.3593821, -0.3771881, -0.4015858, -0.4137115, -0.4041736, -0.3721587, 
    -0.3281645, -0.273591, -0.218464, -0.1665109, -0.1247791, -0.07446986, 
    -0.04886764, -0.03369838, -0.05505255, -0.0861398, -0.1168364, 
    -0.1389556, -0.1221912, -0.0991118, -0.03376365, -0.1082101, -0.1295804, 
    -0.1679919, -0.1136299, -0.0676012, -0.1513089, -0.2084867, -0.2505116, 
    -0.3241607, -0.3784902, -0.4071847, -0.4325592, -0.453604, -0.452839, 
    -0.4298898,
  -0.6230376, -0.5433826, -0.4601307, -0.3649158, -0.2737212, -0.178604, 
    -0.08275443, 0.01293248, 0.1026134, 0.1957774, 0.2803152, 0.3549245, 
    0.4222912, 0.4878022, 0.5497977, 0.6059988, 0.6598887, 0.7046967, 
    0.7397391, 0.7808198, 0.8181896, 0.8543061, 0.89345, 0.9291759, 
    0.9567801, 0.9769461, 0.9886323, 1.002093, 1.011663, 1.017701, 1.005608, 
    1.002744, 0.9910899, 0.960605, 0.9317964, 0.9115328, 0.8749768, 0.822454, 
    0.7843029, 0.7473726, 0.7061941, 0.6574311, 0.6161877, 0.5697359, 
    0.5189221, 0.4690198, 0.4207287, 0.3681898, 0.3130464, 0.258066, 
    0.2037038, 0.1470632, 0.09016216, 0.03514928, -0.01514369, -0.05993539, 
    -0.1101795, -0.1497466, -0.184496, -0.2178619, -0.2500396, -0.2627675, 
    -0.2804433, -0.2957427, -0.3044992, -0.3161203, -0.3131256, -0.3166086, 
    -0.3278879, -0.344994, -0.3616607, -0.3879465, -0.4169341, -0.4494537, 
    -0.486856, -0.529076, -0.5700103, -0.6099843, -0.653718, -0.6969797, 
    -0.7416412, -0.7892811, -0.8324127, -0.8677154, -0.8965729, -0.9185944, 
    -0.9378489, -0.955785, -0.9576731, -0.9479725, -0.9308339, -0.9036855, 
    -0.8638091, -0.8155669, -0.763158, -0.6952544,
  -0.5256057, -0.5305369, -0.5323926, -0.5319043, -0.5290234, -0.5241571, 
    -0.5186558, -0.5117873, -0.504105, -0.4965203, -0.4887569, -0.4819371, 
    -0.4763545, -0.4712272, -0.4688021, -0.4687696, -0.4735875, -0.4819362, 
    -0.4941595, -0.5094752, -0.5262725, -0.5455761, -0.5637238, -0.5800486, 
    -0.5927112, -0.6013377, -0.6039743, -0.5998731, -0.5885937, -0.571373, 
    -0.5472031, -0.5167344, -0.4807, -0.4396355, -0.3951367, -0.3460808, 
    -0.2943883, -0.2410191, -0.1866896, -0.1321161, -0.07790056, -0.02414078, 
    0.02774715, 0.07859349, 0.1281217, 0.1773241, 0.2353969, 0.282696, 
    0.3138158, 0.3240862, 0.3476694, 0.3476045, 0.4245906, 0.494138, 
    0.495163, 0.5070605, 0.5282037, 0.5308731, 0.5063288, 0.5123837, 
    0.4969375, 0.4900854, 0.4868138, 0.4615371, 0.440362, 0.4167125, 
    0.3990202, 0.3735645, 0.3590949, 0.3483202, 0.3328905, 0.315475, 
    0.3009245, 0.193763, 0.234633, 0.2017872, 0.151885, 0.1197236, 
    0.07356405, 0.02792597, -0.02365255, -0.07723379, -0.130815, -0.1807003, 
    -0.2309775, -0.2769408, -0.3184452, -0.3564658, -0.388155, -0.4158731, 
    -0.4400592, -0.4619012, -0.4804235, -0.4965694, -0.5096388, -0.5190623,
  -0.4407261, -0.4203159, -0.3882359, -0.3457554, -0.2985223, -0.2483432, 
    -0.2017287, -0.1608921, -0.1275913, -0.1012892, -0.08143252, -0.06776059, 
    -0.06357765, -0.06616551, -0.07754266, -0.09427434, -0.113057, 
    -0.1317582, -0.1463252, -0.1543328, -0.1598017, -0.1659701, -0.176338, 
    -0.1874218, -0.2004426, -0.2158716, -0.2337596, -0.2515657, -0.2764189, 
    -0.3066761, -0.3327665, -0.3490596, -0.354691, -0.3538938, -0.3461134, 
    -0.3287628, -0.3016796, -0.2654324, -0.2193881, -0.167419, -0.1111851, 
    -0.06357765, -0.0399937, -0.007506847, 0.001705647, -0.0203321, 
    -0.02829051, -0.06512356, -0.09144187, -0.1259634, -0.1179068, 
    -0.1331899, -0.119518, -0.08898425, -0.1106639, -0.03857756, -0.02751017, 
    -0.01263332, 0.004765749, 0.0276823, 0.02664137, 0.01251292, 
    -0.003095627, -0.02571964, -0.04512066, -0.05641618, -0.04941749, 
    -0.0390659, -0.01401711, 0.01988602, 0.06586587, 0.1051887, 0.1271777, 
    0.1579069, 0.1313443, 0.1304002, 0.1103156, 0.08744776, 0.05463523, 
    0.003463149, -0.0154655, -0.0456574, -0.08117175, -0.09889627, 
    -0.1691437, -0.2019398, -0.2577016, -0.3008657, -0.3357453, -0.3637726, 
    -0.3871129, -0.4104521, -0.4276237, -0.4429883, -0.4510776, -0.4512566,
  -0.3804885, -0.4387078, -0.4629754, -0.4615758, -0.4415238, -0.4200394, 
    -0.3866246, -0.3359248, -0.2754105, -0.2163609, -0.1683628, -0.1325718, 
    -0.1025425, -0.07943052, -0.07721698, -0.1031446, -0.1658561, -0.2498245, 
    -0.3312366, -0.3931184, -0.4222529, -0.4170606, -0.3683465, -0.3082879, 
    -0.2829461, -0.2842972, -0.2834834, -0.2733597, -0.2714391, -0.293265, 
    -0.3401725, -0.3996937, -0.459296, -0.5016143, -0.5238967, -0.5337934, 
    -0.5426478, -0.5419798, -0.5186887, -0.4681363, -0.3932662, -0.2797561, 
    -0.1500032, -0.07012033, -0.01351261, -0.01764667, -0.04604835, 
    -0.09290707, -0.1589878, -0.2317417, -0.2976597, -0.3427444, -0.3634312, 
    -0.3661981, -0.3567092, -0.3285842, -0.3094761, -0.3162632, -0.3351761, 
    -0.3740594, -0.424157, -0.4753289, -0.5091995, -0.5082392, -0.4922072, 
    -0.464603, -0.4201043, -0.371976, -0.3150913, -0.2505243, -0.1904656, 
    -0.1401891, -0.1031773, -0.09160507, -0.0914585, -0.09582049, 
    -0.05189148, -0.1331415, -0.158353, -0.1630731, -0.1683789, -0.1609735, 
    -0.1538447, -0.1355828, -0.1019564, -0.04521811, -0.01792312, 
    -0.05675769, -0.06574202, -0.06365848, -0.1110055, -0.1279004, 
    -0.1587434, -0.2101433, -0.2662793, -0.3276564,
  -0.04640603, -0.1181507, -0.2023952, -0.289326, -0.3653677, -0.415612, 
    -0.4533725, -0.4839389, -0.5241407, -0.559948, -0.5680699, -0.550801, 
    -0.4951532, -0.4125522, -0.3327508, -0.2617873, -0.223506, -0.2403031, 
    -0.3292513, -0.4798696, -0.6320512, -0.722904, -0.7110382, -0.6328648, 
    -0.53376, -0.4845413, -0.4724644, -0.4498408, -0.4513871, -0.4661494, 
    -0.4975296, -0.5169307, -0.5135127, -0.5044795, -0.4979364, -0.5072784, 
    -0.5292022, -0.5850296, -0.6615443, -0.7108607, -0.6889362, -0.613627, 
    -0.3825078, -0.1559935, -0.01141262, 0.07024407, 0.05136395, 0.139596, 
    0.1140265, 0.07180646, 0.004065577, -0.1225132, -0.2630894, -0.3726271, 
    -0.4611199, -0.52668, -0.5796908, -0.6832715, -0.631416, -0.5339388, 
    -0.41278, -0.3540883, -0.2654653, -0.224694, -0.1527538, -0.08851171, 
    -0.03146458, 0.01744485, 0.0812633, 0.1336071, 0.1796193, 0.2148087, 
    0.2353973, 0.2483366, 0.2658823, 0.2800421, 0.2527797, 0.2143193, 
    0.169121, 0.1132616, 0.104619, 0.07061831, 0.01568666, -0.01071307, 
    -0.01251966, -0.03454107, -0.05679071, -0.04629242, 0.01365221, 
    -0.002460957, 0.01047873, 0.05487967, 0.07042336, 0.04063821, 0.03661799, 
    0.003968239,
  0.2845831, 0.2837205, 0.2700148, 0.1465611, -0.02482557, -0.1438842, 
    -0.284184, -0.4218788, -0.7010293, -0.7241578, -0.7800975, -0.8146191, 
    -0.8037958, -0.6896193, -0.4708692, -0.2948602, -0.1821161, -0.08558285, 
    -0.04793638, -0.1249707, -0.3583202, -0.6391969, -0.910583, -1.037911, 
    -1.038301, -0.9980175, -0.9648144, -0.8945837, -0.8367221, -0.81265, 
    -0.8026397, -0.7993032, -0.7481153, -0.6570672, -0.5460808, -0.4661982, 
    -0.4607783, -0.5242382, -0.6069695, -0.7055699, -0.7826045, -0.7694697, 
    -0.6337112, -0.4210484, -0.2272007, -0.05449581, 0.08256495, 0.2042608, 
    0.3306769, 0.3388637, 0.2686327, 0.03433901, -0.2226271, -0.4985712, 
    -0.7472039, -0.9646031, -1.203665, -1.344486, -1.380635, -1.27694, 
    -1.102884, -0.9409049, -0.8189646, -0.6993846, -0.5981475, -0.4137561, 
    -0.1703808, -0.06442308, 0.1934869, 0.3670547, 0.3949516, 0.3551238, 
    0.470602, 0.4539844, 0.4301562, 0.5079231, 0.4390914, 0.4241663, 
    0.4164028, 0.3602668, 0.248369, 0.243242, 0.2141242, 0.2000128, 
    0.1907518, 0.1316535, 0.05463529, -0.02005541, -0.06470066, -0.08572924, 
    -0.08913088, -0.1077018, 0.04177809, 0.1056771, 0.1515107, 0.2627573,
  0.09404039, 0.3506968, 0.4144506, 0.4361298, 0.425534, 0.4271128, 
    0.3717256, 0.2362599, 0.2262828, 0.1856089, 0.01228523, -0.09892845, 
    -0.1649456, -0.2073278, -0.2070992, -0.1871119, -0.1532748, -0.105293, 
    -0.1070834, -0.07347333, -0.08416653, -0.08188772, -0.206954, -0.2783084, 
    -0.3586135, -0.3767934, -0.3542676, -0.2976441, -0.2428918, -0.2493529, 
    -0.306921, -0.3549685, -0.326859, -0.2448931, -0.08978224, 0.04276991, 
    0.2131481, 0.3323698, 0.4605274, 0.437269, 0.3499486, 0.1870255, 
    0.09067035, 0.04583001, 0.006702065, 0.1160121, 0.2220667, 0.3281702, 
    0.3932907, 0.419007, 0.3776333, 0.1841112, -0.03778011, -0.2993686, 
    -0.5879755, -0.886771, -1.179252, -1.409492, -1.492256, -1.471716, 
    -1.284688, -1.057263, -0.8221064, -0.6235712, -0.4791374, -0.370739, 
    -0.1879103, -0.04678088, 0.1333298, 0.2638636, 0.3352829, 0.2979945, 
    0.4977177, 0.5758592, 0.6800583, 0.6898402, 0.7041305, 0.74207, 
    0.5262985, 0.5237433, 0.3977831, 0.3561327, 0.369772, 0.4593879, 
    0.5360969, 0.5782355, 0.5648566, 0.4940884, 0.4057746, 0.3397425, 
    0.3092088, 0.2788864, 0.1242318, -0.009134173, -0.1169791, -0.1321323,
  0.7640103, 0.806849, 0.9158659, 1.017071, 1.179067, 1.238377, 1.227943, 
    1.148451, 1.097328, 1.043731, 0.8971651, 0.6464655, 0.319984, 
    -0.01616526, -0.07781935, 0.07187176, 0.1410284, 0.07439494, -0.05317688, 
    -0.2556829, -0.3744497, -0.491442, -0.4107454, -0.2184443, 0.03113317, 
    0.3030894, 0.4712377, 0.5576799, 0.5762019, 0.4714487, 0.3954558, 
    0.3862114, 0.3963504, 0.2342906, 0.328887, 0.290508, -0.2589874, 
    0.1355112, 0.4432745, 0.6489549, 0.7776828, 0.8562632, 0.8042939, 
    0.7319801, 0.6873672, 0.6263962, 0.6451136, 0.7304814, 0.8333298, 
    0.9107387, 0.9556605, 0.9251593, 0.7670376, 0.5958462, 0.4747525, 
    0.3383918, 0.1714973, -0.0254755, -0.2177444, -0.3675491, -0.387715, 
    -0.2178746, 0.126445, 0.4852828, 0.7232062, 0.8005824, 0.7793096, 
    0.7144009, 0.7200812, 0.783102, 0.9296677, 1.164026, 1.467038, 1.732337, 
    1.851982, 1.841028, 1.799638, 1.787643, 1.749769, 1.438864, 1.285186, 
    1.085039, 1.074378, 1.15999, 1.34041, 1.450485, 1.465231, 1.358379, 
    1.196367, 1.081377, 1.004391, 0.9257128, 0.7950487, 0.6878546, 0.669365, 
    0.7009405,
  1.930514, 1.970912, 2.031051, 2.034437, 1.944642, 1.815215, 1.803789, 
    1.938766, 2.144935, 2.248678, 2.291387, 2.303398, 2.262936, 2.162024, 
    2.100175, 2.155352, 2.289727, 2.36375, 2.284811, 2.099329, 1.935722, 
    1.792021, 1.699118, 1.737529, 1.913831, 2.11541, 2.250615, 2.277373, 
    2.173092, 1.996709, 1.798939, 1.663538, 1.703366, 1.835072, 1.904619, 
    1.91292, 1.848466, 1.792591, 1.693047, 1.557809, 1.50374, 1.51943, 
    1.562464, 1.537708, 1.480547, 1.472295, 1.499752, 1.556556, 1.685039, 
    1.825892, 1.929603, 2.008883, 2.093503, 2.149166, 2.136162, 2.035609, 
    1.826787, 1.611129, 1.388083, 1.115036, 0.8796189, 0.7559371, 0.8417933, 
    1.076168, 1.327861, 1.476445, 1.445488, 1.319886, 1.227617, 1.254082, 
    1.340996, 1.393438, 1.498955, 1.680873, 1.849476, 1.988929, 2.089726, 
    2.233753, 2.387383, 2.490849, 2.490182, 2.342086, 2.135478, 2.003349, 
    1.911878, 1.880124, 1.852698, 1.825062, 1.75055, 1.700029, 1.797441, 
    1.948678, 1.994788, 1.990361, 1.961097, 1.937383,
  2.379733, 2.23097, 2.197734, 2.252796, 2.285397, 2.219316, 2.149606, 
    2.154993, 2.241875, 2.354878, 2.496789, 2.685006, 2.926331, 3.120244, 
    3.188033, 3.224378, 3.356018, 3.513586, 3.612333, 3.680449, 3.724459, 
    3.700012, 3.616467, 3.520064, 3.416484, 3.320325, 3.243306, 3.205872, 
    3.030936, 2.786308, 2.550142, 2.394592, 2.327356, 2.346188, 2.378056, 
    2.514482, 2.789303, 3.012056, 3.040654, 2.869885, 2.684973, 2.612398, 
    2.501071, 2.333899, 2.224036, 2.247034, 2.380221, 2.505319, 2.631946, 
    2.819626, 3.072441, 3.290117, 3.436194, 3.50911, 3.502926, 3.368454, 
    3.221627, 3.146123, 3.054505, 2.860836, 2.586292, 2.361634, 2.216614, 
    2.160233, 2.155188, 2.149085, 2.116321, 2.048564, 1.96689, 1.871106, 
    1.843518, 1.819056, 1.727291, 1.690475, 1.849476, 2.166142, 2.353138, 
    2.330692, 2.362838, 2.531246, 2.648319, 2.554049, 2.419543, 2.327633, 
    2.291142, 2.349182, 2.478398, 2.59941, 2.618665, 2.679309, 2.785478, 
    2.850582, 2.85037, 2.758931, 2.657808, 2.534094,
  2.474248, 2.41821, 2.404375, 2.465996, 2.530401, 2.547377, 2.479018, 
    2.415004, 2.454929, 2.522573, 2.529701, 2.446742, 2.466045, 2.623028, 
    2.844268, 2.941761, 3.001771, 3.114923, 3.208022, 3.231345, 3.326918, 
    3.386716, 3.375144, 3.342266, 3.245391, 3.134438, 3.119577, 3.202943, 
    3.146124, 2.946677, 2.715574, 2.548777, 2.394578, 2.194105, 2.001446, 
    1.881654, 1.967543, 2.232289, 2.483315, 2.653741, 2.704067, 2.711667, 
    2.745782, 2.814207, 2.861765, 2.86323, 2.924769, 3.052486, 3.236096, 
    3.414807, 3.530416, 3.59425, 3.546139, 3.485282, 3.445601, 3.4144, 
    3.36396, 3.389156, 3.420991, 3.31829, 3.128365, 2.996041, 2.865589, 
    2.736911, 2.637968, 2.481946, 2.339336, 2.249557, 2.138913, 1.986438, 
    1.943568, 2.03211, 2.005027, 1.878318, 1.866778, 1.924997, 1.837644, 
    1.63569, 1.555758, 1.654749, 1.874135, 1.957028, 1.931214, 1.975501, 
    2.155644, 2.322034, 2.432809, 2.53927, 2.601233, 2.634274, 2.739776, 
    2.903708, 2.966648, 2.897946, 2.756084, 2.594984,
  2.165394, 2.1749, 2.172978, 2.088978, 1.902162, 1.763327, 1.689906, 
    1.59596, 1.500485, 1.479001, 1.482614, 1.408574, 1.318584, 1.30654, 
    1.366061, 1.435608, 1.53494, 1.622961, 1.638814, 1.690084, 1.873905, 
    1.994917, 1.962317, 1.962332, 1.986081, 1.985381, 1.994967, 2.068047, 
    2.172979, 2.195976, 2.106686, 1.903284, 1.735168, 1.669429, 1.674411, 
    1.689434, 1.715508, 1.742835, 1.807208, 1.92721, 2.044951, 2.065834, 
    2.069121, 2.174818, 2.278285, 2.263181, 2.24238, 2.395131, 2.630873, 
    2.832468, 2.960382, 3.115086, 3.215639, 3.164597, 3.106263, 3.035658, 
    2.914809, 2.892282, 2.966925, 2.979766, 2.941713, 2.855011, 2.619105, 
    2.389092, 2.304457, 2.212172, 2.071172, 1.943584, 1.797621, 1.563897, 
    1.439743, 1.46699, 1.41471, 1.329098, 1.23434, 1.048369, 0.8913536, 
    1.018226, 1.125518, 1.067087, 0.9960909, 0.9741664, 0.9258265, 0.9146614, 
    1.047897, 1.246286, 1.431166, 1.508574, 1.456768, 1.488278, 1.635592, 
    1.839808, 2.035853, 2.135202, 2.146351, 2.136276,
  1.06782, 0.9833775, 0.9477825, 0.9607058, 0.9391069, 0.8841753, 0.8247347, 
    0.7067175, 0.526721, 0.3245249, 0.1678348, 0.0939579, 0.02634716, 
    -0.08063507, -0.1108599, -0.01497746, 0.2145967, 0.410511, 0.4498177, 
    0.5413857, 0.7311974, 0.7915659, 0.7149553, 0.7002087, 0.7513313, 
    0.8185358, 0.8712378, 0.8333302, 0.8131151, 0.8970022, 0.958086, 
    0.8304176, 0.6269178, 0.4925423, 0.3778448, 0.3444633, 0.4341278, 
    0.4993944, 0.4524374, 0.4124641, 0.5042276, 0.611455, 0.6055951, 
    0.5834107, 0.6877732, 0.8041148, 0.7525845, 0.675127, 0.8743944, 
    1.279261, 1.604978, 1.944008, 2.26266, 2.423125, 2.535105, 2.634404, 
    2.595651, 2.541582, 2.482289, 2.308444, 2.131588, 1.983591, 1.721725, 
    1.462318, 1.344935, 1.273793, 1.191419, 1.129895, 1.015263, 0.82301, 
    0.7437778, 0.7111773, 0.5663214, 0.4933558, 0.4104466, 0.1249795, 
    -0.03719425, 0.03720284, -0.1416869, -0.4477262, -0.3394418, -0.144259, 
    -0.1661334, -0.2492228, -0.2567587, -0.2145386, -0.1023955, 0.03336287, 
    0.1588674, 0.3186979, 0.519496, 0.6995411, 0.8616347, 1.023565, 1.115214, 
    1.118356,
  -0.0595417, -0.05711746, -0.1242867, -0.1905956, -0.2165403, -0.1770544, 
    -0.1397986, -0.2608104, -0.3854699, -0.4749064, -0.6297402, -0.7556353, 
    -0.844161, -0.8632851, -0.8117065, -0.789392, -0.7442594, -0.5931678, 
    -0.4617548, -0.3779173, -0.3025265, -0.3748245, -0.3916054, -0.2845078, 
    -0.2487011, -0.2344589, -0.1726599, -0.1832056, -0.2573767, -0.3037949, 
    -0.2685909, -0.2886267, -0.382165, -0.4670448, -0.5610061, -0.6160846, 
    -0.7207232, -0.8929892, -0.8715696, -0.8384967, -0.9125528, -0.8877153, 
    -0.7285519, -0.6642289, -0.6866412, -0.6001501, -0.4564338, -0.5171103, 
    -0.4335976, -0.03626728, 0.2888465, 0.552927, 0.9455209, 1.218096, 
    1.414417, 1.616745, 1.629652, 1.553854, 1.431198, 1.209909, 1.062644, 
    0.9330049, 0.8162241, 0.7625623, 0.6243296, 0.4702606, 0.3637176, 
    0.1845021, 0.0860157, -0.03717756, -0.1929393, -0.2798052, -0.3636746, 
    -0.4498901, -0.6212931, -0.7529993, -0.573132, -0.520088, -1.046243, 
    -1.334166, -0.8747747, -0.6063995, -0.6628613, -0.6941767, -0.8052607, 
    -0.9226928, -0.95575, -0.9347215, -0.8785362, -0.812048, -0.7335315, 
    -0.5910997, -0.4026723, -0.2479362, -0.1544313, -0.1002159,
  -0.9864945, -0.9315958, -0.8852253, -0.911983, -1.086316, -1.208988, 
    -1.076957, -0.9689975, -0.9962759, -1.018558, -1.026891, -1.006237, 
    -1.086527, -1.21553, -1.276338, -1.413073, -1.591116, -1.595315, 
    -1.54403, -1.501631, -1.369568, -1.335193, -1.389034, -1.409575, 
    -1.365744, -1.261446, -1.277625, -1.365108, -1.443543, -1.619763, 
    -1.719714, -1.685404, -1.580146, -1.44001, -1.468427, -1.549157, 
    -1.684866, -1.80788, -1.616637, -1.415042, -1.547333, -1.54206, 
    -1.557816, -1.696081, -1.831547, -1.916101, -1.73464, -1.551549, 
    -1.581644, -1.394584, -1.102185, -0.8225298, -0.3381062, 0.07382441, 
    0.3060179, 0.4790163, 0.4342246, 0.2916141, 0.09403849, -0.1218467, 
    -0.07249832, -0.101388, -0.1854377, -0.1999717, -0.367208, -0.4748416, 
    -0.5679898, -0.7931523, -0.8925829, -0.9456749, -1.049516, -1.198751, 
    -1.341378, -1.347595, -1.438887, -1.471243, -0.9079949, -0.5461459, 
    -0.9157751, -0.8693069, -0.3975458, -0.3905958, -0.4853714, -0.6799188, 
    -1.068086, -1.221357, -1.271991, -1.347561, -1.429935, -1.491686, 
    -1.515889, -1.447026, -1.37131, -1.310584, -1.177966, -1.051795,
  -1.895657, -1.780146, -1.675996, -1.604642, -1.652396, -1.800378, 
    -1.772497, -1.476843, -0.9892613, -0.865254, -1.046895, -1.31042, 
    -1.613041, -1.838594, -1.911071, -1.915677, -2.00072, -2.009818, 
    -1.902071, -1.977494, -2.111722, -2.094681, -2.115612, -2.160224, 
    -2.163561, -2.081204, -2.115009, -2.150329, -2.12611, -2.342761, 
    -2.507507, -2.518346, -2.373571, -1.873717, -1.759964, -1.824157, 
    -1.517891, -1.027722, -0.79224, -1.074108, -1.164375, -1.110615, 
    -1.452917, -1.879968, -2.016735, -2.176582, -2.36195, -2.309134, 
    -2.171845, -1.9064, -1.600606, -1.508662, -1.287796, -0.9708366, 
    -0.8494499, -0.7519403, -0.7071478, -0.5889673, -0.5605981, -0.7225285, 
    -0.6639998, -0.6498888, -0.8095891, -0.9116886, -1.068395, -1.118069, 
    -1.092239, -1.187682, -1.315123, -1.505195, -1.533776, -1.53485, 
    -1.69849, -1.599467, -1.300573, -0.867484, -0.2005405, -0.01562858, 
    -0.5596063, -0.6219268, -0.145918, -0.2457716, -0.214668, -0.3533725, 
    -0.7165236, -0.8495152, -1.188122, -1.483662, -1.698148, -1.789489, 
    -1.746162, -1.769404, -1.794567, -1.8494, -1.862063, -1.886819,
  -2.048229, -1.884622, -1.699824, -1.430667, -0.8569856, -0.5604852, 
    -0.5806509, -0.5708203, -0.2958692, -0.2296095, -0.6266308, -1.112487, 
    -1.421927, -1.380082, -1.227413, -1.248376, -1.47961, -1.791117, 
    -1.818021, -1.822692, -1.987113, -2.119421, -2.221862, -2.194176, 
    -2.207165, -2.157816, -2.105147, -2.106547, -1.908175, -1.717273, 
    -1.293363, -1.120967, -1.197351, -0.967044, -0.777819, -0.6359408, 
    -0.6571486, -0.5504428, -0.4825068, -0.9071975, -1.118574, -1.115042, 
    -1.2939, -1.316768, -1.301989, -1.484411, -1.788643, -1.815286, 
    -1.727461, -1.851745, -1.950377, -2.023376, -1.979349, -1.779072, 
    -1.702754, -1.564896, -1.307604, -0.9920119, -0.6808791, -0.6409865, 
    -0.7321324, -0.83223, -1.01916, -1.099401, -1.20793, -1.30959, -1.306823, 
    -1.3446, -1.364424, -1.465612, -1.418867, -1.324808, -1.246113, 
    -1.115156, -0.8694042, -0.2464715, 0.2992315, 0.4645475, -0.2058628, 
    -0.5758493, -0.2691605, -0.2573602, -0.113317, 0.05258441, -0.08966708, 
    -0.3073602, -0.7634636, -0.8729525, -1.062406, -1.376322, -1.525557, 
    -1.781628, -1.909476, -2.008939, -2.119047, -2.131416,
  -1.409574, -1.243558, -0.9083042, -0.4336305, 0.02074862, 0.09477195, 
    -0.04101906, -0.1069371, -0.1569693, -0.1339712, -0.01623058, -0.2922082, 
    -0.7656775, -0.7633824, -0.3385782, -0.3341346, -0.8515177, -1.262796, 
    -1.31763, -1.155457, -1.029593, -1.0481, -1.340417, -1.493428, -1.501729, 
    -1.396846, -1.127331, -0.9539261, -0.6505575, -0.3758664, -0.06990862, 
    -0.209883, -0.5398469, -0.5573599, -0.5819855, -0.3237822, -0.2502639, 
    -0.4066602, -0.5377145, -0.7827667, -0.7444696, -0.8639848, -0.9230995, 
    -0.5626335, -0.3898311, -0.3593946, -0.5694375, -0.7465534, -0.7215538, 
    -1.046537, -1.434134, -1.700361, -1.87043, -1.77196, -1.681987, 
    -1.531839, -1.206645, -1.109899, -1.059411, -1.027543, -1.057686, 
    -1.014034, -1.079593, -1.115466, -1.150459, -1.205065, -1.154968, 
    -1.21213, -1.102233, -0.9539585, -0.8669796, -0.7501495, -0.5242712, 
    -0.3539908, -0.155781, 0.148597, -0.07746112, 0.3699673, 0.1535934, 
    -0.5765007, -0.148799, 0.046839, 0.03448558, 0.3128711, 0.356931, 
    0.2207489, -0.06150961, -0.1992223, -0.4897492, -0.8755401, -1.164993, 
    -1.410762, -1.52878, -1.58721, -1.567549, -1.469471,
  -0.4538293, -0.2386756, -0.02923536, 0.2576628, 0.3809697, 0.1477832, 
    -0.1077182, -0.032897, -0.01740217, 0.09784842, 0.5164845, 0.4091766, 
    -0.1883988, -0.7145867, -0.3370476, -0.04310369, -0.7160034, -1.101159, 
    -0.8861847, -0.5362983, -0.502233, -0.4096222, -0.441165, -0.5824084, 
    -0.5763702, -0.5863314, -0.3164921, 0.009566307, 0.3547482, 0.642086, 
    0.827845, 0.3565885, -0.2765336, -0.1703322, -0.2435257, -0.2540078, 
    -0.1192412, -0.06850886, -0.2714059, -0.4408071, -0.2486525, -0.3569217, 
    -0.4467807, -0.2437377, 0.1443806, 0.4453077, 0.1832638, -0.07755899, 
    -0.02327871, -0.09359121, -0.4674354, -1.083272, -1.536609, -1.467614, 
    -1.320788, -1.436934, -1.418331, -1.316264, -1.339083, -1.27476, 
    -1.119682, -0.923214, -0.9325886, -0.9819703, -0.93573, -0.9450235, 
    -0.8549194, -0.800817, -0.5757689, -0.4951859, -0.4022012, -0.1716838, 
    -0.08784628, 0.07086229, 0.3345509, 0.3706834, -0.3580926, 0.1436813, 
    0.3093879, -0.8123572, -0.2147495, 0.1127734, -0.07671261, -0.03069997, 
    0.001168728, 0.149997, 0.08980823, -0.1559436, -0.344372, -0.5078485, 
    -0.7615106, -0.7425337, -0.8032756, -0.7697959, -0.6989293, -0.6595087,
  0.1966758, 0.2220831, 0.2579393, 0.4800909, 0.5293423, 0.1889941, 
    0.1369435, 0.1180308, -0.05106115, 0.1108365, 0.3712695, 0.312578, 
    0.08145815, -0.4900751, -0.6307163, 0.06540966, -0.2144408, -0.9403682, 
    -0.929121, -0.2774782, 0.05994177, 0.08236885, 0.03406286, -0.02664757, 
    0.1574502, 0.2425575, 0.4724073, 0.7416306, 0.7764454, 0.7769992, 
    1.145765, 1.327861, 0.7430143, 0.2701631, 0.08057952, -0.02386308, 
    -0.05062151, 0.02952123, -0.2821808, -0.3454304, -0.09647226, 0.07751846, 
    0.2593222, 0.2329712, 0.6914186, 1.026266, 0.6827273, 0.542851, 
    0.7301397, 0.9000931, 0.6250443, -0.1461792, -0.8825231, -1.213122, 
    -1.208776, -1.273116, -1.368184, -1.307621, -1.287943, -1.180081, 
    -1.073783, -0.9438353, -0.804822, -0.7771039, -0.6677289, -0.6310902, 
    -0.567028, -0.5113802, -0.3257189, -0.2187204, -0.1573763, -0.001208782, 
    0.1210403, 0.3804655, 0.3815236, 0.3131638, 0.01876283, 0.2438447, 
    0.1741665, -0.3674188, -0.40098, -0.2025912, -0.07176447, -0.1495804, 
    -0.1416862, -0.327575, -0.1580765, -0.07744455, -0.1287632, -0.07632256, 
    -0.2352414, -0.2382693, -0.3117228, -0.20544, -0.05913496, 0.05465031,
  0.3253224, 0.2837858, 0.1331021, 0.3197396, 0.2253222, -0.2028519, 
    0.005611658, 0.1150846, -0.06985974, 0.1728808, 0.2805305, 0.1836554, 
    0.02665651, -0.1616245, -0.5298047, -0.01761436, 0.1138964, -0.6351104, 
    -0.9291377, -0.536885, -0.05762148, 0.1658821, 0.3035607, 0.3907518, 
    0.5662236, 0.6017387, 0.5958798, 0.7753874, 0.9032517, 0.7495571, 
    0.7429002, 1.188718, 1.412676, 0.9070603, 0.6004034, 0.373906, 0.4101689, 
    0.6442836, 0.4600391, 0.4894333, 0.481637, 0.8200822, 1.234275, 1.092429, 
    1.113962, 1.398907, 0.9950814, 0.3765106, 0.3295867, 0.7914357, 
    0.9142714, 0.445456, -0.1998248, -0.6801147, -0.958858, -1.120577, 
    -1.186983, -1.154203, -1.120967, -1.080423, -1.028373, -0.8791695, 
    -0.6707387, -0.5581408, -0.4631705, -0.4160185, -0.3038278, -0.2190299, 
    -0.2365427, -0.1030145, -0.03660917, 0.1081662, 0.2237101, 0.1950159, 
    0.09578133, 0.2705532, 0.3663051, 0.2249806, 0.04571599, 0.002844691, 
    -0.2742385, -0.3441115, -0.1566441, -0.01055026, 0.2309211, -0.3875525, 
    -0.3476758, -0.009378433, -0.08192158, 0.1734004, 0.2373815, 0.2156043, 
    0.2618608, 0.2726192, 0.2466269, 0.3045535,
  0.1789029, 0.1583624, -0.1617059, -0.06149435, 0.14028, -0.06938821, 
    0.01527977, 0.06425434, -0.0003452301, 0.1225225, 0.07638007, 
    -0.02594745, -0.2099482, -0.1378942, -0.3095739, -0.1715205, 0.009387851, 
    -0.4575392, -0.7800002, -0.6880567, -0.2020541, 0.06047857, 0.1485156, 
    0.2201953, 0.3447717, 0.5308886, 0.494593, 0.51069, 0.672051, 0.7840295, 
    0.7412727, 0.6137495, 0.8750942, 1.052991, 1.08997, 0.756279, 0.9225065, 
    1.263815, 1.06279, 1.290963, 1.239873, 1.397702, 1.296628, 1.23818, 
    0.9010708, 0.901201, 0.8495083, 0.09980124, -0.4855337, -0.3654981, 
    0.2142057, 0.2152314, -0.2431183, -0.4963572, -0.6235385, -0.7930703, 
    -0.7749715, -0.7031941, -0.6391635, -0.6392293, -0.6538277, -0.5801625, 
    -0.4768586, -0.242744, -0.05197239, 0.006930351, -0.05229807, 0.04506397, 
    0.04975176, 0.05235577, 0.03149033, 0.09825468, 0.08280945, -0.03493166, 
    0.0171515, 0.1088182, 0.1714484, 0.0835415, -0.002851725, 0.001103342, 
    -0.08330421, -0.1688836, -0.2655471, -0.2127311, 0.1091113, -0.2469273, 
    -0.5028844, -0.1324415, 0.06282187, 0.216012, 0.3287563, 0.3251915, 
    0.3029909, 0.2822881, 0.2500458, 0.2236791,
  0.1557258, 0.03940088, -0.04635739, 0.009599686, 0.09119177, 0.1309863, 
    0.1192349, 0.2473598, 0.3575649, 0.4036424, 0.3095505, 0.2098435, 
    -0.1117873, -0.1179723, -0.1153352, -0.0951364, 0.1474903, -0.1584506, 
    -0.5504755, -0.4951532, -0.07348979, 0.01062483, -0.04342806, 0.1190884, 
    0.09561837, 0.2433071, 0.3222623, 0.2468884, 0.1735482, 0.05815125, 
    0.1483688, 0.22721, 0.4403939, 0.3369925, 0.5074177, 0.5685835, 1.135819, 
    0.8711872, 0.2476201, 0.4492642, 0.7586228, 0.9986621, 0.3816373, 
    0.2785774, -0.1632522, -0.4283399, -0.08983082, -0.1194859, -0.5655634, 
    -0.8840526, -0.4105179, -0.2059114, -0.374352, -0.4377964, -0.4333203, 
    -0.4648471, -0.4017615, -0.2959018, -0.1972213, -0.06497812, -0.08242607, 
    -0.1305218, -0.07272577, 0.1558557, 0.1970663, 0.2625933, 0.2186971, 
    0.1748166, 0.1393352, 0.1044884, 0.1529756, 0.07693386, -0.06575847, 
    -0.1388707, -0.09027036, 0.02318978, 0.02909812, -0.01846045, 
    -0.01214536, -0.06292662, -0.125801, -0.1486525, -0.1974156, -0.5505405, 
    -0.3895704, 0.05234039, -0.3122106, -0.2693884, 0.01391292, 0.07913089, 
    0.2659476, 0.3128388, 0.3389618, 0.4256647, 0.2869271, 0.2207646,
  0.4126431, 0.2411097, 0.1645801, 0.1748667, 0.3865368, 0.219121, 
    0.09599268, 0.2189907, 0.3389776, 0.6402635, 0.9893682, 0.5685353, 
    -0.01911116, -0.02112974, -0.06886721, -0.1363806, -0.03167653, 
    -0.1275586, -0.2873405, -0.3681347, -0.215726, -0.1940463, -0.3038282, 
    -0.1780467, -0.2752142, -0.2664256, -0.2120957, -0.2995791, -0.09344411, 
    -0.04417634, -0.1974316, -0.1984246, 0.2683234, 0.1708138, 0.2346482, 
    0.2748668, 0.1916955, -0.1073441, -0.06906268, 0.06584944, -0.006350994, 
    0.04006815, -0.5599481, -0.6529819, -0.9600457, -1.259671, -1.080277, 
    -0.8768586, -0.9461621, -1.049336, -0.7861362, -0.7245147, -0.6077185, 
    -0.4130082, -0.2376983, -0.07796526, 0.02291369, 0.2533174, 0.3659313, 
    0.4621062, 0.5744433, 0.6001761, 0.5814097, 0.6852348, 0.7238903, 
    0.6424937, 0.5176239, 0.3853159, 0.4005344, 0.254571, 0.1595507, 
    0.1235641, 0.08302051, -0.02026707, -0.1689162, 0.1364387, 0.1596157, 
    0.0400519, -0.0009474456, 0.004065573, 0.009876132, -0.07884455, 
    -0.02505225, -0.2821649, -0.4673861, -0.05986655, -0.2962761, -0.2951858, 
    -0.06728852, 0.0712204, 0.1455693, 0.2521123, 0.3872523, 0.4523402, 
    0.3602179, 0.3855597,
  0.1144009, 0.1897755, 0.1242483, 0.1398402, 0.213587, 0.08220679, 
    0.006865054, -0.0119175, 0.09949201, 0.6299769, 1.148597, 0.3105767, 
    -0.006807804, 0.2153945, 0.1636847, 0.1137985, -0.07736346, -0.2121617, 
    -0.1923374, -0.1585158, -0.03574562, 0.008248508, -0.2366408, -0.2788122, 
    -0.2323114, -0.2834505, -0.3438674, -0.07458025, -0.04604836, -0.1275749, 
    -0.04230487, -0.127689, -0.03361347, 0.08510399, 0.2563768, 0.0988898, 
    -0.06665382, -0.1157424, -0.08597349, -0.01046896, -0.3016473, 
    -0.4457389, -0.7799183, -0.8978219, -1.09696, -1.158695, -1.101957, 
    -1.058939, -1.123994, -1.031742, -0.8471885, -0.8662477, -0.7786174, 
    -0.5697632, -0.3632851, -0.1884317, -0.09482813, 0.07597303, 0.2372036, 
    0.3708463, 0.5939741, 0.7992318, 0.9616995, 1.067852, 1.09972, 1.014499, 
    0.9618454, 0.7306768, 0.7018845, 0.4792121, 0.1929327, 0.09498352, 
    -0.03753614, -0.006643891, -0.13778, 0.06571937, 0.2390265, 0.1631802, 
    0.01122704, 0.0147264, 0.1215135, -0.08050454, -0.0305537, -0.1854203, 
    -0.3069692, -0.2971385, -0.2939808, -0.1597037, -0.0818069, -0.01165718, 
    -0.07711932, 0.1238247, 0.1501756, 0.1444952, 0.1573207, 0.1255827,
  -0.2373729, -0.03428102, 0.1659639, 0.1461719, 0.09114236, 0.05273092, 
    0.01804671, -0.07135761, 0.1277472, 0.7042607, 1.071058, 0.2673633, 
    0.09700155, 0.2658, 0.3540502, 0.3526831, 0.2238252, 0.1488252, 
    0.08489251, 0.08889627, 0.0245409, -0.0194695, -0.04744804, -0.09505552, 
    -0.1293328, -0.141719, -0.2380244, -0.1062047, -0.1599642, -0.3677118, 
    -0.1051792, 0.003007635, 0.06907213, 0.2179825, 0.3776989, 0.2532687, 
    0.1822562, 0.1084285, -0.09655261, -0.1683786, -0.1931677, -0.2598014, 
    -0.2924032, -0.3991899, -0.535388, -0.4065304, -0.3159547, -0.2362995, 
    -0.3324423, -0.2776737, -0.2652383, -0.2527709, -0.2378783, -0.2421103, 
    -0.2939982, -0.3217978, -0.2460489, -0.2011108, -0.07518291, 0.0472126, 
    0.270927, 0.4213505, 0.6177535, 0.7261527, 0.7930958, 0.8674943, 
    0.9493462, 0.8169401, 0.8151984, 0.7169237, 0.5133592, 0.3409796, 
    0.0002408028, -0.09360647, -0.4390979, -0.1019565, 0.2891242, 0.30457, 
    0.1579393, 0.08717102, -0.05737638, -0.05989927, -0.3320508, -0.2359581, 
    -0.2123899, -0.0231328, 0.1119428, 0.150192, 0.1473119, 0.1385218, 
    0.03306948, 0.01975566, -0.02262723, 0.1369758, -0.08742166, -0.2464387,
  -0.1117873, -0.181986, 0.03500617, -0.1835321, -0.02495462, 0.03458316, 
    -0.1469598, -0.1742548, 0.1329067, 0.4287564, 0.4752895, 0.4871881, 
    0.2478647, 0.2144341, 0.5044885, 0.4192834, 0.2784142, 0.1596324, 
    0.1469696, 0.1415496, 0.01658201, -0.007359743, 0.03201175, -0.1232617, 
    -0.2648959, -0.1787144, -0.09420916, -0.1949741, -0.4270549, -0.3117542, 
    -0.1487174, 0.06757486, 0.266875, 0.1580853, 0.2152963, 0.2773566, 
    0.1941524, 0.1659784, 0.1760697, 0.1733193, 0.01832247, -0.1510134, 
    -0.1295114, -0.2213569, -0.2586617, -0.1675487, -0.1656938, -0.1656122, 
    -0.1979036, -0.1176143, -0.06544924, -0.002151966, 0.05377245, 
    -0.05535841, -0.1185417, -0.1798048, -0.2639842, -0.3263216, -0.3120155, 
    -0.3796587, -0.2385945, -0.07264423, 0.07102489, 0.1436319, 0.3006635, 
    0.5093389, 0.6771779, 0.7817028, 0.7943497, 0.6817682, 0.4959443, 
    0.5533496, 0.5034959, 0.1615525, -0.1597364, 0.0836066, 0.7419887, 
    0.2060677, 0.2583463, -0.09912443, -0.2875519, -0.2923045, -0.2266307, 
    -0.1490922, 0.008623123, 0.1984339, 0.2102332, 0.2813268, 0.326282, 
    0.378366, 0.3116502, 0.1944627, 0.1258266, 0.1880667, 0.04250956, 
    -0.04656917,
  -0.1032749, -0.1617222, -0.3675489, -0.4151564, 0.03972626, 0.02361315, 
    -0.1190462, -0.01722336, 0.3468879, 0.5591599, 0.2496058, 0.2291143, 
    0.1355276, 0.01274014, 0.3665166, 0.5102334, 0.4638309, 0.3621874, 
    0.4085097, 0.3086227, 0.3507941, -0.03908181, -0.1998572, -0.2848182, 
    -0.6654663, -0.8460331, -0.5699253, -0.2496774, -0.5367055, -0.3855991, 
    -0.04844093, -0.1440463, 0.003105164, 0.04931378, 0.06300116, 0.1317992, 
    0.128952, 0.09443045, 0.1119919, 0.008410931, -0.07816124, -0.03810596, 
    -0.05356789, -0.1230831, -0.122448, -0.161315, -0.08122063, -0.01015949, 
    0.02493191, -0.02881145, 0.0246706, 0.0294075, 0.09539032, 0.05832958, 
    0.02607059, 0.01723289, -0.07419014, -0.1798048, -0.1948113, -0.1865759, 
    -0.1405144, -0.08050442, -0.02173185, -0.01264954, -0.05179453, 
    0.1494751, 0.3906536, 0.6634898, 0.8280725, 0.8553839, 0.8057423, 
    0.9783978, 0.8042598, 0.07755184, 0.07122052, 0.3900682, 0.3399705, 
    -0.02739549, -0.06369162, -0.3486371, -0.3553419, -0.1979856, -0.2361031, 
    0.0681119, 0.1293907, 0.2121387, 0.2645469, 0.3833456, 0.4590774, 
    0.5951138, 0.5741346, 0.6825324, 0.5373827, 0.2282355, -0.00386095, 
    -0.01261759,
  -0.3150909, -0.3545601, -0.4586458, -0.4084501, -0.2384639, -0.2302766, 
    -0.02497101, 0.2039356, 0.5239874, 0.700371, 0.2906051, -0.1412145, 
    -0.1499059, 0.03126335, 0.1872845, 0.4612584, 0.5212364, 0.6373343, 
    0.5531867, 0.3809209, 0.4403937, -0.2675974, -0.2934763, -0.38765, 
    -0.7665236, -0.7330923, -0.7120639, -0.2605502, -0.4582551, -0.2198114, 
    0.2050095, -0.1700392, -0.3375854, -0.1551466, -0.3264189, -0.434834, 
    -0.4341502, -0.3818717, -0.3026719, -0.2668653, -0.1945996, -0.1537638, 
    -0.07038116, -0.04072571, 0.01938152, 0.01689148, 0.0955534, 0.03269482, 
    0.1429815, 0.1043434, 0.1359339, 0.119626, 0.04356766, 0.003333092, 
    0.0373497, 0.1511354, 0.1157675, -0.01372433, -0.04420948, 0.03448486, 
    0.1037073, 0.1527309, 0.1439748, 0.1949677, 0.2224402, 0.3048301, 
    0.2171843, 0.5032516, 0.9952278, 1.272083, 1.427471, 1.245489, 0.600502, 
    0.09678984, 0.6241336, 0.6477346, 0.329277, 0.2720184, 0.01418877, 
    -0.30163, -0.3273954, -0.2389522, -0.1070185, -0.003535271, 0.06077099, 
    0.2753544, 0.3274865, 0.4604125, 0.5299926, 0.6794877, 0.6481247, 
    0.6486132, 0.3128221, -0.00120759, -0.003094912, -0.1287632,
  -0.5164092, -0.5719922, -0.4584017, -0.3703969, -0.4578483, -0.481205, 
    -0.1506219, 0.1838672, 0.5158982, 0.5540492, 0.4164842, -0.2248082, 
    -0.3998079, 0.1623828, 0.2468066, 0.2394989, 0.2524705, 0.6991179, 
    0.7175102, 0.6427698, 0.4441535, -0.4531124, -0.3074741, -0.2896681, 
    -0.2026076, -0.2329952, -0.5580763, -0.7423209, -0.5359735, -0.1232452, 
    -0.3157752, -0.7149286, -0.8257198, -0.8365107, -0.9938507, -0.8798208, 
    -0.8292508, -0.7476268, -0.7257681, -0.7403188, -0.6113963, -0.5005889, 
    -0.2489285, -0.2793813, -0.1827669, -0.05818987, 0.0943327, 0.02177334, 
    0.09937859, 0.1080213, 0.1032033, 0.1809049, 0.1673636, 0.1458468, 
    0.183672, 0.2270803, 0.1422324, 0.1157675, 0.1610479, 0.06933212, 
    -0.06341505, 0.01995087, 0.02830124, 0.1105113, 0.2096143, 0.1496873, 
    0.1008267, 0.3379523, 0.3181932, 0.1524543, 0.2005662, -0.01234078, 
    -0.06300807, 0.5662079, 0.9823036, 0.7770467, 0.4859018, 0.1661911, 
    -0.1823435, -0.07410812, -0.05244541, -0.1499705, -0.1188507, 
    -0.09162235, 0.1234012, 0.2919884, 0.3471642, 0.5008097, 0.4491334, 
    0.4626417, 0.4636836, 0.3682425, -0.0315299, -0.1397986, -0.2554393, 
    -0.3662791,
  -0.3172724, -0.6032751, -0.7296584, -0.5320017, -0.6150916, -0.6461129, 
    -0.4148467, -0.196846, 0.1265264, 0.2288864, 0.389694, -0.116068, 
    -0.5744333, -0.003209949, 0.3253546, 0.008346081, -0.1098175, 0.39054, 
    0.4047978, 0.4087366, -0.08146507, -0.4343459, -0.2760937, -0.3239455, 
    -0.3959017, -0.21654, -0.2748244, -0.3773797, -0.3996454, -0.1050816, 
    -0.6842811, -1.384509, -1.686869, -1.516377, -1.454936, -1.383435, 
    -1.358761, -1.247775, -1.059981, -0.8965535, -0.6363316, -0.5630412, 
    -0.4799685, -0.4439492, -0.2526083, -0.210144, -0.1115437, -0.03380966, 
    0.03865194, 0.08342648, 0.03962851, 0.0001101494, -0.06621504, 
    -0.1181679, -0.07555676, 0.02330303, 0.1634727, 0.1793742, 0.03215694, 
    -0.07124329, -0.1263051, -0.124938, -0.07111406, 0.1095495, 0.1719527, 
    0.12503, 0.4504358, 0.536113, 0.0665493, -0.1046423, 0.02157879, 
    -0.04687846, 0.151136, 0.7215793, 0.7238088, 0.4982386, 0.3656693, 
    0.2273064, 0.02859306, -0.1571326, -0.2977743, -0.2753782, -0.2444377, 
    -0.170577, -0.0140667, 0.05831289, 0.1640582, 0.2077913, 0.2824173, 
    0.3346634, 0.2125769, 0.1784472, -0.08351541, -0.2109246, -0.2461298, 
    -0.1897161,
  -0.4052281, -0.632962, -0.9615595, -0.9091016, -1.232083, -1.100817, 
    -0.5125522, -0.6066603, -0.1228062, 0.04672509, -0.6835157, -0.9672396, 
    -0.5028028, 0.2234015, 0.3257453, -0.2197137, -0.1557001, 0.315296, 
    -0.0385451, -0.1800653, -0.4442256, -0.4615107, -0.3160029, -0.639847, 
    -0.5594428, -0.206709, 0.04662743, -0.9224811, -0.8453974, 0.0892868, 
    -0.1848016, -0.3205597, -0.4022331, -0.5567739, -0.6957881, -0.9425817, 
    -0.9408396, -1.015026, -1.015579, -0.963138, -0.8504916, -0.8528515, 
    -0.7492383, -0.5650913, -0.4177279, -0.3305371, -0.2140336, -0.1903839, 
    -0.1633332, -0.07029939, -0.0276401, -0.03664088, -0.05140305, 
    0.04327464, 0.1957159, 0.190671, 0.01768899, -0.1612172, -0.2805212, 
    -0.2688675, -0.3529663, -0.3800011, -0.237227, -0.05503249, 0.01978827, 
    0.1963508, 0.4561001, 0.2370246, -0.005472183, 0.1927049, 0.1587856, 
    0.08819646, 0.2364385, 0.3295698, 0.289597, 0.2529271, 0.09955788, 
    -0.007098913, -0.1319854, -0.3410516, -0.2992873, -0.2376335, -0.3442414, 
    -0.3320994, -0.2456574, -0.1585968, -0.04686165, -0.08647776, 
    -0.09691095, -0.1142287, -0.1962767, -0.1059442, -0.2989125, -0.5158072, 
    -0.7020869, -0.6144073,
  -0.7283072, -1.046292, -1.166995, -0.9658726, -1.141068, -0.7372431, 
    -0.4896519, -0.7516312, -0.1395217, -0.01317072, -1.013887, -0.8037795, 
    0.0842088, 0.2336066, -0.2921746, -0.511885, 0.05850893, 0.1343879, 
    -0.1999383, -0.1914748, -0.1704461, -0.1007033, -0.04816425, -0.3646029, 
    -0.116833, 0.342526, 0.153496, -0.8903673, -0.1957064, 0.3347298, 
    -0.1311231, 0.009599566, -0.372155, -0.4887562, -0.3870802, -0.5456415, 
    -0.4858432, -0.6216508, -0.724027, -0.8536168, -0.9249382, -0.8914747, 
    -0.7204947, -0.5017774, -0.3777213, -0.1972039, -0.07737958, -0.05257511, 
    0.01054335, -0.001891613, -0.0570671, -0.1189977, -0.06146181, 0.1383917, 
    0.2845506, 0.1863084, -0.1680861, -0.4139681, -0.4539586, -0.585306, 
    -0.7465202, -0.6727084, -0.4152377, -0.2268101, -0.01185232, 0.2727342, 
    0.2959276, 0.0635708, 0.03987287, 0.06863263, -0.1435581, -0.1885614, 
    -0.04899406, 0.106442, 0.1620408, 0.04565078, -0.1389683, -0.3622756, 
    -0.616605, -0.680456, -0.6085973, -0.6963903, -0.7413935, -0.5864944, 
    -0.4105504, -0.2745966, -0.2420282, -0.3118362, -0.4311396, -0.5784049, 
    -0.6298864, -0.7519724, -0.7431678, -0.609362, -0.7924023, -0.7706414,
  -0.5838251, -0.7386103, -0.7714391, -0.8548701, -1.073701, -0.9587439, 
    -0.5657262, -0.4637077, -0.2728385, -0.4876823, -0.600264, 0.01545879, 
    0.1835578, -0.3874383, -0.7134801, -0.3157912, -0.1013869, -0.3408238, 
    -0.2846065, 0.2181768, 0.3524706, 0.4265918, 0.4624481, 0.3826456, 
    0.2585244, 0.3510375, -0.3202839, -0.3904333, 0.4978485, 0.242477, 
    -0.1865596, 0.1125945, -0.1851922, -0.1450721, 0.219772, -0.01333332, 
    -0.07529628, -0.1158071, -0.09650373, -0.1189485, -0.2038131, -0.2379117, 
    -0.1968794, -0.1037478, -0.05008602, -0.008370399, 0.03456593, 0.1487913, 
    0.1607056, 0.1199508, 0.1918259, 0.1489873, 0.1658006, 0.3338017, 
    0.3175263, 0.1161427, -0.2371128, -0.509948, -0.6259313, -0.7471715, 
    -0.816898, -0.7600946, -0.530163, -0.1892939, 0.05120087, 0.03748029, 
    -0.218314, -0.1638218, 0.2149706, 0.1981738, 0.05580711, 0.1254523, 
    0.1023078, 0.09532535, 0.08002567, -0.08520842, -0.2599318, -0.4870305, 
    -0.6990266, -0.8843453, -1.08817, -1.207685, -1.043216, -0.8318877, 
    -0.7233918, -0.522578, -0.5084991, -0.6279331, -0.6661, -0.7325068, 
    -0.7732295, -0.7895381, -0.700622, -0.5392612, -0.4612014, -0.4790074,
  -0.5819533, -0.6794298, -0.8834012, -0.951386, -0.7079942, -0.4748404, 
    -0.3222692, -0.1905632, -0.3649771, -0.3526726, 0.3136684, 0.314824, 
    -0.3224971, -0.6515008, -0.3212599, -0.1555699, -0.3551466, -0.3609085, 
    0.07952131, 0.3966437, 0.379456, 0.2633271, 0.1575973, 0.2441044, 
    0.1104937, -0.08760071, -0.2663932, -0.1123569, 0.1850712, -0.08869159, 
    -0.04886411, 0.3151333, 0.06659794, 0.07039045, -0.01548171, -0.411006, 
    -0.2479362, -0.06321931, 0.06951094, 0.3132458, 0.5949841, 0.80724, 
    0.8682098, 0.7903123, 0.6727834, 0.6140757, 0.5706348, 0.5217576, 
    0.4097781, 0.4023566, 0.5060678, 0.4830699, 0.4727511, 0.5263143, 
    0.3929644, 0.09397364, -0.2883658, -0.5212927, -0.6307971, -0.7466984, 
    -0.8266306, -0.8084826, -0.4036162, -0.03284848, -0.03094417, -0.1282424, 
    -0.1454625, -0.08766627, 0.2330048, 0.3327605, 0.1998174, 0.2043096, 
    0.2295866, 0.2421516, 0.2767708, 0.1952608, -0.05724621, -0.3641953, 
    -0.5818386, -0.7863975, -0.9357958, -1.081059, -1.238123, -1.282019, 
    -1.217858, -0.9325719, -0.749938, -0.8158722, -0.8227732, -0.7859564, 
    -0.7227564, -0.7069526, -0.685469, -0.6288122, -0.5885777, -0.5698929,
  -0.607522, -0.7441924, -0.8529656, -0.446048, 0.1769823, 0.4642545, 
    0.3818813, 0.2615526, 0.1882777, 0.270895, 0.3716437, -0.008011341, 
    -0.3365593, -0.07840508, 0.1389451, -0.2471389, -0.1395868, 0.1221483, 
    -0.01286155, 0.08582008, 0.1160121, -0.0735873, -0.1790725, -0.00975278, 
    0.07587549, 0.06523097, 0.1866178, 0.04556966, 0.004879385, -0.05418622, 
    -0.03952146, -0.02747726, -0.153926, -0.07394564, -0.09569001, 
    -0.4022827, -0.1140499, 0.5805464, 0.4395967, 0.4703255, 0.5859332, 
    0.6155725, 0.5589328, 0.5189095, 0.5537567, 0.592917, 0.5302219, 
    0.4041963, 0.4667125, 0.6175914, 0.6128879, 0.5862598, 0.688067, 
    0.7363739, 0.5664682, 0.2154746, -0.1472869, -0.4021039, -0.6546426, 
    -0.8482618, -0.9054227, -0.8471873, -0.449922, -0.1270868, -0.1707717, 
    -0.06222677, 0.1661099, 0.2486136, 0.26209, 0.5438932, 0.5579394, 
    0.3923959, 0.4463997, 0.4760706, 0.3829072, 0.1994269, -0.01740146, 
    -0.1835318, -0.2956753, -0.675786, -1.027137, -1.303195, -1.536624, 
    -1.561608, -1.484704, -1.297725, -1.120918, -1.050883, -0.7912793, 
    -0.3662629, -0.2686715, -0.4105823, -0.4944041, -0.5085478, -0.577803, 
    -0.5727574,
  -0.1108263, -0.1122589, 0.08967781, 0.3580532, 0.5204067, 0.65763, 
    0.6730597, 0.6228155, 0.5692186, 0.5253873, 0.3078904, 0.2269986, 
    0.1926886, 0.1761684, 0.03463185, -0.08039069, 0.08915657, 0.235348, 
    0.1519334, 0.07299459, 0.1776821, 0.06399399, 0.06025052, 0.06929995, 
    -0.1655798, -0.1015497, 0.1164193, -0.1424184, -0.2173047, 0.04719758, 
    0.02546883, -0.07791591, -0.06675053, -0.109834, -0.1728058, -0.1625361, 
    0.1265745, 0.4673138, 0.5875945, 0.1425738, -0.006596565, -0.09100342, 
    -0.1499877, -0.1165733, -0.04383564, 0.04970312, 0.1795545, 0.2657847, 
    0.3200979, 0.3606405, 0.3423624, 0.4209108, 0.5546508, 0.5915651, 
    0.428267, -0.01043797, -0.3852744, -0.4993529, -0.6106157, -0.7829947, 
    -0.8263702, -0.7506378, -0.3909212, 0.0683071, 0.3114712, 0.3001595, 
    0.1905079, 0.1687303, 0.2175088, 0.6257777, 0.5208139, 0.3815556, 
    0.4832813, 0.5882294, 0.7967901, 0.3474905, 0.199671, 0.01106524, 
    -0.2765818, -0.6474965, -1.033743, -1.144535, -1.103779, -1.086722, 
    -1.108955, -1.095837, -1.078177, -1.034037, -0.7731318, -0.319665, 
    -0.1354852, -0.1107292, -0.03364563, -0.09541321, -0.2152542, -0.2013869,
  0.1647265, 0.1227993, 0.550078, 0.6211392, 0.6371872, 0.9820117, 1.020846, 
    0.7537241, 0.8535938, 1.107614, 1.21681, 1.166012, 0.7352341, 0.3911261, 
    0.4328578, 0.4203578, 0.3868454, 0.3613246, 0.4164515, 0.4148076, 
    0.2702602, 0.2113247, 0.1923957, 0.02577782, -0.1554559, -0.06522161, 
    0.01910472, -0.07235003, 0.1316538, 0.2150848, 0.0009410381, -0.01569319, 
    -0.09363937, -0.2270379, -0.05526018, 0.1804163, 0.235055, 0.5419405, 
    0.9684539, 1.153675, 1.137756, 1.020634, 0.7892537, 0.5550251, 0.3987269, 
    0.3446577, 0.4568322, 0.6242321, 0.7060843, 0.6594856, 0.6721652, 
    0.6284964, 0.4145966, 0.2205863, 0.1076956, -0.1346548, -0.3727407, 
    -0.4407089, -0.5171249, -0.5973008, -0.466572, -0.2181513, 0.107337, 
    0.4366826, 0.3873664, 0.2624153, 0.2021453, 0.3398075, 0.5011029, 
    0.5338507, 0.3712693, 0.3580046, 0.3664028, 0.3679165, 0.01925111, 
    -0.08535498, -0.12515, -0.1850131, -0.1757032, -0.05192375, -0.5148952, 
    -0.4004581, -0.2438989, -0.2904162, -0.4393582, -0.6210318, -0.8031449, 
    -0.8643594, -0.6376824, -0.2693558, 0.01106405, 0.2291141, 0.4483685, 
    0.5555792, 0.5926559, 0.4171515,
  0.5795054, 0.805205, 1.036064, 0.7501109, 0.4896451, 0.6373498, 0.8306608, 
    0.8986785, 1.141972, 1.264775, 1.117266, 0.8837043, 0.7071254, 0.6428188, 
    0.7442349, 0.8046515, 0.6613898, 0.5572068, 0.5916632, 0.5109667, 
    0.3805143, 0.2674119, 0.1363735, -0.1016474, -0.1379266, -0.1359732, 
    -0.1669626, -0.196146, -0.06287766, -0.1427107, -0.2450385, -0.2577343, 
    -0.3005075, -0.1969268, 0.1310842, 0.2407684, 0.1162565, 0.5336721, 
    1.379309, 2.208085, 1.18276, 0.608135, 0.2817024, 0.1249803, 0.06705379, 
    0.1911589, 0.3331511, 0.4148078, 0.5444627, 0.7314255, 0.8591437, 
    0.8716601, 0.7983853, 0.6702929, 0.5009081, 0.1765751, -0.199971, 
    -0.4129103, -0.4372756, -0.2297721, 0.06049454, 0.2389126, 0.2392217, 
    0.2137661, 0.2368944, 0.2328743, 0.2326956, 0.2757618, 0.2830532, 
    0.2605761, 0.192119, 0.1527309, 0.1061814, 0.03598291, -0.0250361, 
    -0.0470413, -0.09214222, -0.2750199, -0.3335321, -0.2809931, -0.06401694, 
    0.1680305, 0.2055142, -0.08629799, -0.1361842, -0.03011322, 0.09586239, 
    0.2725387, 0.3845992, 0.4466755, 0.56287, 0.7661419, 0.9121377, 
    0.8987105, 0.813473, 0.6545537,
  0.880205, 1.103106, 1.02848, 0.5356737, 0.3755337, 0.5046027, 0.7123663, 
    0.7041959, 0.6555468, 0.5386033, 0.3512661, 0.1690232, 0.2223598, 
    0.3591111, 0.4191697, 0.3621222, 0.3538053, 0.4516895, 0.5661263, 
    0.5082977, 0.3788869, 0.2930467, 0.1371549, -0.007262707, -0.09575534, 
    -0.1469597, -0.1708528, -0.2205112, -0.3373082, -0.4137081, -0.3919792, 
    -0.3174834, -0.2507679, -0.08957028, 0.1078581, 0.2228971, 0.3202928, 
    0.9778936, 0.9850223, 0.9097781, -0.6338413, -1.142223, -0.619144, 
    -0.5260451, -0.2357129, 0.2104785, 0.5965134, 0.7554002, 0.8336552, 
    0.8737106, 0.7646612, 0.6096644, 0.5823534, 0.5624152, 0.2787563, 
    -0.2393265, -0.5469274, -0.3934278, -0.00218448, 0.2774217, 0.3292285, 
    0.08604813, 0.1972458, 0.2709275, 0.3221645, 0.3562467, 0.4089648, 
    0.415166, 0.3641405, 0.3176723, 0.2980109, 0.235755, 0.266354, 0.4196578, 
    0.4934537, 0.4126596, 0.04825503, -0.2335483, -0.3007196, -0.1643751, 
    -0.08445954, -0.02583337, -0.4702182, -0.8190303, -0.5144078, 0.01015306, 
    0.4176724, 0.6830859, 0.7454879, 0.7411423, 0.9097457, 1.142477, 
    1.211732, 1.081849, 0.8733526, 0.7696092,
  0.959518, 0.9498501, 0.7359177, 0.3777471, 0.3454556, 0.1775357, 0.1542283, 
    0.1338507, 0.03868472, -0.02010432, -0.09510434, -0.1502312, -0.1087436, 
    -0.07907245, -0.1403354, -0.2442256, -0.3110387, -0.306644, -0.338968, 
    -0.2975457, -0.2989616, -0.2745314, -0.2340524, -0.2158558, -0.242972, 
    -0.3135452, -0.3460644, -0.3446485, -0.3231481, -0.2971878, -0.3282251, 
    -0.320348, -0.3729191, -0.1419629, 0.1089159, 0.3502736, 0.4549775, 
    0.4018521, 0.03931952, -0.9922396, -1.889587, -1.812944, -0.6036164, 
    -0.3103223, -0.1669626, 0.5142875, 0.8756475, 0.7997363, 0.6638968, 
    0.4058402, 0.1181614, -0.1173859, -0.1040397, -0.1200716, -0.4503614, 
    -0.7229201, -0.7017282, -0.203861, 0.290036, 0.2995086, -0.2227409, 
    0.1109668, 0.4532518, 0.6169074, 0.5179653, 0.3307257, 0.3130825, 
    0.3859015, 0.3569139, 0.2702765, 0.2046026, 0.08424115, 0.04412103, 
    -0.01292682, -0.09556007, -0.2722852, -0.6626337, -0.7342646, -0.61903, 
    -0.5050652, -0.7373893, -0.9651729, -1.220609, -0.8245801, 0.008704126, 
    0.5501104, 0.7465948, 0.7907192, 0.8572557, 0.9589971, 0.9651169, 
    0.8598598, 0.7458298, 0.7428024, 0.7953578, 0.8508917,
  -0.3731642, -0.3558953, -0.1095412, -0.1531773, -0.1724156, 0.03368795, 
    -0.1977736, -0.1688674, -0.1224806, -0.1482944, -0.2143589, -0.2615432, 
    -0.2741245, -0.2801792, -0.2895379, -0.3258986, -0.3497106, -0.4094111, 
    -0.4697138, -0.4699905, -0.4871454, -0.4352249, -0.4120477, -0.4105015, 
    -0.4338901, -0.4877476, -0.4814489, -0.4193394, -0.3463739, -0.2616894, 
    -0.1929722, -0.1622751, -0.0738802, 0.1279752, 0.2740364, 0.2325162, 
    0.06000632, -0.1369175, -0.3525749, -0.5459502, -0.5174019, -0.3332393, 
    -0.2024934, -0.05234694, 0.1738088, 0.3505509, 0.2525198, -0.7036982, 
    -1.260535, -1.528145, -1.546488, -1.397562, -0.6094105, -0.4274933, 
    -0.3362339, -0.3396029, -0.1965206, 0.1098921, 0.2701628, 0.1907841, 
    0.1800095, 0.3172166, 0.4346482, 0.4109991, 0.2560187, 0.1454881, 
    0.1572555, 0.2193651, 0.225729, 0.125908, 0.0582974, 0.01667947, 
    0.06799787, 0.01763979, -0.1349155, -0.3083693, -0.5715204, -0.6857781, 
    -0.7766473, -0.7143263, -0.8873895, -1.220365, -1.11973, -0.4906285, 
    -0.05508173, 0.2589482, 0.2630501, 0.255856, 0.327373, 0.3313607, 
    0.1736621, -0.06416368, -0.1741897, -0.1470413, -0.1419305, -0.256937,
  -1.108858, -0.9628291, -0.7030797, -0.3257521, -0.3084018, -0.4352899, 
    -0.5652052, -0.5823276, -0.5710483, -0.5105667, -0.4277379, -0.3411657, 
    -0.3361363, -0.3918004, -0.4582392, -0.4714554, -0.4048049, -0.5337274, 
    -0.6049352, -0.644014, -0.6729202, -0.603568, -0.5300815, -0.4622267, 
    -0.4579299, -0.4794143, -0.4539422, -0.3987829, -0.2957879, -0.162943, 
    -0.02414083, 0.07125318, 0.1483201, 0.1718065, 0.09342106, -0.05833676, 
    -0.3001661, -0.3846551, -0.3702183, -0.2366245, -0.1692743, -0.1152866, 
    -0.09901065, 0.02512681, 0.232142, 0.4581344, 0.5105925, 0.4201472, 
    0.2468393, 0.1244271, 0.07200181, -0.003828168, 0.006963253, -0.01160789, 
    -0.00408864, 0.03780603, 0.1015592, 0.1429327, 0.1480596, 0.141533, 
    0.1021287, 0.09184226, 0.04949202, -0.02485695, -0.07181334, -0.0557977, 
    0.06140608, 0.1901821, 0.1756964, 0.04421857, -0.07560565, -0.1729852, 
    -0.2297886, -0.195967, -0.1721714, -0.2664585, -0.3553582, -0.4434767, 
    -0.4756219, -0.5752314, -0.6945512, -0.5775099, -0.3074412, -0.05159831, 
    0.1598268, 0.1717417, 0.2935514, 0.3776169, 0.5953407, 0.6270137, 
    0.2418261, -0.03130245, -0.2833204, -0.5239127, -0.7928417, -1.031156,
  -1.083548, -0.9918654, -1.009248, -1.155814, -1.331107, -1.204252, 
    -1.15378, -0.8870639, -0.5578647, -0.3042514, -0.2286818, -0.1179721, 
    -0.2722529, -0.6015823, -0.6979527, -0.6942744, -0.6196813, -0.5767452, 
    -0.5902052, -0.6206579, -0.5691441, -0.4577345, -0.3236851, -0.3033563, 
    -0.344437, -0.3533075, -0.3355341, -0.2331579, -0.1247265, -0.00705111, 
    0.04469037, 0.04286766, 0.002617002, -0.0579136, -0.07114598, -0.1149611, 
    -0.08607119, 0.0414027, 0.1863897, 0.2991829, 0.3657681, 0.3699509, 
    0.4340461, 0.5521939, 0.6794562, 0.7680305, 0.7773241, 0.6392543, 
    0.4775845, 0.3383918, 0.2446092, 0.1562304, 0.1003225, 0.01109719, 
    0.01791692, -0.009687185, -0.01014328, -0.04691088, -0.04240268, 
    -0.08275098, -0.09844095, -0.1009475, -0.1627965, -0.1799512, -0.167663, 
    -0.0138869, 0.1358201, 0.1748989, 0.09543926, 0.007483542, -0.06883481, 
    -0.08291352, -0.04126322, -0.01040381, -0.08017921, -0.0390659, 
    -0.1420119, -0.2220086, -0.458988, -0.6577995, -0.6317581, -0.5207877, 
    -0.2369339, 0.1587367, 0.3535938, 0.3504362, 0.2089159, 0.103854, 
    0.1803514, 0.2088833, 0.1054652, -0.1577346, -0.6748244, -1.160762, 
    -1.23555, -1.178519,
  -0.7408564, -0.7917027, -0.8054233, -0.7912958, -0.7094923, -0.5327346, 
    -0.2734408, -0.07990265, 0.06938112, -0.02230144, -0.1347688, -0.3607455, 
    -0.515954, -0.5563346, -0.4848179, -0.3113967, -0.3059443, -0.2277378, 
    -0.1020217, -0.02755877, 0.01921858, 0.05849266, 0.09054017, 0.1070278, 
    0.04745752, -0.04645526, -0.1251826, -0.1124868, 0.009062529, 0.1921026, 
    0.2653447, 0.3163866, 0.3250617, 0.3429328, 0.3652961, 0.2239873, 
    0.379326, 0.4636196, 0.5976691, 0.6524868, 0.5930467, 0.583102, 
    0.5648729, 0.5630337, 0.5355109, 0.4849412, 0.380384, 0.2603644, 
    0.158216, 0.07649398, 0.01389635, -0.03390646, -0.0472846, -0.05023098, 
    -0.05550432, -0.07765603, -0.1416214, -0.2222852, -0.2872103, -0.3592644, 
    -0.4092643, -0.4203321, -0.300638, -0.3171257, -0.222334, -0.09407899, 
    -0.02464536, 0.01082014, 0.009192526, 0.030742, -0.07648455, -0.1124058, 
    -0.1384637, -0.1702019, -0.2082065, -0.3057325, -0.4280634, -0.6844761, 
    -0.6079137, -0.5154982, -0.4974971, -0.2271678, 0.1441538, 0.4354625, 
    0.3252734, 0.02843082, -0.1554387, -0.1448927, 0.09493446, 0.2347624, 
    0.2810351, 0.2429491, 0.08064434, -0.1286655, -0.5642287, -0.6589715,
  -0.6344435, -0.4731153, -0.2661653, -0.03901672, -0.09503889, -0.211966, 
    -0.1738801, -0.07523084, -0.08943939, -0.1437042, -0.1724641, -0.1860222, 
    -0.1794469, -0.08278346, 0.05642569, 0.1311488, 0.2017542, 0.2210577, 
    0.182223, 0.1465459, 0.1521775, 0.1665003, 0.1336716, 0.08219039, 
    0.1552699, 0.1643357, 0.1972134, 0.2660773, 0.3625454, 0.4358364, 
    0.5552212, 0.5763962, 0.6196579, 0.5598272, 0.5215949, 0.4691535, 
    0.4288214, 0.4042284, 0.3918748, 0.3842577, 0.3563443, 0.3283658, 
    0.2925421, 0.253333, 0.2183558, 0.1986293, 0.1867802, 0.1689906, 
    0.1292119, 0.07955396, 0.005904555, -0.08201826, -0.176338, -0.2598503, 
    -0.3464552, -0.4251173, -0.481351, -0.5081089, -0.4949578, -0.4676465, 
    -0.4251825, -0.3830274, -0.3593946, -0.334232, -0.2698114, -0.3213088, 
    -0.3151401, -0.3350295, -0.3862339, -0.4459832, -0.4907912, -0.5161331, 
    -0.5762731, -0.547253, -0.6586298, -0.6855829, -0.6300002, -0.668135, 
    -0.6118683, -0.4110389, -0.230505, 0.05142879, 0.2097301, 0.1503059, 
    -0.06442401, -0.2598504, -0.3646352, -0.2934771, -0.1232128, -0.01299143, 
    0.03490901, 0.01903963, -0.04375356, -0.1721714, -0.2810418, -0.4172072,
  -0.2511591, -0.1841342, -0.06214523, -0.03081369, 0.08593416, 0.1680632, 
    0.2185838, 0.211341, 0.2268356, 0.2164842, 0.2393681, 0.2690232, 
    0.3074834, 0.3598598, 0.3859502, 0.3979131, 0.377845, 0.3272427, 
    0.2662402, 0.1983691, 0.1287239, 0.08464837, 0.07066727, 0.04988277, 
    0.1590462, 0.2016406, 0.2822396, 0.3800746, 0.4372849, 0.4927048, 
    0.5389614, 0.5544236, 0.5481735, 0.5321091, 0.5112271, 0.498662, 
    0.4876919, 0.4623664, 0.4183885, 0.3538377, 0.2880337, 0.2159959, 
    0.1455369, 0.07087871, -0.007946163, -0.09835958, -0.1996779, -0.2937046, 
    -0.3795282, -0.4608108, -0.5407587, -0.6145706, -0.676566, -0.7057489, 
    -0.6956252, -0.667077, -0.6422561, -0.6054884, -0.5410353, -0.4704624, 
    -0.4149448, -0.3843296, -0.3831577, -0.404284, -0.4313674, -0.4335809, 
    -0.4486036, -0.468672, -0.4887892, -0.5130731, -0.5357782, -0.387536, 
    -0.3745966, -0.3125848, -0.2787145, -0.2455763, -0.2009474, -0.1796421, 
    -0.139668, -0.07733083, -0.04735041, -0.03493172, -0.03524104, 
    -0.0554235, -0.06865501, -0.04793596, 0.02515936, 0.08087206, 0.1024051, 
    0.103301, 0.0566535, -0.06232429, -0.1277866, -0.2154656, -0.2455438, 
    -0.266898,
  -0.1102898, -0.09137702, -0.05342144, -0.01487982, 0.04080045, 0.09923148, 
    0.1419563, 0.181442, 0.215345, 0.2348112, 0.2491829, 0.2566373, 
    0.2606087, 0.2516894, 0.2392708, 0.2185352, 0.1904101, 0.1613085, 
    0.140524, 0.1370084, 0.1515429, 0.1835415, 0.2337532, 0.2829392, 
    0.340231, 0.4024541, 0.4496221, 0.483639, 0.4913539, 0.4961064, 
    0.4958135, 0.4849737, 0.4635546, 0.4311489, 0.3972622, 0.362106, 
    0.3225551, 0.2721971, 0.2262498, 0.1714321, 0.117005, 0.057923, 
    -0.004642107, -0.06077817, -0.1066603, -0.1491571, -0.1887079, 
    -0.2281447, -0.2596877, -0.2880894, -0.3065952, -0.3225946, -0.3440464, 
    -0.3591506, -0.3610549, -0.3624546, -0.360062, -0.3591994, -0.3564813, 
    -0.3521681, -0.3499383, -0.3540724, -0.3603875, -0.3649123, -0.3535516, 
    -0.3302118, -0.303161, -0.2793329, -0.2555373, -0.229577, -0.1997756, 
    -0.1792027, -0.1746616, -0.1633986, -0.1380243, -0.1444207, -0.1152703, 
    -0.0793654, -0.06574236, -0.04285824, -0.03725928, 0.0316698, 0.05046856, 
    0.06521451, 0.02073216, 0.1428676, 0.1436976, 0.1190556, 0.09436488, 
    0.02807271, -0.01154327, -0.04403013, -0.06085956, -0.08773129, 
    -0.1121942, -0.1197789,
  -0.2414748, -0.23223, -0.2139683, -0.1928583, -0.1743361, -0.1545607, 
    -0.1396193, -0.1239781, -0.1023147, -0.08520865, -0.06276405, 
    -0.04036808, -0.01575875, 0.005774498, 0.02533829, 0.04563445, 
    0.06674445, 0.09742481, 0.1212367, 0.1496547, 0.1781865, 0.2067998, 
    0.2423956, 0.2697718, 0.2953578, 0.3165492, 0.340654, 0.3596483, 
    0.3793911, 0.3801235, 0.3790004, 0.3789029, 0.3697231, 0.3584113, 
    0.3466274, 0.3317186, 0.3067023, 0.2824022, 0.2514614, 0.2164679, 
    0.178675, 0.1470018, 0.111699, 0.07628238, 0.03897762, 0.009013474, 
    -0.0231154, -0.05050802, -0.07884455, -0.1069859, -0.1352085, -0.1642124, 
    -0.1871617, -0.2141311, -0.2371128, -0.260534, -0.2770867, -0.2951694, 
    -0.3129591, -0.3212111, -0.3248732, -0.3271355, -0.3256382, -0.32681, 
    -0.3277378, -0.3219436, -0.3107131, -0.301159, -0.2972202, -0.290547, 
    -0.2856968, -0.285827, -0.2830275, -0.2766636, -0.2710809, -0.2723667, 
    -0.2697463, -0.2691766, -0.264424, -0.2618198, -0.257702, -0.2587925, 
    -0.2625197, -0.2670933, -0.2752476, -0.281286, -0.2870314, -0.2927118, 
    -0.298327, -0.2955275, -0.2926304, -0.2865269, -0.2807977, -0.2771194, 
    -0.2673863, -0.2553095,
  -0.2539001, -0.2426858, -0.2346289, -0.230463, -0.2294695, -0.2310971, 
    -0.2358497, -0.2438412, -0.2541113, -0.2663997, -0.2808529, -0.2949967, 
    -0.3095315, -0.3242451, -0.3391535, -0.3541927, -0.3695412, -0.3851988, 
    -0.4004166, -0.4146583, -0.4277442, -0.4395444, -0.4501235, -0.4577248, 
    -0.4627538, -0.4653256, -0.463454, -0.4575946, -0.447015, -0.4318786, 
    -0.4130309, -0.3916442, -0.368711, -0.3428321, -0.3131607, -0.2844341, 
    -0.2555274, -0.2260514, -0.1972918, -0.1697525, -0.1450944, -0.1230241, 
    -0.1048601, -0.09162784, -0.08389676, -0.08158541, -0.06089878, 
    -0.07087588, -0.09332037, -0.1272724, -0.167702, -0.1956804, -0.1107521, 
    -0.1314714, -0.1247821, -0.1832781, -0.2272072, -0.2805927, -0.2823017, 
    -0.258913, -0.3360286, -0.3351173, -0.3989031, -0.3867447, -0.3989356, 
    -0.4064064, -0.4027119, -0.3841572, -0.3731055, -0.3862405, -0.3807716, 
    -0.3649511, -0.3199971, -0.2239194, -0.3246193, -0.3129659, -0.2578714, 
    -0.2143331, -0.2613707, -0.2704692, -0.2653747, -0.2672954, -0.2762146, 
    -0.2837343, -0.2947855, -0.3064561, -0.3160267, -0.3214617, -0.324717, 
    -0.3251567, -0.3219829, -0.3156514, -0.3074484, -0.2951922, -0.2816992, 
    -0.2672954,
  -0.3462826, -0.3361263, -0.324847, -0.3194108, -0.3206966, -0.3306738, 
    -0.3447851, -0.3622495, -0.3828386, -0.4033951, -0.4226498, -0.4408953, 
    -0.4563249, -0.4700618, -0.4813899, -0.4917415, -0.5038674, -0.521348, 
    -0.5453063, -0.5757746, -0.6096613, -0.6447201, -0.6725523, -0.693711, 
    -0.7050231, -0.70696, -0.7036886, -0.694037, -0.6832781, -0.6756124, 
    -0.6753192, -0.6793394, -0.68362, -0.682888, -0.6705012, -0.6416445, 
    -0.5930929, -0.5245218, -0.4404721, -0.3452568, -0.2350032, -0.1629329, 
    -0.1165625, -0.06023121, -0.03363633, -0.02527046, -0.04708028, 
    -0.08013678, -0.1116638, -0.06887388, -0.1241961, -0.1681256, 
    -0.08661485, -0.2283788, -0.1567156, -0.2867451, -0.3169374, -0.3383884, 
    -0.3942485, -0.4294043, -0.4826598, -0.552598, -0.5872657, -0.6001073, 
    -0.6104915, -0.6186458, -0.5979915, -0.5800717, -0.5883723, -0.598171, 
    -0.6090922, -0.5870867, -0.5407488, -0.4710221, -0.4201274, -0.3466082, 
    -0.2562274, -0.1794205, -0.05764323, 0.01691711, 0.07542944, 0.1909895, 
    0.0775454, 0.2169008, 0.1444073, 0.113287, 0.04242229, -0.03443384, 
    -0.1143484, -0.1902447, -0.2537694, -0.3020117, -0.3325293, -0.3525815, 
    -0.3650162, -0.3604101,
  -0.4739681, -0.4670345, -0.4492286, -0.4355241, -0.4128027, -0.3800229, 
    -0.346543, -0.3168229, -0.3013284, -0.3056902, -0.3169369, -0.326556, 
    -0.3266699, -0.3218849, -0.3295672, -0.3583431, -0.412396, -0.48528, 
    -0.5568457, -0.6005635, -0.5929625, -0.5192969, -0.4066179, -0.3205013, 
    -0.3087988, -0.3441667, -0.3731868, -0.3818623, -0.3761331, -0.3798118, 
    -0.4040785, -0.4450946, -0.5052178, -0.5741305, -0.6380639, -0.6808701, 
    -0.679893, -0.6367779, -0.5559015, -0.4428644, -0.3142519, -0.1904073, 
    0.01401997, 0.08566713, 0.1024964, 0.1244693, 0.1120996, 0.07289066, 
    0.02484378, -0.02496105, -0.0790301, -0.1286395, -0.1327736, -0.1050717, 
    -0.06994796, -0.03951192, -0.03659856, -0.0654397, -0.1266214, 
    -0.1982522, -0.277207, -0.338291, -0.3768002, -0.3815852, -0.3623307, 
    -0.320485, -0.2716082, -0.2124772, -0.1504819, -0.08134151, -0.01368189, 
    0.02638984, 0.02948213, -0.02826524, -0.07334995, -0.1361588, -0.1328385, 
    -0.1270931, -0.1204036, -0.06024735, 0.01135096, 0.09868801, 0.159707, 
    0.2239159, 0.2782614, 0.322174, 0.3257229, 0.3196678, 0.2578838, 
    0.1225324, -0.009954453, -0.1709733, -0.3107195, -0.4186623, -0.4754009, 
    -0.4938902,
  -0.7772074, -0.7321715, -0.6632912, -0.6147401, -0.5891055, -0.5747002, 
    -0.5528907, -0.5326107, -0.5180763, -0.5109147, -0.5146093, -0.5163834, 
    -0.480853, -0.4206805, -0.3577248, -0.2964291, -0.274196, -0.2851986, 
    -0.3245542, -0.4330504, -0.4844661, -0.5004816, -0.4681251, -0.4217708, 
    -0.3637955, -0.3451921, -0.3545836, -0.3761005, -0.4017678, -0.4240495, 
    -0.441237, -0.4476985, -0.4486591, -0.4574156, -0.4870863, -0.546299, 
    -0.6366963, -0.7219176, -0.7429795, -0.6754832, -0.5611753, -0.4384375, 
    -0.2422957, -0.03788471, 0.04085922, 0.09181952, 0.2083557, 0.2270899, 
    0.250283, 0.2274479, 0.2278874, 0.198265, 0.1294011, 0.09701157, 
    0.09660482, 0.09387016, 0.0341208, 0.01984692, -0.08541036, -0.2264421, 
    -0.3096128, -0.3874285, -0.4454689, -0.5442319, -0.6492612, -0.671185, 
    -0.6301529, -0.5465431, -0.4356055, -0.3063252, -0.1870379, -0.07676792, 
    0.01100898, 0.05822563, 0.08589494, 0.1235415, 0.1317122, 0.09662092, 
    0.05015302, 0.03275394, -0.007805943, 0.01292972, 0.01338545, 0.06389001, 
    0.1292383, 0.1667383, 0.1940169, 0.189085, 0.08649731, 0.1587627, 
    0.06883788, -0.09978247, -0.3255954, -0.5978293, -0.7796483, -0.838747,
  -0.0505147, -0.05049849, -0.08466196, -0.1022401, -0.05043316, -0.05588579, 
    -0.04118824, -0.04904938, 0.005914211, -0.1173115, -0.2199159, 
    -0.2879009, -0.3032494, -0.2995703, -0.2938738, -0.1436296, -0.01062131, 
    0.06556606, 0.04017582, 0.04251933, -0.1479754, -0.3750749, -0.5167747, 
    -0.5698833, -0.5545835, -0.505609, -0.4597104, -0.4506121, -0.4812274, 
    -0.5111101, -0.5362735, -0.5443625, -0.5114843, -0.4616146, -0.4132748, 
    -0.3979753, -0.3883235, -0.4058691, -0.4295508, -0.419655, -0.3680439, 
    -0.308522, -0.2524838, -0.1899676, -0.1609964, -0.03301787, 0.1748275, 
    0.3688865, 0.4733626, 0.5472722, 0.5871322, 0.6084701, 0.6128321, 
    0.6065333, 0.5395735, 0.4532942, 0.355638, 0.2636133, 0.1365297, 
    0.0363344, -0.05163765, -0.1512303, -0.2258074, -0.2632754, -0.3405054, 
    -0.4084253, -0.4462342, -0.5242128, -0.511306, -0.4947858, -0.3041933, 
    -0.2122006, -0.116514, 0.03726208, 0.1600485, 0.2632712, 0.4361553, 
    0.5278547, 0.4936263, 0.5246322, 0.4484928, 0.4204167, 0.3565495, 
    0.3090235, 0.2555567, 0.1842188, 0.1194727, 0.09655607, 0.1307845, 
    0.1388733, 0.1403058, -0.004909039, 0.102757, 0.06406879, 0.02147436, 
    0.006972313,
  -0.2205176, -0.2438416, 0.1361394, 0.04733706, 0.04369116, 0.1150937, 
    0.1897037, 0.2656965, 0.3530335, 0.436774, 0.4478908, 0.5148177, 
    0.4929094, 0.4005108, 0.2096415, 0.05721664, 0.09058237, 0.05641925, 
    0.04805326, 0.04821587, -0.04218102, -0.1089621, -0.1663189, -0.1373644, 
    -0.1675406, -0.08344173, 0.03517818, 0.0907445, 0.0595603, -0.09678745, 
    -0.2411237, -0.3221784, -0.3136334, -0.2408957, -0.1776958, -0.1412864, 
    -0.1307716, -0.1194761, -0.0544045, 0.03150058, 0.1018944, 0.1005108, 
    0.07334566, 0.05894172, -0.08370125, 0.030882, 0.216543, 0.4961003, 
    0.6817448, 0.788239, 0.7891993, 0.7088607, 0.6642644, 0.7129785, 
    0.7605046, 0.8563868, 0.9747787, 1.05847, 1.026748, 0.9499903, 0.8486718, 
    0.7147201, 0.6520411, 0.5336003, 0.3458887, 0.2155013, 0.1810775, 
    0.2028712, 0.3175033, 0.4287987, 0.3741114, 0.2377507, 0.2257227, 
    0.2277409, 0.3072167, 0.5016667, 0.7519431, 0.9914613, 0.7297429, 
    0.9183658, 0.7873438, 0.7448795, 0.690957, 0.6570378, 0.6115463, 
    0.5120671, 0.3914779, 0.2841211, 0.2554916, 0.306224, 0.3541406, 
    0.3711325, 0.2896059, 0.06511021, -0.209532, -0.2737079,
  1.929662, 1.69431, 1.558584, 1.510798, 1.552481, 1.569326, 1.359138, 
    1.179108, 1.091511, 1.264948, 1.608535, 1.863662, 1.879092, 1.651878, 
    1.2836, 0.8928449, 0.5419662, 0.4089417, 0.4087305, 0.4897685, 0.6558656, 
    0.7367574, 0.6296287, 0.5244367, 0.4373436, 0.5700259, 0.635309, 
    0.8594141, 1.007591, 1.010098, 0.8614972, 0.7661691, 0.6893454, 
    0.4017639, 0.4253318, 0.3901105, 0.2271223, 0.6584373, 0.7722235, 
    0.8225808, 0.732151, 0.691201, 0.6607485, 0.6741116, 0.7407776, 
    0.8678125, 1.048363, 1.255345, 1.479368, 1.704922, 1.893252, 2.006777, 
    1.999062, 1.869912, 1.735537, 1.699844, 1.751243, 1.816722, 1.858177, 
    1.91363, 2.009609, 2.158112, 2.282786, 2.272142, 2.091576, 1.790794, 
    1.464281, 1.214736, 1.065664, 1.008682, 1.004971, 1.015469, 1.010309, 
    0.9915918, 0.9494857, 0.9336491, 1.008079, 1.222272, 1.502822, 1.567715, 
    1.634365, 1.590648, 1.642406, 1.784935, 1.930963, 1.946279, 1.903115, 
    1.868821, 1.758503, 1.736611, 1.800771, 1.829401, 1.90279, 1.977367, 
    2.060537, 2.056891,
  2.864166, 2.837425, 2.771182, 2.754401, 2.889329, 3.071442, 3.169602, 
    3.09942, 2.899632, 2.749827, 2.757135, 2.951455, 3.17984, 3.339248, 
    3.346849, 3.247011, 3.096002, 2.921165, 2.763646, 2.691705, 2.690501, 
    2.726097, 2.769586, 2.78858, 2.724681, 2.552285, 2.439834, 2.462425, 
    2.596295, 2.757624, 2.882835, 2.971133, 3.0121, 3.041998, 3.011416, 
    2.898493, 2.80126, 2.843626, 2.939703, 2.975527, 2.876146, 2.702399, 
    2.548867, 2.422776, 2.366771, 2.391836, 2.434153, 2.494944, 2.585455, 
    2.659414, 2.710976, 2.830719, 2.961253, 3.022255, 3.024371, 2.959755, 
    2.878017, 2.788906, 2.729759, 2.729531, 2.850559, 3.022402, 3.164948, 
    3.256435, 3.244733, 3.148802, 2.95663, 2.68487, 2.392161, 2.103343, 
    1.803652, 1.555344, 1.428733, 1.398183, 1.413157, 1.428456, 1.46568, 
    1.57774, 1.764491, 2.018284, 2.258762, 2.399648, 2.491835, 2.631484, 
    2.751601, 2.783355, 2.713515, 2.567389, 2.45427, 2.39068, 2.389817, 
    2.435374, 2.539541, 2.657998, 2.749079, 2.8232,
  2.39055, 2.42403, 2.324681, 2.192226, 2.159804, 2.252106, 2.419912, 
    2.580247, 2.64291, 2.582346, 2.519717, 2.547663, 2.63404, 2.752854, 
    2.89584, 3.045791, 3.137165, 3.143252, 3.088873, 3.01944, 2.994472, 
    3.014801, 3.101715, 3.240061, 3.346686, 3.350266, 3.25777, 3.200038, 
    3.224355, 3.273167, 3.296247, 3.276276, 3.2461, 3.27294, 3.308356, 
    3.249355, 3.121507, 3.117048, 3.237457, 3.404092, 3.51931, 3.505622, 
    3.349355, 3.144358, 3.005052, 2.91791, 2.835439, 2.748054, 2.698639, 
    2.725608, 2.817942, 2.976862, 3.170449, 3.354661, 3.507965, 3.641559, 
    3.691868, 3.665826, 3.592551, 3.545595, 3.552675, 3.564264, 3.507477, 
    3.402643, 3.411578, 3.391819, 3.281419, 3.16402, 3.054466, 2.882786, 
    2.69291, 2.541038, 2.374062, 2.235781, 2.136416, 2.111562, 2.093903, 
    2.022484, 1.901195, 1.844082, 1.870107, 1.874339, 1.931435, 2.134218, 
    2.428164, 2.635537, 2.669765, 2.587978, 2.474176, 2.356273, 2.250999, 
    2.200788, 2.239427, 2.304108, 2.319896, 2.32307,
  1.857428, 1.887229, 1.903668, 1.860081, 1.716949, 1.563091, 1.513304, 
    1.566753, 1.635195, 1.697141, 1.80484, 1.886318, 1.916233, 1.944407, 
    1.990907, 2.041119, 2.114475, 2.144049, 2.047597, 1.93189, 1.956206, 
    2.053554, 2.145075, 2.302984, 2.478586, 2.573769, 2.572141, 2.479302, 
    2.353034, 2.288629, 2.32442, 2.358323, 2.331549, 2.364003, 2.466412, 
    2.499175, 2.440517, 2.381435, 2.42735, 2.526845, 2.634056, 2.708079, 
    2.729824, 2.767373, 2.795986, 2.707672, 2.530344, 2.34859, 2.199485, 
    2.138011, 2.224599, 2.405084, 2.574111, 2.665892, 2.787474, 2.95082, 
    3.132412, 3.305215, 3.335537, 3.227464, 3.149664, 3.149535, 3.169326, 
    3.183975, 3.261123, 3.34597, 3.338401, 3.294505, 3.255996, 3.208226, 
    3.147841, 3.015779, 2.738597, 2.308632, 1.897581, 1.557037, 1.278749, 
    1.07447, 1.025267, 1.091656, 1.19042, 1.172711, 1.127626, 1.19164, 
    1.410813, 1.658356, 1.81861, 1.890419, 1.935227, 2.000185, 2.020303, 
    1.968431, 1.920498, 1.918886, 1.893106, 1.846914,
  1.255571, 1.162392, 1.075722, 0.978261, 0.848443, 0.761838, 0.7523813, 
    0.7148819, 0.614769, 0.5714579, 0.5778551, 0.5649147, 0.5914125, 
    0.7148819, 0.8481827, 0.9534082, 1.108324, 1.267504, 1.268579, 1.191479, 
    1.216039, 1.263744, 1.223412, 1.23155, 1.353881, 1.462377, 1.493073, 
    1.415209, 1.231762, 1.106534, 1.10655, 1.110489, 1.086547, 1.105899, 
    1.140518, 1.172012, 1.169425, 1.113239, 1.075901, 1.145872, 1.244895, 
    1.239182, 1.180605, 1.173671, 1.201372, 1.199191, 1.162375, 1.1704, 
    1.238173, 1.211024, 1.107883, 1.110829, 1.211643, 1.322386, 1.433583, 
    1.483763, 1.476846, 1.571409, 1.746995, 1.825299, 1.874567, 2.033844, 
    2.181988, 2.228212, 2.236432, 2.199046, 2.187132, 2.247255, 2.328897, 
    2.264215, 2.120465, 1.890224, 1.568252, 1.330752, 1.201275, 0.9552956, 
    0.5900617, 0.4688048, 0.5412812, 0.6901259, 0.7733459, 0.7360735, 
    0.6697488, 0.6897192, 0.7755098, 0.8819227, 1.033567, 1.162521, 1.188775, 
    1.201307, 1.251096, 1.256077, 1.237197, 1.25899, 1.293592, 1.29662,
  0.655654, 0.7149143, 0.7016821, 0.5815163, 0.4203844, 0.2482977, 
    0.05062389, -0.1534615, -0.2843208, -0.3366318, -0.3786731, -0.4258733, 
    -0.422976, -0.3613062, -0.2705994, -0.1304789, 0.059268, 0.2321024, 
    0.3184471, 0.3910379, 0.5025787, 0.5891342, 0.5720119, 0.5758371, 
    0.668643, 0.727644, 0.7111893, 0.6332273, 0.4862537, 0.3261623, 
    0.2079983, 0.05798244, -0.09146404, -0.2191992, -0.401474, -0.5196543, 
    -0.462575, -0.4232349, -0.4679127, -0.4596605, -0.4087009, -0.4303474, 
    -0.5168715, -0.5856371, -0.5186138, -0.2980089, -0.2421494, -0.3435817, 
    -0.338438, -0.1199489, -0.01578188, -0.05370617, -0.03124428, 0.02087116, 
    0.115582, 0.2126846, 0.1985407, 0.2223363, 0.3465066, 0.4194884, 
    0.4233623, 0.4811587, 0.6219134, 0.7917218, 0.8978577, 0.8414779, 
    0.6896873, 0.6781149, 0.7654848, 0.7217021, 0.7226624, 0.7891011, 
    0.7409401, 0.7001033, 0.6617084, 0.3749251, 0.08607388, -0.03738022, 
    -0.3259544, -0.595046, -0.5313091, -0.4431257, -0.5235939, -0.5789981, 
    -0.5045033, -0.4461856, -0.3764429, -0.2841253, -0.195632, -0.141726, 
    -0.1228132, -0.06653118, 0.02995396, 0.1884823, 0.3962126, 0.5665255,
  -0.4184513, -0.3249784, -0.2394638, -0.2283964, -0.2754822, -0.3792744, 
    -0.5400329, -0.7108827, -0.8367128, -0.8742776, -0.8910909, -0.907155, 
    -0.9171162, -0.9205995, -0.9022403, -0.9056902, -0.9145613, -0.8162374, 
    -0.6759062, -0.5558209, -0.5094833, -0.5202088, -0.5068793, -0.4618602, 
    -0.3371363, -0.2129011, -0.1804638, -0.2486267, -0.4011822, -0.6013455, 
    -0.7689075, -0.9750104, -1.192622, -1.329422, -1.428022, -1.495795, 
    -1.589073, -1.761778, -1.80154, -1.730268, -1.77685, -1.88546, -1.857172, 
    -1.789171, -1.723644, -1.554519, -1.338487, -1.571315, -1.789887, 
    -1.639692, -1.502533, -1.637429, -1.691351, -1.648089, -1.505479, 
    -1.258099, -1.085231, -0.9893332, -0.9757752, -1.014398, -0.9959087, 
    -0.9593363, -0.9287376, -0.8388777, -0.7311625, -0.6140237, -0.5827575, 
    -0.5371847, -0.3855896, -0.3829365, -0.3438907, -0.2005472, -0.1310811, 
    -0.1860776, -0.3365173, -0.5977478, -0.6307228, -0.6777279, -1.09363, 
    -1.435019, -1.294655, -1.209092, -1.469883, -1.675091, -1.584694, 
    -1.407627, -1.337136, -1.285654, -1.190619, -1.080886, -1.028575, 
    -0.9512801, -0.843142, -0.7697372, -0.632628, -0.494998,
  -1.20849, -1.055935, -0.9549255, -0.9199324, -0.9729099, -1.015912, 
    -0.8958759, -0.7550232, -0.7960389, -0.7717388, -0.7137634, -0.8486266, 
    -1.228037, -1.576572, -1.74236, -1.971462, -2.104941, -1.978704, 
    -1.826181, -1.666937, -1.545274, -1.530609, -1.561322, -1.613112, 
    -1.57532, -1.419964, -1.401329, -1.456098, -1.506325, -1.698805, 
    -1.862201, -1.906487, -1.917604, -1.890017, -1.876003, -1.905153, 
    -1.993288, -2.061599, -1.940618, -1.702044, -1.767279, -1.916253, 
    -2.14433, -2.246495, -2.251784, -2.299115, -2.167702, -2.022796, 
    -2.383034, -2.578249, -2.578591, -2.681976, -2.638991, -2.54166, 
    -2.506944, -2.380593, -2.307302, -2.1289, -1.967312, -1.935898, 
    -1.850612, -1.856585, -1.822731, -1.723122, -1.718923, -1.600466, 
    -1.516302, -1.512217, -1.388242, -1.357204, -1.326475, -1.276328, 
    -1.298366, -1.268207, -1.338015, -1.309303, -0.9601495, -0.7529397, 
    -1.098187, -1.079372, -0.9807878, -1.178932, -1.325759, -1.43248, 
    -1.403704, -1.263958, -1.287836, -1.361354, -1.491514, -1.531504, 
    -1.503118, -1.487656, -1.420078, -1.443305, -1.460768, -1.340554,
  -1.754469, -1.633978, -1.549212, -1.456618, -1.431146, -1.455283, 
    -1.277484, -0.9269953, -0.7219826, -0.8232194, -1.102728, -1.333229, 
    -1.68362, -2.016578, -2.125059, -2.162689, -2.159027, -2.067002, 
    -2.058945, -2.077712, -2.080576, -2.065325, -1.949326, -1.996673, 
    -2.070713, -2.016107, -2.032367, -2.044183, -2.003102, -2.137819, 
    -2.195713, -2.106113, -1.892653, -1.562819, -1.562656, -1.810361, 
    -1.699961, -1.185736, -0.9584408, -1.090261, -1.016855, -1.173024, 
    -1.703346, -2.047292, -1.989626, -2.069085, -2.252337, -2.296657, 
    -2.528997, -2.66015, -2.478737, -2.42278, -2.330072, -2.296869, 
    -2.338503, -2.212184, -2.107236, -1.933522, -1.818272, -1.909206, 
    -1.912819, -2.052988, -2.137363, -2.024896, -2.015081, -1.875937, 
    -1.867897, -1.962477, -1.94415, -2.058245, -2.029909, -1.934043, 
    -1.89835, -1.706976, -1.559369, -1.144867, -0.4299576, -0.3034277, 
    -0.7004493, -0.7092227, -0.3901465, -0.424961, -0.3397559, -0.5332943, 
    -0.7132098, -0.7785743, -1.042832, -1.130772, -1.232285, -1.366774, 
    -1.388633, -1.555055, -1.622178, -1.630153, -1.735182, -1.799147,
  -1.543467, -1.513861, -1.375938, -1.034662, -0.5431745, -0.4069922, 
    -0.4508888, -0.4496517, -0.3175229, -0.4174418, -0.6814063, -0.9423275, 
    -1.050693, -1.215505, -1.296445, -1.348561, -1.530022, -1.668841, 
    -1.691937, -1.668353, -1.645436, -1.662429, -1.647406, -1.711046, 
    -1.904779, -1.940294, -1.868191, -1.809938, -1.696023, -1.505788, 
    -1.146087, -1.001996, -0.8176374, -0.6449649, -0.5752865, -0.6270443, 
    -0.6892514, -0.4647884, -0.4505146, -0.7232847, -0.6187109, -0.5966086, 
    -0.9433537, -1.216303, -1.409874, -1.651443, -1.86391, -1.922715, 
    -1.938357, -1.842654, -1.62086, -1.487348, -1.3942, -1.312689, -1.376507, 
    -1.322764, -1.34581, -1.385134, -1.362754, -1.496917, -1.433099, 
    -1.378119, -1.45429, -1.406048, -1.427467, -1.429079, -1.595029, 
    -1.771071, -1.75193, -1.827956, -1.800091, -1.793304, -1.751068, 
    -1.562982, -1.249213, -0.4956804, 0.1423731, 0.286188, -0.2601498, 
    -0.4562278, -0.1352962, -0.0889914, -0.1390078, -0.2700136, -0.5404723, 
    -0.4115014, -0.4543886, -0.5323505, -0.6856055, -0.8427019, -0.9263769, 
    -1.152549, -1.285524, -1.35307, -1.398675, -1.452549,
  -1.202614, -1.005691, -0.7297788, -0.2989516, 0.1239486, 0.2914779, 
    0.173558, -0.1244238, -0.3991637, -0.2438738, 0.0253644, -0.1639423, 
    -0.3064227, -0.3934021, -0.641921, -0.7214293, -0.7864037, -0.9294534, 
    -1.106276, -1.176508, -1.158376, -1.12545, -1.16347, -1.192295, 
    -1.224277, -1.13847, -1.015163, -0.8680596, -0.5948501, -0.3446064, 
    -0.3124611, -0.5181091, -0.3898048, -0.4010515, -0.3902116, -0.2088645, 
    -0.145843, -0.2375588, -0.4176047, -0.4798932, -0.3397074, -0.2991147, 
    -0.5039158, -0.5935478, -0.7426529, -0.9406347, -0.9008565, -0.8611426, 
    -0.7893171, -0.7171645, -0.5986261, -0.4344993, -0.4398375, -0.4591246, 
    -0.5698342, -0.6798115, -0.8447528, -0.983685, -0.8545351, -0.869916, 
    -0.9425397, -0.8584087, -0.8801047, -0.865033, -0.958132, -1.094802, 
    -1.16749, -1.28668, -1.2935, -1.359336, -1.318727, -1.236761, -1.011061, 
    -0.8119402, -0.5162535, -0.02927423, -0.01303059, 0.3676822, 0.1778547, 
    -0.3849707, 0.06584311, 0.1434797, -0.08161819, 0.07831025, -0.2352638, 
    -0.2675228, 0.06880522, 0.01825166, -0.1694272, -0.2016699, -0.3176858, 
    -0.497422, -0.7140074, -0.9958272, -1.177728, -1.222422,
  -0.5802178, -0.337347, -0.09193707, 0.1884177, 0.3448632, 0.178587, 
    0.06113911, -0.1935322, -0.2688251, 0.04720664, 0.4649801, 0.3125224, 
    0.3015847, 0.3136454, -0.1507092, -0.3274188, -0.4004822, -0.5284281, 
    -0.7800555, -0.9180603, -0.9917741, -0.9828711, -0.8230405, -0.6195254, 
    -0.5247822, -0.441514, -0.354291, -0.1807556, 0.2022195, 0.4855857, 
    0.3727438, -0.05754566, -0.1894631, -0.0839777, -0.2134862, -0.1975527, 
    -0.06587887, -0.1134539, -0.1707618, -0.2299578, -0.2494569, 
    0.0005106926, 0.2104554, 0.3005428, 0.39955, 0.08761978, -0.03508472, 
    0.2144918, 0.2817283, 0.2985091, 0.1972728, 0.2180085, 0.03014946, 
    -0.1983495, -0.4206967, -0.5507097, -0.4733658, -0.6063251, -0.7006772, 
    -0.6529231, -0.6953874, -0.6188903, -0.719785, -0.8842871, -0.9881284, 
    -1.070599, -0.9619403, -0.8994889, -0.8116803, -0.8309345, -0.7510676, 
    -0.6011653, -0.4376397, -0.1724057, 0.1323304, 0.2515688, -0.163291, 
    0.1501042, 0.2079493, -0.5762632, -0.03415692, 0.2625225, -0.1515237, 
    0.09766221, -0.1238217, -0.4102314, -0.1469665, -0.1507421, -0.2982521, 
    -0.2920184, -0.4486756, -0.4867454, -0.5573339, -0.6457458, -0.7659769, 
    -0.7840919,
  -0.09691763, 0.02442026, 0.2755437, 0.7072819, 0.8039615, 0.1141176, 
    0.0068748, -0.1166601, -0.2352149, 0.05485654, 0.3711488, 0.3214258, 
    0.1550684, 0.01512623, -0.1750586, -0.3418231, -0.3884053, -0.3412371, 
    -0.6962829, -1.007953, -1.031, -0.8892355, -0.6161556, -0.3392191, 
    -0.1303163, 0.05809498, 0.2468324, 0.3695865, 0.4618225, 0.5914452, 
    0.8894432, 1.032152, 0.8764389, 0.5697651, 0.3382549, 0.1887596, 
    0.07689452, 0.01926088, -0.1123471, -0.08598042, -0.1172466, 0.1016827, 
    0.8006897, 1.137441, 1.436008, 1.197809, 0.8790107, 1.137978, 1.010765, 
    0.9362211, 0.837327, 0.5835671, 0.1459208, -0.1396909, -0.1587987, 
    -0.2343197, -0.1777768, -0.3929133, -0.6851826, -0.7026792, -0.7465262, 
    -0.7331481, -0.710557, -0.7945738, -0.7612081, -0.6382093, -0.5211854, 
    -0.5079851, -0.4041114, -0.3390079, -0.2441998, -0.07628012, -0.02632761, 
    0.1951885, 0.3286359, 0.2775129, 0.209349, 0.2473855, 0.1264549, 
    -0.2117286, -0.224082, 0.1096749, -0.09154642, -0.01547265, 0.008160114, 
    -0.3595481, -0.1695738, -0.1684184, -0.3171973, -0.3227639, -0.3957462, 
    -0.3681412, -0.4530864, -0.3770123, -0.3365989, -0.2401304,
  0.05397749, 0.06646132, 0.1109602, 0.7106999, 1.072093, 0.2263575, 
    0.1651918, 0.2966535, 0.05298495, 0.0780499, 0.2205795, 0.4999088, 
    0.5215722, 0.7387595, 0.6618547, 0.1781964, -0.3971291, -0.3854103, 
    -0.4439878, -0.6935325, -0.7956805, -0.787087, -0.6677999, -0.3377376, 
    -0.01968765, 0.1838603, 0.3578188, 0.4403222, 0.6412823, 0.9026107, 
    1.176292, 1.541966, 1.665208, 1.054645, 0.7640524, 0.5116279, 0.1912336, 
    0.3307519, 0.2518783, 0.1150942, 0.149014, 0.4257715, 1.019131, 1.39068, 
    1.768366, 1.861074, 1.330915, 1.228425, 0.8820866, 0.5250065, 0.4690819, 
    0.3606346, -0.06667662, -0.4657977, -0.4108658, -0.2561951, -0.2233982, 
    -0.3805766, -0.5062113, -0.551621, -0.5853286, -0.6620708, -0.5999775, 
    -0.4837179, -0.3850036, -0.2662535, -0.1001244, 0.03374672, 0.02077436, 
    0.1002989, 0.07549429, 0.1163635, 0.2116604, 0.2579327, 0.3365297, 
    0.3129622, 0.3680892, 0.1972232, -0.04691744, -0.0281837, -0.1665788, 
    -0.05173528, -0.1046973, -0.02548194, -0.03596377, -0.4325624, 
    -0.2215106, -0.168972, -0.2694764, -0.1974382, -0.176312, -0.202126, 
    -0.1331482, -0.05212641, -0.02867222, 0.03827095,
  0.01917958, -0.01633465, -0.21736, 0.02012348, 0.56236, 0.5680564, 
    0.5570375, 0.5433497, 0.4068258, 0.3019757, 0.1748111, 0.4317123, 
    0.7776107, 1.194766, 0.9547917, 0.3877831, -0.324245, -0.6288021, 
    -0.3734313, -0.2123146, -0.1994569, -0.1971457, -0.2537215, -0.032318, 
    0.2520406, 0.4936914, 0.6874252, 0.7094792, 0.7619041, 0.8218652, 
    0.8262272, 0.7472885, 0.7624414, 0.6307352, 0.7941303, 0.6007876, 
    0.2817123, 0.2013737, 0.2119369, -0.04681993, -0.04231125, 0.1957097, 
    0.1938054, 0.4676336, 0.7656478, 0.8243717, 0.2737207, 0.07419273, 
    -0.174082, -0.4983496, -0.5860943, -0.382497, -0.3012636, -0.6182551, 
    -0.7724383, -0.5548277, -0.3240495, -0.1962829, 0.005654335, -0.01957369, 
    -0.1377058, -0.1407981, -0.1458597, -0.03314829, 0.1474185, 0.2617903, 
    0.2342019, 0.2832904, 0.2595601, 0.3719788, 0.3555398, 0.2910709, 
    0.3017478, 0.1558332, 0.268968, 0.2275781, 0.07572269, -0.02805335, 
    -0.04330409, 0.01135096, -0.0132747, -0.07185233, -0.1775814, 0.0135479, 
    -0.0523864, -0.3111591, -0.1057229, 0.09995747, 0.1545477, 0.1857486, 
    0.2561588, 0.1927967, 0.1786032, 0.1159892, 0.08423471, 0.03625321,
  0.08327472, -0.0498144, -0.01939464, 0.1261778, 0.3100652, 0.4715234, 
    0.5409245, 0.6766829, 0.7997462, 0.6209863, 0.2592839, 0.1279199, 
    -0.04966793, 0.02886397, -0.08959311, -0.09953785, -0.1386004, 
    -0.2901954, -0.2213966, -0.0939225, -0.03025067, -0.073138, -0.2444433, 
    -0.1762956, -0.04607117, 0.05514979, 0.06330383, 0.01989555, 0.1929584, 
    -0.02862358, -0.1641214, -0.1797464, -0.001669884, 0.1325747, 0.3180401, 
    0.2587304, 0.2648501, -0.114219, 0.1077864, 0.1460026, -0.1788672, 
    -0.3597754, -0.9616637, -0.8557554, -0.4880469, -0.3614843, -0.519248, 
    -0.7134863, -1.021852, -1.025693, -0.7102474, -0.5029886, -0.1893167, 
    -0.162396, -0.3792582, -0.4447691, -0.3525164, -0.285573, -0.1042743, 
    0.05497074, 0.07822943, 0.1528711, 0.193284, 0.1612368, 0.1692448, 
    0.3448305, 0.4291563, 0.4105201, 0.420661, 0.3600321, 0.2896547, 
    0.181061, 0.1017315, 0.06359673, 0.04605147, 0.1309471, 0.0351465, 
    -0.06724614, -0.008277968, -0.01752275, -0.007252753, -0.0768978, 
    -0.1372331, -0.2347429, -0.469769, -0.2383075, -0.1913996, -0.03412461, 
    0.09717417, 0.1215231, 0.2865622, 0.2545149, 0.2252667, 0.2794821, 
    0.2956283, 0.1561098,
  0.339134, 0.1845931, 0.1446513, 0.4180074, 0.6282127, 0.1736393, 0.1180079, 
    0.498086, 0.9986556, 1.061383, 0.744684, 0.2795632, -0.1658466, 
    -0.1592545, -0.08233404, -0.03607762, -0.199424, -0.4063576, -0.4231384, 
    -0.3803486, -0.4798601, -0.5873631, -0.7260023, -0.7306085, -0.7491145, 
    -0.7599545, -0.716172, -0.6707621, -0.2263771, -0.2851824, -0.5685807, 
    -0.6737403, -0.2456642, -0.005706549, 0.08296537, -0.05655289, 
    -0.09675491, -0.2438086, -0.01340491, 0.02253259, -0.5106057, -0.7136166, 
    -1.136452, -1.131748, -0.9564714, -0.8111914, -0.8198503, -0.9430436, 
    -1.145225, -1.186826, -0.8533633, -0.7284608, -0.4286883, -0.2129006, 
    -0.1901305, -0.08949566, 0.05466127, 0.1526594, 0.1978903, 0.224632, 
    0.2887759, 0.3434632, 0.3988669, 0.4544497, 0.4700911, 0.4938865, 
    0.5464256, 0.5030336, 0.5558331, 0.4940329, 0.4595444, 0.3138082, 
    0.1158594, 0.1081282, -0.1622656, 0.09292632, 0.1231022, -0.007529259, 
    0.009576857, 0.05495429, 0.05381513, -0.04699874, 0.008404791, 
    -0.07723957, -0.4592057, -0.3697852, -0.3163347, -0.3624616, -0.09953773, 
    0.01942384, 0.07315111, 0.1669662, 0.2915429, 0.4263412, 0.4458399, 
    0.3302474,
  0.2789614, 0.3015194, 0.1338117, 0.3239486, 0.3436261, 0.01449203, 
    -0.007659473, 0.04279625, 0.3741114, 1.103717, 1.215697, 0.1420474, 
    0.02293921, 0.1576717, 0.2004297, 0.2384342, -0.0613053, -0.3256119, 
    -0.5064551, -0.6252864, -0.7001566, -0.7806414, -0.9067156, -0.8632096, 
    -0.720078, -0.7003189, -0.5314548, -0.165179, -0.1365494, -0.1819599, 
    -0.08851904, -0.1724056, -0.03791662, 0.170091, 0.1992253, 0.001438841, 
    -0.09206702, -0.1080338, -0.2487077, -0.4248959, -0.676263, -0.7441179, 
    -0.9667096, -0.8568463, -0.8691831, -0.9193132, -0.9962502, -1.066498, 
    -1.062331, -1.136924, -0.971283, -0.9440694, -0.8174419, -0.6087179, 
    -0.4467216, -0.1805921, 0.03451157, 0.2521224, 0.4537988, 0.5492411, 
    0.660049, 0.7507713, 0.8445702, 0.8651435, 0.8823147, 0.8495015, 
    0.7917054, 0.7178288, 0.6587467, 0.5412826, 0.5022364, 0.4815819, 
    0.3334697, 0.1867249, -0.1788838, 0.1066959, 0.1686426, 0.05487309, 
    -0.0001887679, 0.1449121, 0.1036196, 0.05728185, 0.03887367, -0.09271812, 
    -0.2979269, -0.3528094, -0.2302508, -0.1743751, 0.01330408, 0.00690759, 
    -0.05009115, 0.1107975, 0.0780338, 0.1513247, 0.242975, 0.2910702,
  0.0694561, 0.2183983, 0.2012596, 0.2507715, 0.1319889, 0.03996414, 
    0.033877, 0.0153223, 0.2506412, 1.075299, 1.651634, 0.2158267, 
    0.06916332, 0.2855048, 0.3766336, 0.3473206, 0.1701887, 0.03596032, 
    -0.2756608, -0.437054, -0.5913509, -0.7804459, -0.802386, -0.7849543, 
    -0.5359963, -0.319216, -0.316514, -0.2182227, -0.441237, -0.3438736, 
    -0.1853287, -0.01906897, -0.02032232, 0.06804013, 0.0857811, -0.08607769, 
    -0.1706316, -0.192409, -0.2709739, -0.3177676, -0.3126564, -0.3478289, 
    -0.4869399, -0.3590107, -0.2592874, -0.2690039, -0.2519956, -0.3100362, 
    -0.3877707, -0.3811789, -0.3384218, -0.3545189, -0.3776145, -0.3989358, 
    -0.3780212, -0.3112082, -0.07691431, 0.08882427, 0.2300196, 0.3621488, 
    0.4736714, 0.5248919, 0.5750718, 0.6547427, 0.7702863, 0.8248926, 
    0.760716, 0.6995345, 0.6359115, 0.6299381, 0.5045311, 0.4689356, 
    0.2419333, -0.1695898, -0.5134537, -0.1790625, 0.09631189, 0.2308333, 
    0.1158431, 0.2700422, 0.07772422, -0.05598325, -0.2658958, -0.2314715, 
    -0.2797303, -0.1743913, 0.08242846, 0.1310284, 0.1905172, 0.1382227, 
    0.1433659, 0.1262758, -0.03467822, 0.06060219, -0.1182554, -0.008879662,
  0.08436525, 0.01265275, 0.1308171, 0.2091699, 0.2084863, -0.04608738, 
    0.00912115, 0.2669497, 0.3196678, 0.584821, 1.060765, 0.486546, 
    -0.01430082, 0.08374643, 0.3592186, 0.2374413, 0.1150129, -0.1012793, 
    -0.224668, -0.3815691, -0.8173601, -0.8029884, -0.5364681, -0.6846777, 
    -0.5387467, -0.2291438, -0.1501887, -0.319948, -0.5845642, -0.6887302, 
    -0.4962668, -0.1410416, 0.1092029, -0.05520201, 0.07494116, 0.03617191, 
    0.1009827, 0.06493139, -0.05912399, -0.06358433, -0.1016865, -0.2040467, 
    -0.1943297, -0.1609635, -0.08397865, -0.0908637, -0.08375072, 0.04064703, 
    0.04137945, 0.002984047, -0.1112247, -0.1373806, -0.1568627, -0.2787867, 
    -0.1920519, -0.1844506, -0.09024525, -0.04052114, -0.0319767, 
    -0.04732466, 0.08377886, 0.2270894, 0.2431378, 0.3849835, 0.5021224, 
    0.5546286, 0.6464095, 0.6753483, 0.5349833, 0.4158753, 0.1066632, 
    0.1400129, 0.1397037, -0.1059181, -0.2408631, 0.02660158, 0.3702703, 
    0.4461324, 0.4885478, 0.02481079, -0.1518166, -0.2406023, -0.2087507, 
    -0.1378036, -0.07304049, -0.04537153, -0.0128355, 0.06330347, 0.1414127, 
    0.2660869, 0.3425847, 0.2646224, 0.2373924, 0.3236556, 0.09969723, 
    0.1020408,
  0.1364812, 0.2740136, 0.4373274, 0.4763249, 0.2531315, 0.03347009, 
    0.1917869, 0.3673894, 0.4028711, 0.3916081, 0.3839258, 0.2120831, 
    -0.01363301, -0.055902, 0.2277246, 0.316494, 0.412132, 0.1702213, 
    0.129873, -0.2380632, -0.3608661, -0.1228938, -0.2544377, -0.5472429, 
    -0.6110123, -0.9316019, -1.24931, -0.7333601, -0.6330996, -0.7410259, 
    -0.5078878, -0.2813735, -0.1292255, -0.04877305, 0.12468, 0.04927397, 
    0.1179585, 0.1143293, 0.08110905, -0.000287056, -0.02919388, -0.2332301, 
    -0.235558, -0.1401472, -0.1197367, -0.07818413, -0.04800797, 
    -0.006520271, -0.05175018, -0.1107187, -0.09431267, -0.1725035, 
    -0.1810493, -0.2446232, -0.2169218, -0.08825874, -0.06638432, 
    0.005865097, 0.1330462, 0.1522522, 0.2232642, 0.3167052, 0.3777237, 
    0.4895082, 0.4906473, 0.4988832, 0.5619206, 0.5583723, 0.4855859, 
    0.4179263, 0.1860905, 0.07370424, -0.1008883, -0.256927, 0.0001367629, 
    0.2155502, 0.1772363, 0.2927799, 0.2380271, -0.1338315, -0.07149506, 
    -0.0422802, -0.2207136, 0.01056862, -0.02823353, -0.07313919, 
    -0.01814175, 0.08752251, 0.07212496, 0.2242088, 0.2497296, 0.4415593, 
    0.6145082, 0.4894271, 0.3025293, 0.3071192,
  0.3397853, 0.4558493, 0.4512928, 0.2175844, -0.005707026, -0.04431319, 
    0.1432843, 0.08159804, 0.267373, 0.4071517, 0.1774313, 0.0110091, 
    -0.08580112, 0.02604795, 0.1943426, 0.3265042, 0.3516178, 0.2485905, 
    0.3509831, 0.149795, 0.3055723, -0.2129986, -0.410476, -0.6828711, 
    -0.9315529, -0.8503678, -0.8951436, -0.2798763, -0.3980567, -0.4935489, 
    -0.2588806, -0.301784, -0.2447524, -0.1240826, -0.1421814, -0.1210384, 
    -0.0411725, -0.05756235, 0.05327702, -0.02593851, -0.01107836, 
    -0.1251087, -0.1825304, -0.1791124, -0.1143179, -0.03501987, 0.02370453, 
    0.0234766, 0.07718849, -0.0462656, -0.1270599, -0.2052174, -0.2306566, 
    -0.2332621, -0.2806578, -0.1464777, -0.1088963, 0.04186821, 0.1631899, 
    0.2649307, 0.3534398, 0.3863664, 0.4484267, 0.4315329, 0.4204812, 
    0.4268131, 0.3035057, 0.3421775, 0.6241763, 0.8107486, 1.054498, 
    0.9668519, 0.1933167, -0.1151304, 0.3465223, 0.5116282, 0.5660553, 
    0.596508, 0.2759504, -0.05871677, -0.07144547, -0.05364037, -0.01882601, 
    -0.01889133, -0.1949162, -0.1216741, -0.1344509, -0.1129336, -0.06788158, 
    0.1041403, 0.1951072, 0.4431706, 0.3877018, 0.114557, 0.1020246, 0.2634665,
  0.3899965, 0.2806542, 0.1101301, -0.07854247, -0.1394143, -0.1113381, 
    -0.08034801, -0.02681661, 0.1899153, 0.1292057, 0.1410871, -0.06005204, 
    -0.2007589, 0.02292299, 0.1834698, 0.1877503, 0.202106, 0.3952048, 
    0.3990299, 0.4038477, 0.2351626, -0.5268008, -0.3105404, -0.4453382, 
    -0.4525162, -0.3514748, -0.3406514, -0.7736914, -0.7856706, -0.266937, 
    -0.509336, -0.4827411, -0.38834, -0.3449802, -0.3850851, -0.3390241, 
    -0.2345967, -0.1651306, -0.1052351, -0.1714616, -0.23528, -0.3074808, 
    -0.3468366, -0.4143014, -0.2320423, -0.2009058, -0.1118431, -0.1105566, 
    -0.04641342, -0.04808903, -0.1308699, -0.2176371, -0.401639, -0.4413843, 
    -0.4473248, -0.3860788, -0.3754501, -0.2255478, -0.1081648, 0.01427937, 
    0.07640553, 0.195611, 0.2348361, 0.2320375, 0.2968001, 0.2230856, 
    0.2362691, 0.4229883, 0.4645572, 0.1574772, 0.13194, 0.1550357, 
    -0.3075947, -0.06651402, 0.4636779, 0.6679258, 0.6677637, 0.2523184, 
    -0.1643333, -0.08087015, -0.06688881, -0.1636009, -0.2683702, -0.4363227, 
    -0.462738, -0.4289498, -0.4899359, -0.4025164, -0.3144469, -0.1907001, 
    0.004401207, 0.1988344, -0.04047203, -0.01501656, 0.1585677, 0.350446,
  0.2741601, 0.1659732, 0.01471996, -0.0788672, -0.2192645, -0.3338313, 
    -0.3446393, -0.2603619, -0.09838223, -0.1046649, 0.2227601, 0.01410145, 
    -0.3646746, -0.1011494, 0.08841801, -0.1458595, -0.1867452, 0.05591473, 
    -0.3631608, -0.3482845, -0.1433366, -0.3194433, -0.2910254, -0.5029397, 
    -0.3606057, -0.2684176, -0.3051855, -0.3734798, -0.4672625, -0.2393818, 
    -0.6574807, -1.06264, -1.149798, -0.8672137, -0.5497823, -0.4893165, 
    -0.459857, -0.4297624, -0.5005145, -0.5727477, -0.5972762, -0.6584249, 
    -0.6602478, -0.6530538, -0.5680113, -0.6879334, -0.5691504, -0.4876242, 
    -0.475482, -0.4202094, -0.5085878, -0.6264429, -0.6303811, -0.5179462, 
    -0.6417909, -0.6632428, -0.5004339, -0.3789334, -0.2643003, -0.0941186, 
    -0.05082417, 0.04735327, 0.03721333, 0.07230473, 0.1627831, 0.168349, 
    0.4961003, 0.6296127, 0.4177963, -0.07396811, -0.1988869, -0.06153321, 
    -0.4378521, -0.2894301, -0.1568623, -0.1189222, -0.01207066, -0.03449917, 
    0.003961563, -0.2068949, -0.5966568, -0.6980572, -0.8219175, -0.9258404, 
    -1.079323, -1.247747, -1.106879, -1.016254, -0.9621525, -0.7154722, 
    -0.5042906, -0.2118263, -0.1185484, -0.07608414, 0.06805658, 0.2510643,
  0.05449867, -0.08218777, -0.1921161, -0.2531348, -0.4423275, -0.4236914, 
    -0.4174253, -0.6121029, -0.2434668, -0.08034843, -0.3552507, -0.5935318, 
    -0.5025489, 0.04992515, 0.2854883, -0.2552343, -0.3417089, -0.1557066, 
    -0.4575132, -0.2895769, -0.1938088, -0.4304788, -0.6813411, -0.7554293, 
    -0.1599383, -0.1789812, 0.187132, -0.6276956, -1.093207, -0.3036882, 
    -0.4972755, -0.5760031, -0.3929137, -0.5251243, -0.5976827, -0.6441338, 
    -0.6111588, -0.6646258, -0.7309505, -0.8592218, -0.9245219, -0.9407001, 
    -0.8766706, -0.7826765, -0.7637305, -0.8767838, -0.9011817, -0.8787045, 
    -0.7951431, -0.7503676, -0.7903743, -0.8959732, -0.9708757, -0.9626076, 
    -0.9579525, -0.8372169, -0.6705666, -0.4708924, -0.2725358, -0.1349869, 
    -0.04457331, 0.08729506, 0.09598613, 0.04665351, 0.07186496, 0.2012759, 
    0.3481998, 0.2943913, 0.186237, 0.003245413, -0.1576597, -0.2810971, 
    -0.4358823, -0.2674253, -0.1860449, -0.1662207, -0.1508238, -0.2740984, 
    -0.469281, -0.8588808, -1.032627, -1.151638, -1.415749, -1.556781, 
    -1.691791, -1.661094, -1.493044, -1.541497, -1.393174, -1.02042, 
    -0.8615003, -0.496592, -0.1089129, 0.05360317, 0.1664939, 0.1678612,
  -0.09117186, -0.07876956, -0.1165137, -0.1763281, -0.4313248, -0.3177018, 
    -0.4136329, -0.7333595, -0.3170996, -0.177549, -0.7546973, -0.7069433, 
    -0.124261, 0.3054916, 0.07471353, -0.3862404, -0.1873958, -0.07056659, 
    -0.178542, 0.06463873, -0.00292325, -0.4410905, -0.5476822, -0.2338316, 
    0.05456352, 0.4994043, 0.2123433, -1.322129, -0.7419212, 0.08822274, 
    -0.2598243, -0.1211036, -0.2440692, -0.415586, -0.5513445, -0.7598242, 
    -0.7134213, -0.7743753, -0.9152607, -0.9814879, -0.9453877, -1.023008, 
    -1.091302, -1.03585, -0.9725847, -0.8778581, -0.7964454, -0.8122819, 
    -0.8354102, -0.8949316, -0.930023, -1.007529, -1.141693, -1.225889, 
    -1.196413, -1.059889, -0.9133399, -0.5545346, -0.274196, -0.1505144, 
    0.004596353, 0.08200526, 0.1349185, 0.1474186, 0.1750391, 0.2215879, 
    0.1976789, 0.09133142, 0.1559636, -0.1835384, -0.5610937, -0.6319108, 
    -0.5008237, -0.2258235, -0.1976334, -0.4059505, -0.6502539, -0.8919369, 
    -1.176393, -1.345729, -1.33974, -1.50901, -1.683636, -1.811989, 
    -1.908782, -1.821917, -1.810801, -1.635752, -1.300612, -1.031911, 
    -0.6601825, -0.2823668, -0.07640982, 0.1396222, 0.3135157, 0.08239567,
  0.2824119, 0.3219139, 0.1923242, 0.05217111, -0.236696, -0.3845638, 
    -0.4941183, -0.7678811, -0.689056, -0.5596455, -0.438861, 0.08872718, 
    0.3502832, -0.06001949, -0.5848408, -0.6014095, -0.3796647, -0.3510517, 
    -0.2364359, 0.2276756, 0.3383362, 0.4058163, 0.2764225, 0.06707954, 
    0.1387267, 0.3710842, -0.3005476, -0.4401957, 0.3579001, 0.1932518, 
    -0.2320088, 0.1335022, 0.1606997, 0.2890527, 0.2749089, -0.1126562, 
    -0.1769143, -0.2764909, -0.469053, -0.5647886, -0.5577247, -0.587168, 
    -0.6781838, -0.69542, -0.7365496, -0.7232847, -0.6002214, -0.4797301, 
    -0.461875, -0.5685806, -0.7482356, -0.988942, -1.056715, -1.06609, 
    -1.148414, -1.098919, -0.9191672, -0.6470636, -0.4233335, -0.1137958, 
    0.203945, 0.2606183, 0.3310286, 0.3228254, 0.2885807, 0.350999, 
    0.2937077, 0.3405664, 0.2925196, -0.1216731, -0.3247982, -0.2209082, 
    -0.1290625, -0.1529559, -0.2488868, -0.507432, -0.6714458, -0.7387142, 
    -0.9571226, -1.243288, -1.443809, -1.536761, -1.493467, -1.635199, 
    -1.766188, -1.654974, -1.543353, -1.249587, -0.9063576, -0.6028417, 
    -0.03469397, 0.398981, 0.4118392, 0.4246158, 0.3943424, 0.2827539,
  0.5360575, 0.3660867, 0.1478252, 0.07028627, -0.1625261, -0.4123309, 
    -0.4504657, -0.4484799, -0.4172137, -0.1847429, 0.236416, 0.2052799, 
    -0.2736589, -0.6376078, -0.5848405, -0.4031347, -0.42667, -0.4615495, 
    -0.2474544, 0.1644597, 0.6232483, 0.5949123, 0.102529, 0.1251526, 
    0.115273, -0.2306092, -0.1126726, 0.2566146, 0.3455791, 0.2366765, 
    0.3152083, 0.4605534, 0.367015, 0.643903, 0.6034408, 0.4271054, 
    0.2057357, 0.05599594, 0.2229557, 0.3483629, 0.2173886, 0.1431866, 
    0.009022713, -0.131309, -0.1442647, -0.07483101, -0.1209249, -0.2432394, 
    -0.3219337, -0.3742776, -0.4171162, -0.55128, -0.6808534, -0.7116475, 
    -0.6625748, -0.4920015, -0.3433042, -0.1510196, 0.09852552, 0.3035219, 
    0.3625226, 0.4242251, 0.473639, 0.2728903, 0.2187891, 0.3403711, 
    0.3022038, 0.3424057, 0.4060774, 0.2617252, 0.1892642, 0.1984439, 
    0.1444727, 0.0542382, 0.02803385, 0.02113271, -0.05962896, -0.2867937, 
    -0.6120543, -0.7651954, -0.7512956, -0.9493265, -1.278298, -1.542458, 
    -1.524359, -1.252467, -0.9541113, -0.6936135, -0.299082, 0.2493553, 
    0.6775613, 0.7537659, 0.7615299, 0.87123, 0.8820376, 0.6741276,
  0.540257, 0.4156966, 0.2043357, 0.02531576, -0.1208107, -0.07440782, 
    0.1674057, 0.2910873, 0.1782292, 0.2103906, 0.295791, 0.0276432, -0.3907, 
    -0.2165625, 0.1099024, 0.2197657, 0.3479069, 0.07155597, -0.222666, 
    0.1985904, 0.7297262, 0.4936263, 0.1417221, 0.3029525, 0.5706608, 
    0.2268457, 0.7414778, 0.9577051, 0.7128156, 0.7404197, 0.7763574, 
    0.3600489, 0.2538312, 0.3802474, 0.4153709, 0.603457, 0.5946679, 
    0.447093, 0.5888567, 0.7853088, 0.6809311, 0.5124898, 0.3239317, 
    0.2152085, 0.2160378, 0.2018938, 0.1287661, 0.02072573, 0.003993511, 
    0.01554918, -0.1180773, -0.2391057, -0.2097759, -0.1468043, 0.009169102, 
    0.2372127, 0.3871479, 0.4949117, 0.5785866, 0.5427957, 0.5083556, 
    0.5937397, 0.4373106, 0.1186426, 0.2501693, 0.4168522, 0.3613346, 
    0.5715878, 0.7029686, 0.4954653, 0.1572331, 0.1073632, 0.165485, 
    0.1201885, 0.02389908, 0.008078814, -0.06762052, -0.1172791, -0.155283, 
    -0.210557, -0.3000264, -0.4718194, -0.604486, -0.6148858, -0.5655699, 
    -0.388031, -0.1307225, 0.1040425, 0.4475322, 0.9317935, 1.16542, 
    1.087425, 1.064134, 1.012181, 0.8069237, 0.6600809,
  0.3134017, 0.1573143, -0.05352497, -0.1026141, -0.03863277, 0.03221682, 
    0.1247299, 0.1699121, 0.1992903, 0.307933, 0.2258529, 0.1242741, 
    -0.02051754, 0.1865461, 0.529824, 0.6834698, 0.8315166, 0.5619206, 
    0.3050847, 0.3444564, 0.5568587, 0.4494043, 0.6268457, 0.9488673, 
    0.365013, -0.002402306, 0.8134177, 1.143333, 0.6513084, 0.4724669, 
    0.4485576, 0.4054096, 0.5274477, 0.394619, 0.160358, 0.353164, 0.8001361, 
    0.8984599, 1.014068, 0.888711, 0.8679914, 0.6917548, 0.4764872, 
    0.4983788, 0.4538965, 0.2226787, 0.07088852, -0.04771519, -0.1968203, 
    -0.2754016, -0.2937441, -0.2423282, -0.08500433, 0.03355026, 0.2298889, 
    0.6035867, 0.830719, 0.8703022, 0.8353906, 0.7445049, 0.6470118, 
    0.4694238, 0.2796128, 0.2562077, 0.6252669, 0.6383691, 0.3862041, 
    0.3843975, 0.3866436, 0.05197597, -0.2101175, -0.09711289, 0.01149738, 
    0.0370506, 0.05929995, 0.09222651, 0.02036715, 0.06388974, 0.08216786, 
    0.0895896, 0.1397686, 0.3202863, 0.4548402, 0.462018, 0.5705953, 
    0.8248434, 0.999176, 0.9973698, 1.080557, 1.264069, 1.222451, 1.132168, 
    1.149909, 1.013678, 0.7049708, 0.5132062,
  0.03127253, -0.07193363, -0.143532, -0.2363216, -0.3224055, -0.3167416, 
    -0.3294532, -0.267181, -0.1077083, 0.02385095, 0.1046289, 0.1120834, 
    0.2093002, 0.4385484, 0.8488181, 0.8790427, 0.7495668, 0.7241927, 
    0.8176658, 0.8636618, 0.7184147, 0.420612, 0.3704818, 0.3551172, 
    0.05650061, 0.1640689, 0.5566635, 0.7277573, 0.4480371, 0.382656, 
    0.4516503, 0.444098, 0.3458235, 0.2287986, 0.1831932, 0.3981998, 
    0.5656149, 0.8880923, 1.101259, 1.236155, 1.292991, 1.163678, 1.079238, 
    1.136953, 1.037637, 0.8327699, 0.8058338, 0.7167544, 0.3878317, 
    0.1762433, 0.2572002, 0.4274154, 0.5037007, 0.4781961, 0.5739808, 
    0.7481675, 0.7365456, 0.6133528, 0.6340234, 0.7473371, 0.7312562, 
    0.573395, 0.4412337, 0.3987207, 0.3676172, 0.3722233, 0.2915103, 
    0.1856995, -0.04940748, -0.1326923, -0.1367774, -0.0441016, -0.03264332, 
    0.06486642, -0.04512715, -0.06047529, -0.09821939, -0.06609082, 
    0.1062565, 0.3925354, 0.492568, 0.7860091, 1.050364, 1.177708, 1.334414, 
    1.439231, 1.361058, 1.242503, 1.265794, 1.399665, 1.347044, 1.205638, 
    1.050283, 0.7858138, 0.4294822, 0.1627181,
  -0.2948178, -0.2632424, -0.3930111, -0.6187761, -0.8512468, -0.7868916, 
    -0.5916276, -0.3710221, -0.1052506, -0.1382422, -0.2178972, -0.113291, 
    0.1553776, 0.4024642, 0.6188216, 0.6716537, 0.6098047, 0.5558334, 
    0.6300196, 0.7119369, 0.6860743, 0.5276758, 0.3480534, 0.2972069, 
    0.42748, 0.6226459, 0.6756248, 0.4250226, 0.2681053, 0.2496481, 
    0.1789939, 0.001764297, -0.1328876, 0.008860588, 0.2496319, 0.2643945, 
    0.1641501, 0.5068425, 1.025364, 2.038987, 1.850641, 1.790305, 2.060293, 
    2.357249, 2.214215, 1.796002, 1.400852, 1.088743, 0.8767147, 0.9007063, 
    1.073118, 1.213369, 1.248834, 1.263271, 1.323949, 1.288922, 1.040599, 
    0.7662497, 0.6724837, 0.674567, 0.6296287, 0.4920801, 0.2392806, 
    0.05871403, 0.03174484, 0.05405903, 0.08599281, -0.2081642, -0.3044374, 
    -0.1857519, -0.1523212, -0.1257259, -0.03449866, -0.03174818, -0.1455339, 
    -0.2029884, -0.1433204, -0.07191741, -0.006699383, 0.103164, 0.3294987, 
    0.4227766, 0.8875389, 1.071881, 1.296816, 1.451862, 1.507379, 1.510114, 
    1.473997, 1.398965, 1.318187, 1.083942, 0.6329002, 0.1723371, -0.1548433, 
    -0.284466,
  -0.9759539, -1.049033, -0.8685481, -0.7436296, -0.6490333, -0.5483986, 
    -0.3634539, -0.04556638, 0.1185775, 0.1009831, -0.01150062, 0.03111006, 
    0.1620508, 0.2476465, 0.3426172, 0.3634993, 0.38194, 0.376048, 0.3693261, 
    0.380654, 0.3714906, 0.3521061, 0.3096744, 0.2968487, 0.2409242, 
    0.1058818, 0.01649392, 0.04338193, 0.008372068, -0.1249124, -0.2035089, 
    -0.09525752, 0.01024389, 0.0712142, 0.1904522, 0.3279521, 0.5572493, 
    1.000104, 1.192486, 1.333291, 0.8791894, 0.7305241, 1.07766, 1.741885, 
    1.947565, 1.942536, 1.88736, 1.879173, 1.881582, 1.864687, 1.70069, 
    1.367308, 1.031696, 0.842845, 0.7945051, 0.8016503, 0.7275944, 0.7655338, 
    0.852806, 0.8807683, 0.7452862, 0.323346, 0.1131575, 0.03913415, 
    0.06405258, 0.02837563, -0.04779649, -0.0754981, -0.0301857, 0.05189457, 
    0.06058598, 0.07018884, 0.1615463, 0.28111, 0.231354, 0.0797264, 
    0.09178713, -0.0104264, -0.1091571, -0.008001328, 0.09826493, 0.138418, 
    0.1556705, 0.3909732, 0.872272, 1.265013, 1.46402, 1.432559, 1.322093, 
    1.254319, 1.124094, 0.7864323, 0.2392807, -0.2316505, -0.516807, 
    -0.7894144,
  -1.385541, -1.207074, -0.8696387, -0.5353613, -0.4518815, -0.4845149, 
    -0.1773535, -0.1765397, -0.04904944, -0.02426103, -0.0347428, 0.04484706, 
    0.1808334, 0.2744532, 0.2863672, 0.2593164, 0.2318097, 0.2022525, 
    0.1142969, 0.1086491, 0.003180385, -0.09546912, -0.07684946, -0.06918335, 
    -0.1607685, -0.303249, -0.3074481, -0.1861917, -0.1943457, -0.2706155, 
    -0.2309833, -0.01260757, 0.02329683, 0.03675747, 0.1945374, 0.5792053, 
    0.8631245, 0.8356836, 0.5583886, -0.07465172, -0.5389261, -0.1156187, 
    0.4493715, 0.5643779, 0.6244364, 1.244505, 1.619473, 1.954955, 2.172012, 
    1.87141, 1.322923, 0.7742248, 0.41013, 0.204417, 0.115973, 0.3030987, 
    0.4102927, 0.5681055, 0.6456118, 0.5937889, 0.1590722, 0.186123, 
    0.1014388, 0.05226886, 0.02647132, -0.07250321, -0.1577897, -0.1058365, 
    0.03636724, 0.1306055, 0.1270736, 0.149209, 0.1803286, 0.1885806, 
    0.1015851, 0.02658516, -0.1312761, -0.2654721, -0.2085875, -0.01166368, 
    0.1537172, 0.2382878, 0.07134426, 0.2192611, 0.4589096, 0.5511296, 
    0.418545, 0.2853093, 0.2207584, 0.1467838, -0.02925795, -0.3507586, 
    -0.7008725, -0.9596454, -1.143793, -1.270371,
  -1.02833, -0.7313411, -0.3525651, -0.3182552, -0.3622331, -0.2689062, 
    -0.2780696, -0.1284765, 0.01745447, 0.09509119, 0.1104883, 0.1246648, 
    0.153099, 0.1830469, 0.2266504, 0.2124252, 0.1095443, -0.001474738, 
    -0.1426532, -0.2448665, -0.3399349, -0.415472, -0.4495052, -0.4228126, 
    -0.3892838, -0.3906836, -0.3214291, -0.2448177, -0.1856544, -0.1069274, 
    0.04056597, 0.1840234, 0.2183168, 0.2569236, 0.3845929, 0.5174055, 
    0.4123436, 0.1256413, -0.1738056, -0.2860289, -0.08484054, 0.1989322, 
    0.2534244, 0.1426008, 0.09870434, 0.1540592, 0.1892641, -0.1809995, 
    -0.6245544, -0.8321388, -0.82903, -0.7801697, -0.3754985, -0.3066019, 
    -0.1705015, -0.04094434, 0.08431613, 0.2060285, 0.1640687, 0.09367514, 
    0.04670233, -0.009287071, -0.01366535, -0.003362566, -0.04048824, 
    -0.06768566, 0.008697927, 0.1567121, 0.2581934, 0.2747136, 0.268252, 
    0.2153874, 0.1266016, -0.02269852, -0.1535091, -0.1583105, -0.1801692, 
    -0.04193681, 0.1017155, 0.2817936, 0.3987858, 0.4882878, 0.3981837, 
    0.3057519, 0.09284496, -0.2155696, -0.5001563, -0.4990332, -0.4823502, 
    -0.5726662, -0.8236427, -1.095176, -1.252288, -1.298659, -1.291042, 
    -1.224066,
  -0.6637957, -0.5304297, -0.3712826, -0.1742447, -0.145192, -0.05378577, 
    -0.06898759, 0.04613285, 0.08651371, 0.1702051, 0.2441309, 0.2515691, 
    0.216657, 0.1805404, 0.1757226, 0.1528385, 0.04045236, -0.07523763, 
    -0.2192643, -0.31876, -0.3455341, -0.3326433, -0.3600359, -0.3534928, 
    -0.3443457, -0.3441503, -0.3419695, -0.3001726, -0.2306576, -0.133278, 
    -0.03326178, 0.01636386, 0.03099597, 0.02463222, 0.003619831, -0.1132096, 
    -0.275791, -0.2559831, -0.1695085, 0.1063705, 0.2583399, 0.2015039, 
    -0.0913021, -0.4058529, -0.5149517, -0.457644, -0.3824155, -0.4330177, 
    -0.5873797, -0.7115011, -0.7093689, -0.4663022, -0.3378034, -0.1719174, 
    -0.04066765, 0.04802048, 0.1391667, 0.1582259, 0.1698958, 0.1543522, 
    0.1317448, 0.1202865, 0.07930341, 0.06989568, 0.08975261, 0.172972, 
    0.2695866, 0.338418, 0.3558334, 0.293724, 0.1659245, 0.02805015, 
    -0.04668942, -0.05884764, -0.05484372, -0.008684859, 0.1163151, 
    0.1913965, 0.3004948, 0.4071842, 0.4092675, 0.4934148, 0.4157777, 
    0.1367741, -0.2527118, -0.5099056, -0.6535256, -0.8199158, -0.4716082, 
    -0.3900657, -0.6965756, -0.54363, -0.6446387, -0.7344173, -0.7948503, 
    -0.7630956,
  -0.5191016, -0.3280372, -0.1506934, 0.03732747, 0.2366602, 0.266364, 
    0.418431, 0.4863835, 0.527334, 0.5179915, 0.4490787, 0.3085189, 0.193073, 
    0.110114, 0.09435877, 0.02848953, -0.06954098, -0.2184834, -0.3403584, 
    -0.4172952, -0.4647725, -0.439707, -0.3889096, -0.3675064, -0.3877051, 
    -0.4164811, -0.4309345, -0.3673766, -0.2745706, -0.1826109, -0.1188574, 
    -0.1186296, -0.1491308, -0.1483496, -0.08777014, -0.09834957, 0.01502934, 
    0.1960189, 0.3952538, 0.5935447, 0.6256411, 0.423444, 0.1242253, 
    -0.1969987, -0.4469335, -0.6100684, -0.7905046, -0.9062435, -0.9917741, 
    -0.850791, -0.7322689, -0.510638, -0.2489681, -0.0725522, 0.07638979, 
    0.1696842, 0.2213767, 0.2297914, 0.1150616, 0.1190171, 0.1280013, 
    0.1698958, 0.1154037, 0.09769535, 0.06944013, 0.1048566, 0.129987, 
    0.1274805, 0.1011133, -0.01394202, -0.01262364, -0.09087884, -0.1116146, 
    -0.1122168, -0.1049576, -0.04055333, -0.05414382, 0.003977925, 
    0.03721344, 0.03835249, 0.06540346, 0.1051659, -0.06163096, -0.3879168, 
    -0.5464616, -0.5134864, -0.4398698, -0.2278417, -0.2118912, -0.1706315, 
    -0.3060808, -0.5197201, -0.7903581, -0.9682878, -0.8287858, -0.6982358,
  0.4866765, 0.7849511, 1.048151, 1.247532, 1.368773, 1.397109, 1.287669, 
    0.8990949, 0.4567446, 0.03999674, -0.2131773, -0.3795998, -0.4555762, 
    -0.4415137, -0.3155534, -0.2395605, -0.2997168, -0.3062271, -0.3301692, 
    -0.4179947, -0.4093196, -0.3844987, -0.3524837, -0.3295833, -0.3299902, 
    -0.3341569, -0.2990661, -0.2270445, -0.1039977, 0.06524062, 0.1896875, 
    0.234121, 0.241836, 0.2718815, 0.3420801, 0.3608464, 0.4015365, 
    0.4095769, 0.3957585, 0.279808, 0.07741538, -0.1133236, -0.2626073, 
    -0.3422136, -0.4117448, -0.5108497, -0.6419858, -0.7644954, -0.8182877, 
    -0.7776628, -0.6525, -0.5046489, -0.3636656, -0.2478614, -0.1897724, 
    -0.1569111, -0.142344, -0.1680927, -0.1372334, -0.1155211, -0.1225197, 
    -0.1401956, -0.06498408, -0.1632259, -0.1624773, -0.164349, -0.1634538, 
    -0.1493425, -0.1767187, -0.2847102, -0.3192968, -0.3513769, -0.3653417, 
    -0.2976171, -0.1837174, -0.1054623, -0.05923843, -0.1081315, 0.01605451, 
    0.05222009, 0.03972006, -0.03601265, -0.05023789, -0.05079126, 0.0466373, 
    0.09846032, 0.1013246, 0.161725, 0.1886783, 0.1048567, -0.1296813, 
    -0.2927995, -0.4012305, -0.4351498, -0.2977475, 0.05265953,
  0.5416404, 0.7099673, 0.860065, 0.7783105, 0.4613996, 0.02512026, 
    0.09027338, -0.09644556, -0.2352474, -0.406276, -0.5227474, -0.5653093, 
    -0.5132748, -0.3941342, -0.2683366, -0.181504, -0.1519792, -0.197194, 
    -0.2597754, -0.2913347, -0.3040788, -0.2769141, -0.1822038, -0.1266374, 
    0.0198307, 0.08653, 0.1436589, 0.2083562, 0.2755762, 0.3177963, 0.418431, 
    0.464785, 0.4573469, 0.450625, 0.4232324, 0.3143458, 0.2238672, 
    0.1423243, 0.0345605, -0.07484704, -0.182562, -0.252858, -0.2946875, 
    -0.3054622, -0.3015887, -0.2812762, -0.2902117, -0.3044533, -0.3040951, 
    -0.3056252, -0.3003678, -0.3033466, -0.2955667, -0.2963969, -0.3066508, 
    -0.3275328, -0.3527769, -0.3681902, -0.3754655, -0.3857845, -0.396071, 
    -0.402077, -0.3993261, -0.4260516, -0.4108171, -0.4512467, -0.4380794, 
    -0.4283789, -0.4159928, -0.411989, -0.3962825, -0.3405859, -0.2879167, 
    -0.2157649, -0.2062924, -0.2013118, -0.1882096, -0.1994565, -0.2478938, 
    -0.2346616, -0.2039485, -0.1491961, -0.1031513, -0.07660484, -0.1163183, 
    -0.1294045, -0.119297, -0.1323833, -0.1981058, -0.2410581, -0.2437272, 
    -0.2141213, -0.1171973, 0.01235986, 0.1867416, 0.3633366,
  0.1104719, 0.06310868, 0.008404613, -0.1641052, -0.2149186, -0.2663183, 
    -0.2912045, -0.3046486, -0.2849545, -0.2430274, -0.1841732, -0.1051042, 
    -0.01735997, 0.06174159, 0.09795558, 0.1072004, 0.09790677, 0.07295555, 
    0.05770493, 0.04933894, 0.05550766, 0.08088207, 0.1220767, 0.1889713, 
    0.2718651, 0.2328191, 0.2560612, 0.3535547, 0.3548729, 0.3601627, 
    0.3572005, 0.3065332, 0.2800195, 0.2609277, 0.2421777, 0.2183006, 
    0.1911684, 0.1580305, 0.116071, 0.07303712, 0.04079428, -0.007203728, 
    -0.06753904, -0.1111588, -0.1681738, -0.2059342, -0.2425065, -0.2835709, 
    -0.3191666, -0.3522232, -0.3698828, -0.3762468, -0.3758398, -0.3763606, 
    -0.3736588, -0.3706803, -0.3657324, -0.3525488, -0.3204199, -0.2847265, 
    -0.247552, -0.2362565, -0.2479427, -0.2537207, -0.2481054, -0.2349869, 
    -0.216595, -0.203802, -0.1866471, -0.1804459, -0.1070572, -0.09087896, 
    -0.07818377, -0.1068945, -0.1182227, -0.1541767, -0.174131, -0.1594664, 
    -0.1998798, -0.2240335, -0.1851335, -0.1586686, -0.1079363, -0.08694041, 
    -0.09683609, -0.1369729, -0.1259055, -0.09709692, -0.06880856, 
    -0.02419615, 0.02144194, 0.03739214, 0.03368163, 0.03893864, 0.06891932, 
    0.1047429,
  -0.1002539, -0.07055011, -0.05188155, -0.02046877, 0.008925736, 0.04487938, 
    0.0918358, 0.1247784, 0.1737044, 0.2178288, 0.2579329, 0.2849674, 
    0.2990136, 0.2970605, 0.2913474, 0.2941144, 0.3090557, 0.3225974, 
    0.3241762, 0.3306215, 0.339362, 0.3510644, 0.3559473, 0.368138, 
    0.3857324, 0.4054915, 0.4386458, 0.4670149, 0.447614, 0.4290918, 
    0.4108301, 0.3864974, 0.3575259, 0.3271712, 0.3057683, 0.297793, 
    0.2775782, 0.2573145, 0.2417545, 0.2154851, 0.1744532, 0.1402084, 
    0.1042872, 0.06605473, 0.03677412, 0.00995121, -0.02071285, -0.05490882, 
    -0.0806738, -0.09659176, -0.108636, -0.1208919, -0.1401302, -0.1535091, 
    -0.1588151, -0.162054, -0.1642838, -0.1674902, -0.1685644, -0.1580501, 
    -0.1492447, -0.1414485, -0.1229427, -0.1015397, -0.08620764, -0.06718095, 
    -0.05354162, -0.02566077, 0.004531294, 0.03003585, 0.04183596, 
    0.04525393, 0.05291986, 0.04512373, 0.02821293, 0.03234705, 0.03286787, 
    0.0003646165, 0.0046615, -0.008880138, -0.01903659, 0.007428408, 
    -0.004078746, 0.00122726, -0.02461922, 0.02487624, -0.006504297, 
    -0.04159534, -0.06314456, -0.1114681, -0.1396908, -0.150319, -0.1534279, 
    -0.1521419, -0.142718, -0.1262793,
  -0.0244889, 0.01540369, 0.05666345, 0.110293, 0.1599838, 0.1913475, 
    0.2266504, 0.2605859, 0.2910547, 0.3178449, 0.344375, 0.3630598, 
    0.3801823, 0.394196, 0.4097721, 0.4246484, 0.4435123, 0.4554427, 
    0.4600814, 0.4581283, 0.4612858, 0.4667871, 0.4692448, 0.47722, 
    0.4868717, 0.4871973, 0.4902572, 0.4874903, 0.4820541, 0.4799382, 
    0.4648015, 0.4451075, 0.4317286, 0.4157129, 0.3997135, 0.3790592, 
    0.3569564, 0.3312728, 0.306696, 0.2839258, 0.2518946, 0.2168034, 
    0.1823633, 0.1482812, 0.1179752, 0.08841795, 0.05586588, 0.01582682, 
    -0.02652347, -0.06358403, -0.1042415, -0.1427344, -0.176735, -0.2074805, 
    -0.2399349, -0.267474, -0.2920182, -0.3022884, -0.314349, -0.3302018, 
    -0.3386653, -0.3406673, -0.3350034, -0.3138444, -0.2880794, -0.2643652, 
    -0.2394466, -0.212347, -0.1903092, -0.1626399, -0.1356868, -0.1105729, 
    -0.09387368, -0.08072263, -0.06954098, -0.05821288, -0.05555981, 
    -0.05344394, -0.05642247, -0.06490231, -0.07816732, -0.09286457, 
    -0.1090918, -0.1262304, -0.145485, -0.160345, -0.1722916, -0.1817155, 
    -0.1851334, -0.1818782, -0.1770117, -0.1652278, -0.1447851, -0.1212988, 
    -0.09346676, -0.05886389,
  0.3235765, 0.336791, 0.3453357, 0.3496006, 0.3488519, 0.3447505, 0.3380772, 
    0.3291417, 0.3193111, 0.3095129, 0.3003983, 0.2935134, 0.2892329, 
    0.2873123, 0.2878003, 0.2891352, 0.2914293, 0.2947991, 0.2991769, 
    0.3040926, 0.3105214, 0.3184967, 0.3285069, 0.3411369, 0.356648, 
    0.3753169, 0.3965893, 0.4197018, 0.4431715, 0.4663324, 0.4874916, 
    0.5055413, 0.5211818, 0.5314684, 0.5320544, 0.5293856, 0.5208572, 
    0.5051836, 0.4824132, 0.4543535, 0.4218014, 0.3852942, 0.3454828, 
    0.3027257, 0.257983, 0.2105708, 0.1534255, 0.1042717, 0.06922936, 
    0.0389235, 0.004907131, -0.003605366, -0.06065345, -0.1993415, 
    -0.1571536, -0.2418542, -0.3087649, -0.3321366, -0.2986903, -0.272486, 
    -0.2933683, -0.3768477, -0.337688, -0.3516364, -0.343971, -0.3389416, 
    -0.3380628, -0.3461027, -0.3489022, -0.3329678, -0.3287525, -0.3222585, 
    -0.3053637, -0.2919195, -0.2522719, -0.2721443, -0.2171311, -0.3092375, 
    -0.2213941, -0.2069416, -0.1791902, -0.1491609, -0.1116934, -0.07736731, 
    -0.03773594, 0.001212597, 0.03902197, 0.07577419, 0.1118083, 0.1457934, 
    0.1781831, 0.2095957, 0.2380953, 0.2636156, 0.2864671, 0.3066001,
  -0.06721246, -0.04561406, -0.02276245, -0.008276779, -0.002531335, 
    -0.00803265, -0.02362508, -0.04287964, -0.05953002, -0.06610554, 
    -0.05889517, -0.03858268, -0.008716226, 0.02512157, 0.0556879, 
    0.08299911, 0.1072669, 0.1280189, 0.1427319, 0.1450102, 0.139509, 
    0.1230869, 0.1030831, 0.08319473, 0.07154131, 0.07360888, 0.08719921, 
    0.1124921, 0.1466556, 0.182919, 0.2160087, 0.24192, 0.2587652, 0.2636971, 
    0.2582612, 0.2445726, 0.2250576, 0.2022219, 0.1782465, 0.158438, 
    0.136531, 0.1253658, 0.1275631, 0.1190343, 0.1269119, 0.1628659, 
    0.1198311, 0.1381421, 0.1447992, 0.1193595, 0.1187739, 0.241138, 
    0.06395578, 0.160686, -0.03597951, 0.2277102, 0.183228, 0.1087484, 
    0.0121665, -0.07609797, -0.1562419, -0.2365975, -0.3299248, -0.3996019, 
    -0.4685472, -0.5283126, -0.5525314, -0.5350508, -0.5259849, -0.4690516, 
    -0.3998463, -0.3373303, -0.2956963, -0.2196546, -0.2293866, -0.1846437, 
    -0.1494389, -0.1027104, -0.02873582, 0.003751278, 0.03776765, 0.126049, 
    0.0541091, 0.1761949, 0.123137, 0.1154222, 0.09229374, 0.05873251, 
    0.0227952, -0.0126543, -0.04722452, -0.07559395, -0.09812093, -0.1052828, 
    -0.09746981, -0.08433449,
  -0.6191818, -0.5667566, -0.4816004, -0.3991459, -0.3138595, -0.2266036, 
    -0.1512944, -0.0977298, -0.07466668, -0.081047, -0.1140548, -0.1543705, 
    -0.1794356, -0.1810145, -0.1644783, -0.1551359, -0.1581798, -0.1706948, 
    -0.1902585, -0.2096753, -0.2162204, -0.202548, -0.1631434, -0.1129805, 
    -0.08601117, -0.1001714, -0.1581627, -0.2136155, -0.2463791, -0.2545004, 
    -0.2352464, -0.1842053, -0.1162357, -0.06380987, -0.03184366, 
    -0.007184982, 0.02928734, 0.07914066, 0.1289949, 0.1684799, 0.1889887, 
    0.1964612, 0.1492925, 0.1393628, 0.07134557, 0.06594181, 0.08018357, 
    0.1069739, 0.1372147, 0.1732337, 0.2084224, 0.2459224, 0.281111, 
    0.3056066, 0.3105384, 0.2898679, 0.2577063, 0.2093012, 0.1323156, 
    0.03985143, -0.06744003, -0.1612229, -0.2240159, -0.2551843, -0.2658126, 
    -0.2722089, -0.2849694, -0.2840255, -0.2546473, -0.2110927, -0.1581635, 
    -0.1181734, -0.08687472, -0.06094623, -0.04810429, -0.05038297, 
    -0.05511904, -0.01037669, -0.05977419, -0.06633342, -0.05173379, 
    -0.01605666, -0.02510631, -0.01898658, -0.002384901, 0.02530026, 
    0.005004168, 0.02915788, 0.02372265, -0.06657648, -0.2149329, -0.3599033, 
    -0.5050859, -0.6037526, -0.6479099, -0.6503829,
  -0.7646241, -0.7029061, -0.6860116, -0.6488049, -0.6060798, -0.5584069, 
    -0.4850996, -0.3899823, -0.3002853, -0.2454513, -0.2387293, -0.2746342, 
    -0.3183679, -0.3572676, -0.3935958, -0.4165612, -0.4429123, -0.5189381, 
    -0.6640556, -0.7678623, -0.7332263, -0.6515374, -0.6050372, -0.5843838, 
    -0.5422286, -0.4408615, -0.3670334, -0.3589115, -0.3884201, -0.4314051, 
    -0.4858484, -0.534123, -0.5737065, -0.6074471, -0.6320724, -0.6191652, 
    -0.5733805, -0.5067949, -0.4274321, -0.3231354, -0.2032003, -0.03659725, 
    0.02798653, 0.1241302, 0.1009521, -0.005266428, -0.0621345, -0.03929925, 
    0.01696748, 0.04177204, 0.0757727, 0.08923299, 0.09449008, 0.1128495, 
    0.09658992, 0.05127728, 0.007396221, -0.01342082, -0.01794505, 
    -0.04340029, -0.01787949, -0.08545756, -0.08137226, -0.09587431, 
    -0.07928896, -0.1039641, -0.109709, -0.1244876, -0.1563728, -0.1753349, 
    -0.1827726, -0.1856046, -0.1789474, -0.1790777, -0.1701256, -0.1408615, 
    -0.1000737, -0.02894741, -0.01442912, 0.02569132, 0.08037889, 0.1063717, 
    0.1020748, 0.1272213, 0.1600338, 0.177205, 0.1427321, 0.06763458, 
    -0.06823778, 0.002480984, -0.08910418, -0.2571206, -0.5132403, 
    -0.7378979, -0.8256588, -0.8015866,
  -0.439395, -0.4631581, -0.4934816, -0.3927803, -0.340909, -0.2129464, 
    -0.1914301, -0.2135653, -0.2950268, -0.2022533, -0.1390219, 0.004433632, 
    0.1416273, 0.1857004, 0.1689204, 0.1885984, 0.2121162, 0.2246819, 
    0.2407955, 0.113647, -0.2430415, -0.5496488, -0.8138924, -0.9704013, 
    -1.008113, -0.9050052, -0.7598403, -0.6603277, -0.629648, -0.6475837, 
    -0.673691, -0.6813245, -0.6691329, -0.6339439, -0.5983807, -0.5788496, 
    -0.5655031, -0.5647545, -0.5566492, -0.484286, -0.3256762, -0.1535084, 
    -0.004403353, 0.05467868, 0.02108502, -0.02468324, -0.05832565, 
    -0.02601779, 0.09606874, 0.239998, 0.3606359, 0.4110754, 0.4097571, 
    0.390177, 0.3370521, 0.2589432, 0.209692, 0.2012937, 0.1719316, 
    0.1110103, 0.0413487, -0.0387466, -0.08192635, -0.006600618, 0.05811286, 
    0.107836, 0.1758537, 0.2285066, 0.2393792, 0.1497469, 0.2016187, 
    0.06869245, 0.002058506, -0.001457214, 0.02401495, 0.08296669, 0.2003822, 
    0.2161373, 0.1396073, 0.1445227, 0.1991289, 0.2686439, 0.3133866, 
    0.3841711, 0.4068762, 0.3942134, 0.3600012, 0.3170813, 0.3371335, 
    0.3817948, 0.3523998, 0.09422898, 0.03464413, -0.1656489, -0.3591552, 
    -0.4261627,
  -1.163078, -1.161759, -1.021233, -0.9735427, -0.7975178, -0.5633378, 
    -0.320972, -0.3939221, -0.2990003, -0.2515554, -0.221118, -0.05635548, 
    0.2715421, 0.4479747, 0.373446, 0.1941643, 0.08588004, -0.09353068, 
    -0.1044193, -0.08155143, 0.001016378, -0.02036858, 0.0884366, 0.04906178, 
    -0.01648045, -0.03560448, -0.01351738, -0.01172638, -0.1165771, 
    -0.2619386, -0.4125404, -0.545125, -0.5701904, -0.5834217, -0.6032143, 
    -0.6404543, -0.6453707, -0.6240489, -0.6084888, -0.5150156, -0.4184165, 
    -0.2514091, -0.1722424, -0.09558153, -0.08996642, -0.1650313, -0.1563399, 
    -0.0788497, 0.02298951, 0.1796789, 0.3327388, 0.4477617, 0.4927812, 
    0.5238521, 0.5348059, 0.5003983, 0.4915929, 0.4753495, 0.4705644, 
    0.4263098, 0.3608964, 0.3360754, 0.3921301, 0.4233151, 0.4247636, 
    0.5323971, 0.7870194, 1.09698, 1.379907, 1.557299, 1.61975, 1.372973, 
    1.192211, 1.085555, 0.9303789, 0.8525305, 0.8255611, 0.7825598, 0.692179, 
    0.6979896, 0.4848547, 0.4028559, 0.3741451, 0.4012935, 0.4216874, 
    0.4134191, 0.3611079, 0.3487545, 0.3705644, 0.460164, 0.5295975, 
    0.4527421, 0.3079667, -0.02566028, -0.437607, -0.8791099,
  0.9000565, 0.514298, 0.2079991, -0.003296375, -0.1261647, -0.1270118, 
    -0.05074143, 0.145792, 0.4370844, 0.7545812, 1.0566, 1.438224, 1.751717, 
    1.842635, 1.647566, 1.220173, 0.740454, 0.2256253, -0.08977199, 
    -0.08942938, 0.156339, 0.4933182, 0.743953, 0.7980223, 0.7534742, 
    0.7448153, 0.6900144, 0.7878497, 0.9669025, 1.015698, 1.061092, 
    0.9255295, 0.7042727, 0.604322, 0.3787522, 0.03402424, -0.5813081, 
    -0.5985932, -0.608309, -0.6367593, -0.6370852, -0.5116301, -0.272682, 
    -0.004501581, 0.1675857, 0.3547928, 0.4384354, 0.5046136, 0.5743891, 
    0.634822, 0.7387283, 0.8837638, 1.030053, 1.140209, 1.207299, 1.289493, 
    1.344978, 1.348591, 1.301358, 1.243969, 1.18269, 1.178751, 1.152546, 
    1.053458, 0.9143301, 0.8008211, 0.7768955, 0.8762119, 1.135522, 1.453637, 
    1.746232, 1.950284, 2.053344, 2.043334, 1.929841, 1.817472, 1.803784, 
    1.863631, 1.996866, 2.058846, 1.962394, 1.598087, 1.430769, 1.533357, 
    1.7017, 1.720499, 1.63199, 1.44021, 1.326603, 1.263663, 1.274959, 
    1.297208, 1.352612, 1.40284, 1.294441, 1.155037,
  2.122648, 2.088728, 2.000138, 1.870646, 1.698381, 1.512866, 1.41643, 
    1.401131, 1.391268, 1.333243, 1.327612, 1.505818, 1.855786, 2.281372, 
    2.620419, 2.847729, 2.958667, 2.909823, 2.695044, 2.38959, 2.158016, 
    2.100073, 2.164461, 2.216853, 2.171622, 2.034252, 1.906258, 1.882495, 
    1.859284, 1.76656, 1.627367, 1.531567, 1.581714, 1.746183, 1.844506, 
    1.775643, 1.645125, 1.563598, 1.502742, 1.408504, 1.282331, 1.155395, 
    1.100253, 1.105086, 1.067619, 1.012541, 0.9742265, 1.02032, 1.166495, 
    1.304679, 1.371444, 1.372501, 1.39244, 1.456502, 1.542798, 1.595598, 
    1.621086, 1.605444, 1.558195, 1.513143, 1.487053, 1.45271, 1.389087, 
    1.325741, 1.237134, 1.170744, 1.114282, 1.045842, 0.9581139, 0.9249916, 
    1.027921, 1.2851, 1.604338, 1.85704, 1.969279, 1.93466, 1.862655, 
    1.891268, 2.043661, 2.255656, 2.373072, 2.305656, 2.150464, 2.075041, 
    2.124927, 2.197307, 2.230672, 2.228279, 2.233276, 2.182853, 2.101847, 
    2.034871, 2.013517, 1.995011, 2.026359, 2.086434,
  1.934124, 1.764804, 1.593889, 1.47553, 1.363616, 1.206113, 1.060637, 
    0.9692311, 0.8891206, 0.7701411, 0.6404867, 0.6220121, 0.7075758, 
    0.8349676, 0.9824448, 1.152318, 1.374957, 1.654759, 1.913239, 2.002985, 
    1.926196, 1.831681, 1.802612, 1.833097, 1.870386, 1.865388, 1.845451, 
    1.80621, 1.753411, 1.612232, 1.430592, 1.254126, 1.165243, 1.157415, 
    1.205104, 1.291204, 1.401799, 1.525807, 1.597323, 1.604827, 1.591025, 
    1.60984, 1.647047, 1.700155, 1.794832, 1.865063, 1.894914, 1.918954, 
    1.979419, 2.080233, 2.154288, 2.169915, 2.110914, 2.066545, 2.061728, 
    2.023933, 1.909318, 1.785653, 1.677742, 1.615568, 1.532577, 1.505542, 
    1.539657, 1.523624, 1.448168, 1.413012, 1.421704, 1.363582, 1.180021, 
    1.007137, 0.9457922, 1.041903, 1.240097, 1.428997, 1.546525, 1.603736, 
    1.63803, 1.657089, 1.722861, 1.873382, 2.047519, 2.119524, 2.085735, 
    2.071152, 2.143824, 2.163306, 2.140048, 2.128851, 2.139218, 2.184921, 
    2.258797, 2.352905, 2.418889, 2.381811, 2.240292, 2.084969,
  1.718449, 1.739542, 1.675268, 1.575886, 1.42408, 1.192781, 0.9308176, 
    0.7292862, 0.5892487, 0.4781313, 0.3942289, 0.3312407, 0.2799387, 
    0.3611889, 0.5713615, 0.7707262, 0.8372145, 0.8252363, 0.8472242, 
    0.885685, 0.9236078, 0.9607334, 1.026473, 1.140682, 1.26018, 1.349372, 
    1.390762, 1.389475, 1.392226, 1.430817, 1.460196, 1.40764, 1.296507, 
    1.198119, 1.117781, 1.058568, 1.096638, 1.23399, 1.404172, 1.523102, 
    1.603799, 1.669001, 1.745774, 1.832641, 1.910114, 1.936839, 1.905638, 
    1.844749, 1.809804, 1.83959, 1.932039, 2.061677, 2.101131, 2.002352, 
    1.958894, 1.959009, 1.894588, 1.803589, 1.7545, 1.696167, 1.556453, 
    1.462899, 1.513583, 1.566105, 1.483391, 1.312606, 1.170663, 1.076978, 
    0.9956627, 0.8962002, 0.8397384, 0.8601809, 0.9614348, 1.041577, 
    1.040617, 0.984611, 0.8897715, 0.7641687, 0.6338301, 0.6955657, 
    0.9660892, 1.14174, 1.169735, 1.192798, 1.330004, 1.553101, 1.745092, 
    1.832901, 1.834659, 1.807592, 1.746931, 1.728865, 1.735196, 1.695125, 
    1.619637, 1.641952,
  0.9765854, 0.9469633, 0.8720446, 0.7400951, 0.5871983, 0.4743729, 
    0.4374094, 0.3707104, 0.2595778, 0.1546459, 0.09082603, 0.02878284, 
    -0.0948658, -0.2533464, -0.3373137, -0.2934828, -0.1238537, 0.06447792, 
    0.1352139, 0.1210852, 0.1498451, 0.1814213, 0.1698647, 0.2316322, 
    0.3970785, 0.5725012, 0.7431231, 0.8709068, 0.9375248, 0.9863033, 
    1.039054, 1.044328, 1.035522, 1.030087, 0.9190025, 0.7010174, 0.5209064, 
    0.4586496, 0.5063705, 0.5949287, 0.6240473, 0.5969296, 0.6174698, 
    0.7082253, 0.7782125, 0.7918053, 0.8101635, 0.9339275, 1.109252, 1.21062, 
    1.222207, 1.258064, 1.329028, 1.318448, 1.29353, 1.320271, 1.322144, 
    1.290861, 1.347079, 1.488159, 1.596363, 1.613745, 1.533667, 1.429679, 
    1.343204, 1.228149, 1.095386, 1.024227, 1.022535, 0.9734788, 0.822876, 
    0.6418705, 0.482707, 0.2951908, 0.1333094, 0.07017469, 0.03965664, 
    0.006095886, -0.1007881, -0.1152587, 0.04545164, 0.2532969, 0.432529, 
    0.5072999, 0.6131096, 0.8479891, 1.046002, 1.116462, 1.144912, 1.225234, 
    1.274079, 1.251472, 1.19851, 1.137572, 1.074534, 1.011172,
  0.2803946, 0.2850981, 0.3367434, 0.3384676, 0.2635498, 0.1727457, 
    0.0903244, -0.02989006, -0.1379628, -0.1877027, -0.2906647, -0.4563217, 
    -0.5979724, -0.7347088, -0.8845606, -0.9866619, -0.9721766, -0.8779221, 
    -0.7840738, -0.6578054, -0.4642181, -0.3777599, -0.4871187, -0.5488863, 
    -0.4447193, -0.2455006, 0.01314259, 0.263176, 0.4148197, 0.4998608, 
    0.5783596, 0.606144, 0.6187897, 0.5716047, 0.368659, 0.1358633, 
    -0.02053356, -0.1725674, -0.2947035, -0.2825451, -0.2564058, -0.3755465, 
    -0.5124931, -0.4989185, -0.3441648, -0.1899981, -0.1181393, -0.1053305, 
    -0.0168047, 0.1536865, 0.2358003, 0.2279539, 0.2828207, 0.3959227, 
    0.5071044, 0.639575, 0.7324963, 0.714983, 0.6497812, 0.6467376, 
    0.7600517, 0.8555593, 0.8670015, 0.9249754, 0.9943767, 0.9635172, 
    0.871623, 0.8250732, 0.7752042, 0.6019778, 0.4120364, 0.3064542, 
    0.1480718, -0.06537199, -0.2217035, -0.3298588, -0.3731048, -0.3721774, 
    -0.4633212, -0.6390538, -0.7620358, -0.7624912, -0.6290278, -0.485733, 
    -0.2598867, 0.0267334, 0.2205324, 0.2653732, 0.3236399, 0.4634361, 
    0.5547924, 0.5516834, 0.5173588, 0.4953365, 0.4634027, 0.3764887,
  -0.1411052, -0.05389786, 0.02386999, 0.07974529, 0.1297131, 0.1102467, 
    0.0160408, -0.2070875, -0.465714, -0.5660882, -0.580493, -0.6750078, 
    -0.7831945, -0.8983636, -0.9822507, -1.051001, -1.209008, -1.330085, 
    -1.308292, -1.253083, -1.1878, -1.126326, -1.082804, -0.9938226, 
    -0.7938881, -0.545989, -0.3529377, -0.2379808, -0.184124, -0.1639404, 
    -0.1435947, -0.1984959, -0.3065348, -0.3624759, -0.4043703, -0.4609132, 
    -0.5762935, -0.8282475, -1.028019, -1.071298, -1.151831, -1.314721, 
    -1.400154, -1.292699, -1.075153, -0.943644, -0.8937745, -0.9308019, 
    -0.9201894, -0.7423573, -0.4958568, -0.4562898, -0.535017, -0.5430737, 
    -0.4054432, -0.1896391, -0.008405685, 0.1058359, 0.1005135, -0.01273537, 
    -0.0407629, -0.0377841, 0.02225828, 0.1552005, 0.2671313, 0.3194098, 
    0.3142176, 0.2719979, 0.2497158, 0.136158, -0.008780479, -0.09641075, 
    -0.1841874, -0.18365, -0.2281489, -0.4767346, -0.7069099, -0.8652918, 
    -1.039056, -1.114901, -1.134465, -1.249455, -1.337297, -1.325578, 
    -1.192895, -1.001586, -0.811759, -0.6645741, -0.5195222, -0.426115, 
    -0.3409262, -0.2792888, -0.1790285, -0.07072735, -0.07406425, -0.1468992,
  0.03560448, 0.01674032, 0.02486229, -0.009334564, -0.1108003, -0.2070892, 
    -0.1924405, -0.1688399, -0.3184657, -0.3952724, -0.3331629, -0.2921801, 
    -0.2616625, -0.3083098, -0.4791267, -0.7580006, -1.059204, -1.248837, 
    -1.387965, -1.476295, -1.509839, -1.473902, -1.360489, -1.314851, 
    -1.284855, -1.224047, -1.211564, -1.164379, -1.034496, -0.9837642, 
    -0.9592524, -0.869132, -0.8042722, -0.7434974, -0.7064691, -0.8385334, 
    -1.021948, -1.191187, -1.287313, -1.219866, -1.26202, -1.412411, 
    -1.615569, -1.723332, -1.634302, -1.556747, -1.530787, -1.423658, 
    -1.492311, -1.536011, -1.394557, -1.247959, -1.131764, -1.08357, 
    -1.074944, -0.9608161, -0.8170662, -0.678622, -0.6112881, -0.6972582, 
    -0.7384367, -0.8314054, -0.9247489, -0.9200447, -0.8811779, -0.6499116, 
    -0.5193284, -0.5615487, -0.423317, -0.3146901, -0.2889578, -0.3601, 
    -0.5121837, -0.5907645, -0.7220471, -0.8738046, -0.8503507, -0.8716233, 
    -1.223365, -1.200448, -1.395679, -1.766708, -1.840976, -1.82452, 
    -1.69148, -1.424098, -1.163371, -0.8757076, -0.7556067, -0.7196856, 
    -0.5921464, -0.5579667, -0.475235, -0.2599354, -0.1141672, -0.02258205,
  -0.4691336, -0.5966557, -0.5879482, -0.6917729, -0.7882247, -0.827987, 
    -0.8348231, -0.7160568, -0.6450769, -0.4996179, -0.3258549, -0.3881921, 
    -0.5444746, -0.621916, -0.6481367, -0.7742435, -0.9633224, -1.177173, 
    -1.353345, -1.42815, -1.497958, -1.583944, -1.573983, -1.542229, 
    -1.520223, -1.523869, -1.52618, -1.535686, -1.500073, -1.601082, 
    -1.673902, -1.496461, -1.292522, -1.061858, -0.931454, -1.047909, 
    -1.004354, -0.727808, -0.838306, -1.040829, -1.062427, -1.265373, 
    -1.486109, -1.794849, -1.941985, -1.922209, -2.006568, -2.062671, 
    -2.033147, -1.977466, -1.801685, -1.693091, -1.605347, -1.52758, 
    -1.471672, -1.38357, -1.255038, -1.082919, -0.9999111, -1.082301, 
    -1.168596, -1.303134, -1.417115, -1.370175, -1.412265, -1.307968, 
    -1.280282, -1.426424, -1.335556, -1.310962, -1.251815, -1.165975, 
    -1.166431, -1.119426, -1.082642, -0.7747318, -0.2882409, -0.4267665, 
    -0.7950444, -0.6754807, -0.6778407, -1.270826, -1.56635, -1.719426, 
    -1.622795, -1.217457, -1.132561, -1.060035, -0.9448981, -0.9208906, 
    -0.8184495, -0.7503672, -0.624244, -0.4302661, -0.3712168, -0.3546157,
  -0.6912682, -0.7221113, -0.7033612, -0.7036383, -0.4475996, -0.2029708, 
    -0.2541265, -0.3107019, -0.3927006, -0.4677981, -0.3247321, -0.3194587, 
    -0.3790455, -0.4027596, -0.3880301, -0.5454676, -0.872112, -1.190129, 
    -1.312574, -1.294052, -1.362086, -1.470484, -1.533391, -1.588111, 
    -1.586272, -1.534873, -1.469052, -1.429924, -1.313957, -1.169345, 
    -0.9711676, -0.7392174, -0.645923, -0.5725835, -0.5148199, -0.573495, 
    -0.6404058, -0.5083582, -0.542782, -0.7858648, -0.9263759, -1.270858, 
    -1.489608, -1.630136, -1.805966, -1.881568, -2.038046, -2.156243, 
    -2.123805, -2.044964, -1.90525, -1.761858, -1.598674, -1.27649, 
    -1.041887, -1.055803, -1.125969, -1.177434, -1.168791, -1.169377, 
    -1.138013, -1.109123, -1.150676, -1.168043, -1.314315, -1.388013, 
    -1.490373, -1.6705, -1.688062, -1.795647, -1.809107, -1.752157, 
    -1.601555, -1.272079, -1.038192, -0.6088953, -0.009123266, 0.1079504, 
    -0.5186936, -0.5039471, -0.2889898, -0.654175, -0.8894289, -1.19939, 
    -1.463583, -1.218628, -1.089332, -1.076425, -0.9573653, -0.8698001, 
    -0.9005294, -0.929224, -0.8479903, -0.708342, -0.6707605, -0.6661218,
  -0.8255954, -0.6897225, -0.6052167, -0.3497002, 0.1217523, 0.2317133, 
    0.1921139, -0.006307382, -0.3341721, -0.4401457, -0.5401621, -0.7413812, 
    -0.7315345, -0.6325765, -0.4682045, -0.4188061, -0.4585037, -0.4605222, 
    -0.5772538, -0.6779046, -0.7195063, -0.7882409, -0.8493247, -0.9056396, 
    -0.8337812, -0.7216058, -0.678751, -0.7252192, -0.5986896, -0.4049067, 
    -0.2526789, -0.2647712, -0.332057, -0.3780849, -0.3794196, -0.1424892, 
    -0.03109586, -0.07341361, -0.2349217, -0.5314867, -0.811012, -1.101228, 
    -1.291788, -1.440975, -1.624178, -1.650529, -1.627645, -1.534595, 
    -1.329077, -1.242733, -1.160929, -0.8950925, -0.6909261, -0.5908124, 
    -0.4922123, -0.5926037, -0.6094656, -0.6545341, -0.7216892, -0.692538, 
    -0.6818609, -0.5832928, -0.5869551, -0.7034264, -0.9229576, -1.033472, 
    -1.095175, -1.299374, -1.464299, -1.675627, -1.687916, -1.594963, 
    -1.398804, -1.14646, -0.7907314, -0.3631269, -0.04530489, 0.4480383, 
    0.07049927, -0.4808193, -0.2667727, -0.3065026, -0.3482343, -0.4573491, 
    -0.9012944, -1.004175, -0.7971442, -0.7312262, -0.7292895, -0.5813403, 
    -0.5369716, -0.5430262, -0.6642989, -0.7381597, -0.7945236, -0.8982027,
  -0.4770427, -0.2792883, -0.05640554, 0.1926343, 0.1821365, 0.0447669, 
    0.13129, -0.1872158, -0.4954355, -0.5151125, -0.7009366, -0.7935953, 
    -0.7268469, -0.5010333, -0.3025632, -0.2257566, -0.1620684, -0.005899906, 
    -0.1260486, -0.308959, -0.3769274, -0.5296946, -0.5826244, -0.5338449, 
    -0.5184808, -0.4318104, -0.3127351, -0.2614985, -0.06032705, 0.1437588, 
    0.2681072, 0.157022, 0.05498791, 0.1352139, 0.08335781, 0.01870966, 
    0.0784905, 0.1570392, 0.1354566, -0.07697892, -0.5073652, -0.5704837, 
    -0.507966, -0.6081123, -0.7008209, -0.6788483, -0.5996003, -0.5164461, 
    -0.47683, -0.3963776, -0.3453851, -0.1445713, 0.02875233, -0.1270261, 
    -0.2262611, -0.4304442, -0.4666419, -0.4954512, -0.6077731, -0.4836195, 
    -0.4229424, -0.3336844, -0.4201915, -0.6175063, -0.8201916, -1.062477, 
    -1.260947, -1.45512, -1.434661, -1.510864, -1.511646, -1.46316, 
    -1.333862, -1.081861, -0.5618746, -0.02688038, -0.05874884, 0.2223384, 
    0.006339103, -0.3694911, -0.1646897, -0.1603606, -0.3346605, -0.1744227, 
    -0.3000414, -0.483619, -0.6113689, -0.6100836, -0.7474203, -0.7090259, 
    -0.7098875, -0.6496825, -0.6984296, -0.73842, -0.684123, -0.6398683,
  -0.1720943, -0.008796692, 0.2509997, 0.3850825, 0.06156373, -0.1068125, 
    0.02966213, -0.2938566, -0.2941012, -0.2982508, -0.4336184, -0.3228601, 
    -0.217245, -0.0786221, 0.0448637, 0.07253504, -0.06467295, -0.1546292, 
    -0.1949615, -0.3424392, -0.2779365, -0.1999745, -0.2606678, -0.2913647, 
    -0.2696037, -0.1265044, 0.02427673, 0.007853508, 0.2208095, 0.4909916, 
    0.6501713, 0.8621836, 0.5882902, 0.2810473, 0.3243899, 0.4418221, 
    0.4032462, 0.5103264, 0.1907294, 0.198267, 0.2371674, 0.4050374, 
    0.5420504, 0.3415456, 0.211256, 0.2176032, 0.4698329, 0.6219163, 
    0.5564704, 0.5773034, 0.5708256, 0.3805914, 0.283277, 0.1554451, 
    0.02189875, -0.2551522, -0.3387132, -0.3893807, -0.5427177, -0.6607027, 
    -0.8324802, -0.8269465, -0.8276777, -0.9085696, -0.9857337, -1.129419, 
    -1.209724, -1.264722, -1.181193, -1.217113, -1.204434, -1.156469, 
    -0.9667397, -0.603101, -0.3228273, 0.05609488, 0.3437903, 0.5518306, 
    -0.08003786, -0.2156825, -0.01975143, -0.1468513, -0.2628994, -0.2774997, 
    -0.218857, -0.2724535, -0.2789955, -0.3030024, -0.4719315, -0.5776281, 
    -0.6690831, -0.7306881, -0.7460036, -0.6596918, -0.5363522, -0.3434811,
  0.07530165, 0.2201729, 0.395483, 0.7697343, 0.5190992, -0.137363, 
    0.05449986, -0.08689094, -0.1399183, -0.04955268, 0.06693481, 0.2608475, 
    0.07630992, 0.08824015, 0.04465199, 0.01252508, -0.1929274, -0.3190184, 
    -0.1710038, -0.1988521, -0.1770096, 0.09664011, 0.03713512, -0.08283615, 
    -0.02964592, 0.1290455, 0.3407965, 0.3440681, 0.6064053, 1.02491, 
    1.21464, 1.439119, 1.515079, 0.7333407, 0.7370198, 0.6912682, 0.5869708, 
    1.173625, 0.6730714, 0.9142179, 1.041757, 1.162264, 1.381877, 1.318579, 
    1.219621, 0.7282143, 0.5189197, 0.7246485, 0.8826406, 0.6728587, 
    0.5003817, 0.1831124, -0.1968842, -0.2701104, -0.2564049, -0.4744883, 
    -0.5332932, -0.623023, -0.7271409, -0.8641195, -0.9497967, -0.9383869, 
    -0.9238524, -1.006193, -1.015339, -0.9392648, -0.8492584, -0.7710686, 
    -0.769896, -0.7791247, -0.7196846, -0.627677, -0.4878821, -0.272078, 
    -0.1243579, 0.1190506, 0.3663814, 0.4314529, -0.06400621, -0.1121505, 
    -0.0452885, -0.2466402, -0.1748947, -0.2038012, -0.3580329, -0.3537204, 
    -0.2668858, -0.4168534, -0.5707912, -0.6081128, -0.61975, -0.5877352, 
    -0.4624748, -0.2811599, -0.1815996, -0.06545353,
  0.02064538, 0.05573678, 0.1420487, 0.7207435, 0.8483639, 0.2703035, 
    0.28977, 0.2762928, 0.02414489, 0.08674264, -0.08404177, 0.1113197, 
    0.2179277, 0.1068764, 0.2103755, 0.2737048, 0.1803784, 0.1136305, 
    0.3047106, 0.3743565, 0.2199287, 0.4434311, 0.5456138, 0.5787354, 
    0.4700279, 0.5855372, 0.8336332, 0.6956611, 0.5147202, 0.6254468, 
    0.9080472, 0.901423, 1.226408, 1.421216, 1.572045, 0.9355707, 0.8039141, 
    1.480982, 0.8589425, 1.485734, 1.710506, 1.377319, 1.300171, 1.365015, 
    1.628198, 1.286482, 0.6513586, 0.3422279, 0.2723873, -0.3171151, 
    -0.6918547, -0.7242932, -1.015732, -1.029452, -0.7489498, -0.7332273, 
    -0.5752358, -0.5170326, -0.4624915, -0.5137935, -0.4867916, -0.44628, 
    -0.4524975, -0.4867425, -0.4503489, -0.4142489, -0.4528227, -0.4095283, 
    -0.380671, -0.2799873, -0.2758379, -0.2517653, -0.152986, -0.1387949, 
    -0.07707572, 0.1158118, 0.1880774, 0.04811966, -0.03928256, -0.01691937, 
    0.03008585, -0.1081953, -0.1867437, -0.2129645, -0.339479, -0.4051852, 
    -0.18855, -0.2163973, -0.1766353, -0.1337314, -0.2456131, -0.1940832, 
    -0.1496329, -0.1232333, 0.008993149, 0.02372217,
  0.1419506, 0.1631262, 0.1470292, 0.2804604, 0.5932369, 0.5557693, 
    0.4286209, 0.5386469, 0.3787348, 0.3501867, 0.004922986, 0.03550565, 
    0.1556717, -0.1118579, 0.1495519, 0.2894607, 0.3227454, 0.2139238, 
    0.2024492, 0.230037, -0.005037904, 0.03179479, 0.09743631, 0.2845777, 
    0.2595291, 0.402563, 0.3956457, 0.07451952, -0.1662196, -0.211288, 
    0.1460199, 0.2702875, 0.3995359, 0.6511635, 1.044018, 1.019311, 1.225692, 
    1.370922, 0.2765214, 0.3377681, 0.8952223, 0.7740308, 0.5410721, 
    0.4812252, 0.5767004, 0.5630774, 0.1848059, -0.3029871, -0.3665937, 
    -0.5068605, -0.7111253, -0.8112881, -0.9618907, -1.113877, -0.8879476, 
    -0.8700929, -0.6660404, -0.520792, -0.3569574, -0.3328362, -0.2524323, 
    -0.2227612, -0.2361236, -0.1980863, -0.1373768, -0.1100821, -0.06576252, 
    -0.09004736, -0.1347079, -0.1632729, -0.1702709, -0.1832113, -0.1406016, 
    -0.06062078, -0.05184782, 0.1133868, 0.03011823, -0.1040449, -0.05324748, 
    -0.02380413, -0.1011479, -0.1197026, -0.1380619, -0.2303144, -0.4812596, 
    -0.3939874, -0.2479906, -0.2624111, -0.2619889, 0.07369041, 0.2300372, 
    0.1696863, 0.1567307, 0.1851149, 0.1727281, 0.1334054,
  0.07228962, 0.005264878, 0.1513096, 0.1746824, 0.5623121, 0.371069, 
    0.2772538, 0.6188879, 0.6850013, 0.4941969, 0.3297927, 0.2357824, 
    0.3031979, 0.01781386, 0.1754309, 0.257511, 0.2371496, 0.03596115, 
    -0.2070889, -0.3680587, -0.4978113, -0.3657964, -0.3070236, -0.07093942, 
    -0.1554122, -0.1693934, -0.2275963, -0.2964604, -0.2541264, -0.3189212, 
    -0.369312, -0.4205328, -0.2617437, -0.06760287, 0.1058182, 0.252205, 
    0.1294674, 0.01429814, -0.02689657, 0.09237427, 0.06483519, -0.2472579, 
    -0.4649337, -0.4239506, -0.5683028, -0.4938561, -0.5919846, -0.8395429, 
    -0.8267499, -0.6913823, -0.5437752, -0.4587166, -0.3148854, -0.3851976, 
    -0.2995374, -0.3753674, -0.2922289, -0.2198493, -0.1642666, -0.1319425, 
    -0.005053997, 0.0681715, 0.03064013, -0.01887226, 0.03072119, 
    -0.002514362, -0.01825285, -0.05363703, -0.0482831, -0.1692474, 
    -0.1053152, -0.08217049, -0.07064641, 0.05951285, 0.1608313, 0.2522213, 
    -0.121037, -0.03226766, -0.03140503, -0.03145373, -0.04816926, 
    -0.1107181, -0.1110273, -0.06678915, -0.2261151, -0.2149823, -0.1240971, 
    -0.1582451, -0.1093998, 0.1386795, 0.3269281, 0.2947996, 0.2850337, 
    0.2822016, 0.1582272, 0.1444412,
  0.006274223, -0.055884, 0.06416774, 0.2891679, 0.1119217, -0.009106755, 
    -0.007365331, 0.05601358, 0.3120032, 0.7778233, 0.7843173, 0.3722082, 
    0.6056392, 0.4080482, 0.3567459, 0.3398189, 0.08941221, -0.0005946159, 
    -0.2794032, -0.6195726, -0.7640386, -0.8238531, -0.7718188, -0.5645273, 
    -0.4982506, -0.3323328, -0.4281663, -0.172209, -0.1692631, 0.03155071, 
    -0.02845907, -0.1684981, -0.09924358, -0.08682513, -0.1081791, 
    -0.05397987, -0.04538614, -0.1363855, -0.1334884, 0.1675533, -0.2761154, 
    -0.646672, -0.9692304, -1.055591, -1.151327, -0.9321053, -0.7831149, 
    -0.7463794, -0.6460378, -0.5880461, -0.3223062, -0.2112713, -0.1403885, 
    -0.07038498, 0.1275477, 0.1834073, 0.3648195, 0.4863033, 0.5305419, 
    0.5608146, 0.6415107, 0.6881254, 0.7344637, 0.5726149, 0.4913814, 
    0.3810624, 0.3036535, 0.2659258, 0.1980382, -0.004305363, -0.1233972, 
    -0.1993575, -0.1606205, -0.2019943, -0.01420128, 0.2648514, -0.01481998, 
    -0.01574748, -0.01874226, 0.01151487, 0.0419836, -0.1592373, -0.1045499, 
    -0.01952362, -0.02987492, 0.07085729, 0.1887609, 0.2512935, 0.2607174, 
    0.1452551, 0.2506751, 0.322599, 0.2194902, 0.2300533, 0.2144119, 0.1809486,
  -0.1496997, -0.100693, -0.1302667, 0.1329178, 0.04852659, 0.01792765, 
    0.03238077, 0.01135212, 0.2010331, 0.7641842, 1.163452, 0.3470616, 
    0.3329992, 0.3894286, 0.4038001, 0.4415442, 0.1916418, 0.04921007, 
    -0.4310632, -0.8109949, -0.9510665, -1.130949, -1.097844, -0.9980071, 
    -0.7684171, -0.304924, -0.3576585, -0.2111902, -0.4027105, -0.1702071, 
    -0.2564376, -0.05339397, -0.09898317, -0.4136477, -0.4344159, -0.4195397, 
    -0.3187752, -0.3507903, -0.3607345, -0.3072681, -0.5206635, -0.4487557, 
    -0.4024663, -0.33676, -0.2183504, -0.02276182, 0.0312748, 0.08134031, 
    0.1658778, 0.07305527, 0.1385179, 0.1569586, 0.1110601, 0.006323814, 
    -0.01410246, -0.04961681, -0.01600695, 0.04978085, 0.1441493, 0.2633224, 
    0.3266683, 0.3196037, 0.4549711, 0.543009, 0.6710041, 0.6619705, 
    0.5647537, 0.4517493, 0.2978918, 0.1308182, 0.05518365, 0.03936315, 
    -0.08142114, -0.5349371, -0.3354254, 0.08399212, -0.007381618, 
    0.01766729, 0.1160559, 0.07482868, 0.02040172, 0.005102098, -0.1779873, 
    0.1804934, 0.3275805, 0.4711821, 0.6435459, 0.6257237, 0.5816972, 
    0.3305742, 0.3021725, 0.1497796, -0.05710506, 0.003310919, 0.08973718, 
    0.03511477,
  -0.0673424, -0.07743382, 0.03631949, 0.1717361, 0.2690017, 0.1258866, 
    0.228035, 0.414591, 0.2562251, 0.2530513, 0.7645912, 0.4453691, 
    0.2524979, 0.5899646, 0.5288486, 0.4524165, 0.2736893, -0.006730556, 
    -0.2901454, -0.626864, -1.075724, -1.308944, -1.451978, -1.29939, 
    -1.062102, -0.5744877, -0.1185308, -0.3908289, -1.340358, -1.456616, 
    -1.222291, -0.3565841, -0.1322515, -0.6061288, -0.6107011, -0.2901621, 
    -0.3170824, -0.284384, -0.22963, -0.1711502, -0.1699619, -0.1459875, 
    -0.04645967, 0.0288825, 0.1716566, 0.2455335, 0.2509041, 0.3197355, 
    0.3720469, 0.4196057, 0.4104419, 0.3904715, 0.3936939, 0.2218676, 
    0.04045534, -0.1292877, -0.3387928, -0.4362864, -0.38837, -0.3496499, 
    -0.3257885, -0.1958899, -0.04453945, 0.07969451, 0.2034905, 0.1848547, 
    0.1635331, 0.06032676, -0.05751181, -0.1926518, -0.2959233, -0.2194914, 
    -0.1747808, -0.3037033, -0.174732, 0.05632284, 0.191658, 0.1834549, 
    0.2010005, -0.08640182, 0.02549529, -0.02813387, -0.06808996, 0.2556243, 
    0.4601321, 0.5770268, 0.6710532, 0.6224678, 0.6172928, 0.5192298, 
    0.4112219, 0.106925, -0.1058364, -0.1959887, -0.01397359, 0.02948362,
  0.00720185, -0.002189636, 0.09837997, 0.150203, 0.131632, 0.03815877, 
    0.09717569, 0.06296343, 0.07084106, 0.2171627, 0.4244543, 0.2002517, 
    -0.0922935, 0.1568596, 0.2383375, 0.3850011, 0.3600336, 0.160522, 
    0.07422638, -0.3746018, -0.5529046, -0.362834, -0.7304777, -1.04161, 
    -1.176571, -1.261451, -1.452889, -1.635669, -2.038518, -2.052743, 
    -1.836158, -1.029257, -0.3585371, -0.334823, -0.5954666, -0.3076425, 
    -0.1675048, -0.2210689, -0.2205482, -0.2492423, -0.2009673, -0.1805573, 
    -0.126586, -0.01984787, 0.05506897, 0.02154064, 0.03055859, 0.1092205, 
    0.1134186, 0.1320066, 0.2130127, 0.2487707, 0.2081137, 0.1106682, 
    -0.04135036, -0.2441168, -0.4582119, -0.5534263, -0.4910722, -0.3658276, 
    -0.3313551, -0.2301502, -0.09491301, 0.0419035, 0.02661991, -0.08905578, 
    -0.08739495, -0.1614344, -0.1334232, -0.1315191, -0.1306238, -0.1527102, 
    -0.2901618, -0.08562088, 0.01200315, 0.09707804, 0.09112072, 0.03296685, 
    0.09808826, -0.1054435, -0.0468998, -0.1098871, -0.01231194, 0.4190035, 
    0.5337658, 0.650806, 0.7624435, 0.7378664, 0.7793362, 0.8154047, 
    0.7284745, 0.5159414, 0.4159918, 0.3059807, 0.1043046, 0.06966901,
  0.1188228, -0.08742717, -0.2741785, -0.3050053, -0.4581627, -0.5681888, 
    -0.4101331, -0.4444587, 0.05951297, 0.444474, 0.2197018, -0.02585495, 
    -0.2855231, -0.1665297, 0.06885457, 0.2821043, 0.3010168, 0.2130448, 
    0.218546, -0.03029823, 0.1211333, -0.03054231, -0.5410569, -1.096086, 
    -1.275936, -1.210784, -1.506503, -1.10258, -0.5975345, -0.7498945, 
    -0.9315031, -0.9552982, -0.7615814, -0.4699309, -0.41962, -0.3912511, 
    -0.3758535, -0.4685946, -0.3818269, -0.3587799, -0.3729076, -0.2833896, 
    -0.1513758, -0.0649662, 0.02855587, 0.02670097, 0.03963947, 0.06973267, 
    0.10567, 0.09237289, 0.1201239, 0.1379776, 0.07069302, -0.1003847, 
    -0.3329353, -0.4472904, -0.5475836, -0.5559654, -0.5041103, -0.3818598, 
    -0.2990966, -0.1986074, -0.04813576, 0.03431845, 0.02958202, -0.0164156, 
    -0.06983304, 0.02603322, 0.346606, 0.3958899, 0.675024, 0.9139401, 
    0.1300373, -0.1465731, -0.09434271, -0.263648, -0.1719971, -0.1525307, 
    -0.06267166, -0.05601597, 0.04945469, 0.1048918, 0.3104095, 0.4344816, 
    0.4702563, 0.5808196, 0.6540289, 0.7328377, 0.8451095, 0.9344153, 
    0.9908936, 0.9444414, 1.115567, 0.7093012, 0.40214, 0.2778398,
  -0.3635988, -0.3800541, -0.3846447, -0.4040942, -0.5258396, -0.6487226, 
    -0.297014, 0.01099324, 0.3255774, 0.3318273, 0.444181, 0.2178788, 
    -0.3618736, -0.1194913, 0.1577713, 0.1442297, 0.2211829, 0.2357174, 
    0.310945, 0.376163, 0.3256583, -0.4318446, -0.7051681, -0.744117, 
    -0.6470299, -0.4830165, -0.522258, -0.9704839, -0.8349695, -0.5763929, 
    -0.4817152, -0.3936286, -0.5127697, -0.5201092, -0.6351151, -0.6330314, 
    -0.6815348, -0.6801348, -0.6444082, -0.6466055, -0.5687084, -0.4664297, 
    -0.3925209, -0.4104571, -0.2988853, -0.2431078, -0.1665134, -0.08428574, 
    -0.006112099, 0.1051846, 0.1639738, 0.1313057, -0.01014996, -0.2636967, 
    -0.5110598, -0.6062756, -0.7787037, -0.7918053, -0.7385345, -0.6449137, 
    -0.5246501, -0.4182367, -0.2849522, -0.217309, -0.06423378, 0.06201911, 
    0.1524488, 0.3605383, 0.4790606, 0.2300859, 0.1246986, 0.3743404, 
    -0.4377367, -0.4724364, -0.2378001, -0.2298431, -0.1524668, -0.2839289, 
    -0.3186131, -0.1660714, -0.0299387, 0.02956629, 0.2125578, 0.2983165, 
    0.4790783, 0.5476818, 0.6158128, 0.6897554, 0.786809, 0.8938398, 
    0.8676677, 0.8298417, 0.4334223, 0.03457785, -0.1915133, -0.2966235,
  -0.52522, -0.6491133, -0.7038332, -0.5456953, -0.5205331, -0.5466884, 
    -0.3814542, -0.1547451, 0.107283, 0.1541419, 0.6103266, 0.0840735, 
    -0.8667738, -0.3122642, -0.03487184, -0.3230554, -0.1865645, 0.06559992, 
    -0.06623673, -0.2307549, -0.08306623, -0.3577398, -0.704452, -0.5770922, 
    -0.4628832, -0.2798426, -0.1176518, -0.5582117, -0.5287195, -0.2368419, 
    -0.2235608, -0.8015718, -1.151425, -1.012884, -1.060572, -1.014722, 
    -1.084725, -1.084497, -1.05087, -0.9778562, -0.766902, -0.754272, 
    -0.7434964, -0.7288971, -0.6135979, -0.6564693, -0.6339436, -0.4997306, 
    -0.3663154, -0.217927, -0.1512613, -0.1601806, -0.3349195, -0.5591707, 
    -0.8409252, -1.073918, -1.122257, -1.02779, -0.9692783, -0.8615303, 
    -0.7739816, -0.7062907, -0.5206947, -0.3344164, -0.1229093, 0.0486728, 
    0.4183673, 0.5992755, 0.5607661, 0.1392981, 0.03420353, -0.2500736, 
    -0.8128183, -0.7211666, -0.547648, -0.4631095, -0.5040927, -0.5527253, 
    -0.3173742, -0.2070713, -0.1186438, 0.04790926, 0.2038989, 0.233326, 
    0.2841558, 0.2744226, 0.4024501, 0.4382572, 0.4908619, 0.6172123, 
    0.5407147, 0.478523, -0.01120663, -0.4069593, -0.6118908, -0.5965903,
  -0.5591881, -0.6764571, -0.8218347, -0.5343183, -0.5719973, -0.424162, 
    -0.14537, -0.276083, -0.08348837, -0.001994252, -0.3150965, -0.9808354, 
    -0.9628016, 0.01057088, 0.1204994, -0.5327722, -0.636923, -0.204973, 
    -0.09537077, -0.2492278, -0.1922615, -0.2713629, -0.4320723, -0.1212327, 
    -0.09473515, -0.1472579, 0.02137828, -0.6784258, -0.4082768, -0.01123917, 
    -0.1980389, -0.4885176, -0.444247, -0.5296962, -0.6756921, -0.6638107, 
    -0.866138, -1.032805, -1.0344, -1.037216, -0.9940689, -1.046803, 
    -1.059986, -1.199553, -1.271493, -1.192716, -1.062605, -1.016544, 
    -0.8653398, -0.7059975, -0.748836, -0.8205643, -1.020288, -1.217179, 
    -1.405558, -1.557316, -1.552677, -1.453605, -1.308259, -1.148592, 
    -1.046769, -0.8174233, -0.5726981, -0.4214282, -0.1243575, 0.1551347, 
    0.3605049, 0.5728432, 0.3695064, 0.09421346, -0.2598882, -0.6337173, 
    -0.7917719, -0.5896401, -0.6852131, -0.7521892, -0.7405841, -0.6503658, 
    -0.4933844, -0.4878349, -0.3089445, -0.1954515, -0.1179776, -0.01260662, 
    0.07985783, 0.1072178, 0.0677495, 0.009644032, 0.01617098, 0.04859257, 
    0.04711151, 0.1361895, -0.186076, -0.6173424, -1.018319, -0.9207277,
  -0.6883226, -0.7476486, -0.7248948, -0.4273198, -0.3659753, -0.1330003, 
    0.001114488, -0.3687586, -0.247144, -0.1280846, -0.8256921, -1.121265, 
    -0.3324467, 0.2859615, -0.1748948, -0.6489832, -0.2666752, 0.1486727, 
    -0.09055257, -0.3343673, -0.1836674, -0.291838, -0.114185, 0.4381578, 
    0.01055467, -0.1332278, -0.2368577, -0.8568776, -0.1454678, 0.3023676, 
    0.1465733, 0.2464271, 0.191528, 0.1529862, -0.002873063, -0.1737553, 
    -0.4134037, -0.5322025, -0.5978112, -0.7928308, -0.9954839, -1.19467, 
    -1.271737, -1.424114, -1.558439, -1.511158, -1.432593, -1.441464, 
    -1.372242, -1.366888, -1.406601, -1.374212, -1.490959, -1.663958, 
    -1.812867, -1.908326, -1.895045, -1.693417, -1.333163, -1.033993, 
    -0.8002365, -0.5595785, -0.3798752, -0.1885665, 0.1401112, 0.1452382, 
    0.04709387, 0.130167, 0.2382889, -0.1278244, -0.52719, -0.7027106, 
    -0.5495203, -0.2966232, -0.4242926, -0.5734951, -0.7404221, -0.6205979, 
    -0.5320723, -0.4960209, -0.374325, -0.4576095, -0.4007736, -0.3398035, 
    -0.3386639, -0.3224045, -0.4386809, -0.4766529, -0.5436287, -0.664511, 
    -0.6913173, -0.6317797, -0.4828371, -0.5061121, -0.6315026, -0.6828048,
  -0.4416752, -0.3704186, -0.4378341, -0.5159753, -0.4848556, -0.3225672, 
    -0.3074141, -0.434058, -0.4579024, -0.4217694, -0.5611253, -0.269556, 
    0.3418696, 0.06476998, -0.6693443, -0.6828212, -0.1684819, 0.03050923, 
    -0.07238817, 0.1610265, 0.2782304, 0.1601632, 0.2246161, 0.1394453, 
    -0.2958899, -0.1108475, -0.3760648, -0.5496017, -0.002727032, 0.3037999, 
    0.2201736, 0.3434975, 0.3414302, 0.4854568, 0.4356197, 0.2388913, 
    0.07572389, -0.1167405, -0.3988694, -0.7168705, -0.9923588, -1.279127, 
    -1.492684, -1.592912, -1.569133, -1.557642, -1.613192, -1.603817, 
    -1.589559, -1.626734, -1.566008, -1.597502, -1.735393, -1.762671, 
    -1.834644, -1.877499, -1.682382, -1.328329, -0.9758386, -0.6255131, 
    -0.2061771, 0.01983196, 0.1525469, 0.344913, 0.3142662, 0.3248932, 
    0.4268309, 0.5706297, 0.4945226, 0.1282466, -0.06537318, -0.1164149, 
    -0.1233647, -0.1184493, -0.101506, -0.1264733, -0.2193121, -0.218596, 
    -0.1410739, -0.1033778, -0.1648202, -0.3089607, -0.2864189, -0.3800383, 
    -0.5384688, -0.6770267, -0.8496669, -0.8885338, -1.028768, -1.182675, 
    -1.244865, -1.29703, -1.179192, -0.9454514, -0.5797285, -0.4752527,
  -0.6766686, -0.6766362, -0.7000901, -0.5886968, -0.2981369, -0.2035406, 
    -0.1402756, -0.2466561, -0.415992, -0.2495537, 0.01188922, 0.08986795, 
    0.009708166, -0.3577886, -0.4607995, -0.2869226, -0.3400964, -0.2268965, 
    0.3330644, 0.5798092, 0.4288318, 0.05716896, -0.2078376, -0.2765865, 
    -0.09807062, -0.1149833, -0.08819294, 0.1278723, 0.3661046, 0.05542764, 
    -0.2559819, -0.08182815, 0.03016734, 0.06543738, -0.1147709, -0.3093024, 
    -0.3274826, -0.3617271, -0.5546966, -0.7549076, -1.066056, -1.267392, 
    -1.331584, -1.394621, -1.353834, -1.200301, -1.187264, -1.311499, 
    -1.452157, -1.492309, -1.482495, -1.62522, -1.756877, -1.730965, 
    -1.677613, -1.448821, -1.065894, -0.687216, -0.2796314, 0.1112704, 
    0.4563549, 0.6994531, 0.6848214, 0.4478097, 0.2772532, 0.5438881, 
    0.7031489, 0.6601152, 0.4547931, 0.2674718, 0.2399817, 0.1640377, 
    0.1143632, 0.01535594, -0.1029221, -0.07220912, 0.06841612, 0.04305792, 
    -0.02762938, 0.03749132, 0.1566162, 0.2210045, 0.08581543, -0.1791592, 
    -0.3883715, -0.5913007, -0.7060633, -0.7847257, -1.044524, -1.200903, 
    -1.30092, -1.421102, -1.396509, -1.306975, -0.9672937, -0.6696701,
  -0.6516039, -0.6508057, -0.2322843, 0.3908114, 0.8047438, 0.7139235, 
    0.447729, 0.2246822, -0.01927924, 0.009952307, 0.05983841, 0.09437621, 
    0.1646234, 0.2505937, 0.2940995, -0.02015829, -0.2304773, -0.08210504, 
    0.2417395, 0.1095617, -0.1608975, -0.3836511, -0.4330815, -0.424748, 
    -0.1315678, 0.03522915, 0.3778397, 0.5884192, 0.5620846, 0.2156003, 
    0.04824984, -0.05057836, -0.1894129, -0.3023362, -0.2992437, -0.282789, 
    -0.231503, -0.1855233, -0.210165, -0.06167746, -0.06550264, -0.2592864, 
    -0.4213781, -0.5381589, -0.6262121, -0.6315832, -0.6660881, -0.6785722, 
    -0.7308021, -0.8656979, -1.09908, -1.337443, -1.364559, -1.267667, 
    -1.079223, -0.6744704, -0.2705646, 0.1151776, 0.6184168, 0.9185958, 
    1.123251, 1.319344, 0.8800037, 0.2178791, 0.2546954, 0.6587316, 0.463647, 
    0.4225335, 0.6920156, 0.8542068, 0.7776606, 0.6604894, 0.5205805, 
    0.3075274, -0.008781433, -0.04540253, 0.04784274, 0.1303618, 0.2509193, 
    0.3431883, 0.3698487, 0.3695717, 0.2618079, -0.007722855, -0.291512, 
    -0.4456463, -0.427124, -0.6147709, -0.9183187, -0.928133, -0.8774498, 
    -0.9044526, -0.842082, -0.6923265, -0.5116458, -0.463599,
  0.1532629, 0.3534091, 0.7891183, 0.9245032, 0.7914628, 0.6069412, 
    0.6274004, 0.5492102, 0.3756424, 0.2907629, 0.2507564, 0.3938065, 
    0.4035885, 0.3454667, 0.2875567, 0.1011633, 0.0854243, 0.239705, 
    0.1836828, -0.06664266, -0.04794149, 0.3114498, 0.4766353, 0.509578, 
    0.3155026, 0.1667232, 0.2579501, 0.3494707, 0.1427813, -0.0359627, 
    0.1350987, 0.2676833, 0.2252514, 0.194653, 0.05441833, 0.05246568, 
    0.4684005, 0.7679927, 0.6988513, 0.7410061, 0.7888429, 0.6670332, 
    0.51578, 0.5196047, 0.5314054, 0.4093676, 0.1693935, -0.04138136, 
    -0.2420001, -0.431746, -0.6675858, -0.898982, -0.9207597, -0.6931391, 
    -0.3580966, 0.05411005, 0.3946214, 0.8628016, 1.362509, 1.600252, 
    1.744735, 1.726164, 1.035798, 0.3962318, 0.8478758, 1.061059, 0.6166581, 
    0.6232986, 1.141901, 1.064021, 0.6015538, 0.3593991, 0.1190344, 
    -0.03013563, -0.02037001, 0.1525464, 0.09406662, 0.1132886, 0.2531648, 
    0.2969797, 0.1395249, 0.05834031, 0.1221912, 0.07840848, 0.02355909, 
    0.1155677, 0.1687903, -0.07276154, -0.2667232, -0.2208409, -0.1367102, 
    0.0218997, 0.1515865, 0.04328537, 0.05464554, 0.2211664,
  0.6300048, 0.5779213, 0.7555904, 0.7897376, 0.6469641, 0.7010656, 
    0.7240149, 0.4786698, 0.3063391, 0.3837642, 0.6819901, 0.8219967, 
    0.6461014, 0.2154862, 0.03174615, 0.03101325, 0.1335037, 0.1079665, 
    0.08487082, 0.114705, 0.1820227, 0.1480546, 0.09242309, 0.1006099, 
    0.007234395, 0.001146913, 0.267244, 0.5902745, 0.6431227, 0.6789467, 
    0.8040116, 0.7895577, 0.7301013, 0.6027739, 0.3930733, 0.4284899, 
    0.8282132, 1.385424, 1.382332, 1.152758, 1.20362, 1.333162, 1.504451, 
    1.55787, 1.427303, 1.255216, 1.130737, 0.9141846, 0.6391201, 0.4879155, 
    0.4802499, 0.4600019, 0.5195236, 0.6991787, 0.8727951, 1.092994, 
    1.421623, 1.766398, 2.005689, 1.971118, 1.832495, 1.527823, 0.968888, 
    0.5407954, 0.7548416, 0.9183185, 0.8644117, 1.042943, 1.164655, 0.615128, 
    -0.02950072, -0.3475346, -0.4876062, -0.4134851, -0.1821536, 0.01013136, 
    0.1059483, 0.15712, 0.1720777, 0.09126747, -0.09637928, -0.1788826, 
    -0.06018114, 0.0189364, 0.2439523, 0.6007073, 0.7102458, 0.5092204, 
    0.3779707, 0.377954, 0.4572997, 0.6080647, 0.6427326, 0.5963452, 
    0.7537186, 0.8516839,
  1.213908, 1.310197, 1.533472, 1.262313, 0.8669672, 0.6928298, 0.5104406, 
    0.2384517, 0.1689042, 0.2435462, 0.3318113, 0.3388423, 0.1543861, 
    -0.1329025, -0.3394455, -0.251734, -0.06216663, 0.003458142, 0.1095455, 
    0.3170814, 0.3344641, 0.1640539, 0.07171996, 0.2032466, 0.319783, 
    0.5777587, 0.8657631, 0.763598, 0.502351, 0.5145422, 0.6588619, 
    0.5986073, 0.4047601, 0.3425697, 0.5318103, 0.7290441, 0.7720619, 
    0.7266029, 0.8865963, 1.328767, 1.490583, 1.532495, 1.528279, 1.528426, 
    1.423835, 1.30572, 1.295027, 1.377774, 1.510229, 1.682397, 1.820044, 
    1.940503, 2.104712, 2.197176, 2.169751, 2.22465, 2.433228, 2.555704, 
    2.396427, 1.993464, 1.534692, 1.010636, 0.4157792, 0.1243404, 0.1904538, 
    0.334643, 0.6218829, 0.8006263, 0.5130448, -0.0661543, -0.3452396, 
    -0.2945072, -0.1269617, -0.03928262, -0.08492059, -0.2166914, -0.1869226, 
    -0.1486577, -0.1534265, -0.1985762, -0.2015548, -0.02010942, 0.06021279, 
    -0.01683807, -0.01882398, 0.01387477, -0.01729441, -0.141464, 
    -0.06343675, 0.2666414, 0.6891024, 1.018968, 1.141772, 1.207901, 
    1.338711, 1.303035,
  1.501424, 1.772176, 1.70743, 1.280411, 0.9550533, 0.8505122, 0.6130773, 
    0.2396399, 0.1083736, 0.1251379, 0.1111893, 0.06991333, -0.03430218, 
    -0.1470299, -0.2148686, -0.09359579, 0.1065344, 0.2389074, 0.3682367, 
    0.4987544, 0.5200596, 0.5078037, 0.5403072, 0.5393472, 0.4956785, 
    0.4192461, 0.3531163, 0.3040605, 0.2211341, 0.242586, 0.2921951, 
    0.2815669, 0.2107012, 0.2632076, 0.5888425, 0.8685297, 0.7567785, 
    0.5202226, 0.4395909, 0.6314855, 0.6446204, 0.5000241, 0.466528, 
    0.8179765, 1.224324, 1.560424, 1.838859, 2.173152, 2.515031, 2.676977, 
    2.572192, 2.423413, 2.366576, 2.400707, 2.388028, 2.415518, 2.530492, 
    2.358227, 1.929321, 1.399226, 0.8563554, 0.2814205, -0.1133549, 
    -0.1123621, -0.001196623, 0.1705805, 0.215714, 0.01931095, -0.217489, 
    -0.3203211, -0.2234949, -0.08361857, -0.008439541, 0.00651814, 
    -0.1574793, -0.2279871, -0.2320072, -0.1731693, -0.1922448, -0.2261642, 
    -0.1341069, -0.01470584, 0.1330318, 0.1042883, -0.007039845, -0.1024174, 
    -0.1852789, -0.1054122, 0.1620356, 0.5464431, 0.9334388, 1.260359, 
    1.439314, 1.365405, 1.291251, 1.285766,
  1.533911, 1.555737, 1.140909, 0.6087316, 0.5107175, 0.7590899, 0.6879146, 
    0.2294836, -0.01861207, -0.008244231, 0.06748819, -0.001408294, 
    -0.06203655, -0.08536012, -0.09193563, -0.05150592, 0.01104289, 
    0.0556066, 0.1705317, 0.3031327, 0.3843664, 0.3986895, 0.5756587, 
    0.6363031, 0.5211016, 0.3126382, 0.278442, 0.3042068, 0.2649981, 
    0.2417722, 0.2950594, 0.3796623, 0.4318113, 0.4425535, 0.5341712, 
    0.5992917, 0.4526769, 0.2508378, 0.05277473, -0.3931403, -0.5780199, 
    -0.2427011, 0.2091547, 0.5195714, 1.071883, 1.666903, 1.981519, 2.143872, 
    2.264623, 2.188338, 2.028572, 1.857657, 1.746655, 1.594979, 1.640633, 
    1.717293, 1.715161, 1.322696, 0.6753335, 0.09403396, -0.400627, 
    -0.3197841, -0.2805749, -0.09458858, 0.1795976, 0.2811275, 0.1556718, 
    -0.03817587, -0.09232627, -0.0663498, -0.07286012, -0.2289148, 
    -0.3097416, -0.3744877, -0.450627, -0.4855228, -0.4417565, -0.3379318, 
    -0.240894, -0.1696213, 0.006208837, 0.2242264, 0.4271725, 0.7335199, 
    0.9192297, 0.7774164, 0.578507, 0.5953527, 0.8378332, 1.149015, 1.362963, 
    1.422029, 1.451961, 1.392586, 1.244669, 1.316772,
  0.776163, 0.6056719, 0.2285234, 0.09256957, 0.05537882, 0.1463944, 
    -0.01410361, -0.1007898, -0.06814006, 0.01037557, 0.04792439, 0.01740681, 
    -0.05383342, -0.07121623, -0.07964722, -0.1178634, -0.1622481, 
    -0.1344324, -0.01717979, 0.09128368, 0.1314203, 0.1384515, 0.1179925, 
    0.1164954, 0.1339922, 0.1284419, 0.1478105, 0.154744, 0.09982848, 
    0.08405733, 0.1538652, 0.2790607, 0.3451411, 0.3675371, 0.3661212, 
    0.3164953, 0.2373612, 0.1647376, 0.0776931, 0.1284089, 0.2315991, 
    0.3101797, 0.4305253, 0.6388097, 0.8629959, 0.9455483, 0.825187, 
    0.1791899, -0.07841063, -0.1130791, -0.04538655, -0.02681518, 0.3162837, 
    0.07940221, -0.01177597, 0.02217579, 0.09261858, 0.02650535, -0.07220912, 
    -0.187883, -0.1945398, -0.1328862, -0.03330934, 0.08143675, 0.2355709, 
    0.2737707, 0.1216385, -0.006730497, -0.1061283, -0.2467533, -0.4247969, 
    -0.5283289, -0.5424565, -0.547795, -0.5801029, -0.59231, -0.5878829, 
    -0.3954023, -0.1893803, -0.003117278, 0.1243404, 0.2610103, 0.3081295, 
    0.4603919, 0.4584548, 0.4464757, 0.2525792, 0.247143, 0.4505122, 
    0.6941156, 0.805216, 0.8185132, 0.8072339, 0.7820387, 0.7785883, 0.8071039,
  -0.3442957, -0.5071049, -0.5956953, -0.594198, -0.4506921, -0.3482345, 
    -0.2981693, -0.2201257, -0.1774174, -0.1740645, -0.1868575, -0.2142013, 
    -0.2570886, -0.2934819, -0.3040613, -0.3160567, -0.2760665, -0.1994065, 
    -0.0508222, 0.09727323, 0.2052486, 0.2271724, 0.1389074, 0.03016722, 
    -0.03086787, -0.04473519, -0.03820843, -0.05430549, -0.1110274, 
    -0.1398686, -0.06641471, 0.05936652, 0.1414954, 0.1343339, 0.08503377, 
    0.02119914, -0.03602737, -0.03099805, 0.01830208, 0.03041136, 0.0809322, 
    0.1697506, 0.2341385, 0.3587966, 0.4660232, 0.4980867, 0.4299226, 
    0.3273184, 0.2310457, 0.2343173, 0.2069738, 0.1983966, 0.0345453, 
    -0.01296437, 0.009626985, 0.06161237, 0.1291093, 0.1170487, 0.08472461, 
    0.07713997, 0.1232662, 0.1966224, 0.1942134, 0.1642331, 0.1353757, 
    0.07464969, 0.02028781, -0.07025599, -0.2123133, -0.3519129, -0.4737065, 
    -0.467017, -0.3408289, -0.1973881, -0.07186728, -0.002108157, 0.08596146, 
    0.1843014, 0.2401119, 0.2259029, 0.1714107, 0.2638098, 0.3835039, 
    0.403604, 0.2401111, 0.03242922, 0.06413507, -0.1139896, 0.1500568, 
    0.1310625, -0.1470788, -0.1499276, -0.2158128, -0.1751552, -0.1505783, 
    -0.2060797,
  -1.020549, -1.145679, -1.216968, -1.184612, -1.062688, -0.7419194, 
    -0.5482507, -0.4240971, -0.4000086, -0.4675867, -0.5876551, -0.6623458, 
    -0.6871179, -0.672795, -0.672323, -0.5003015, -0.2776452, -0.05500543, 
    0.1315669, 0.1948806, 0.1469966, 0.09170693, 0.07404745, 0.06529093, 
    0.07491007, 0.08037883, 0.05741328, 0.02163869, -0.03715056, -0.05842322, 
    -0.03269085, 0.01092894, -0.0002038628, -0.03103068, -0.1113692, 
    -0.1228276, -0.0565027, 0.06807411, 0.158927, 0.2347734, 0.2726477, 
    0.2849524, 0.2855384, 0.2649003, 0.1949946, 0.1481521, 0.09151185, 
    0.04748476, 0.003913999, -0.02048385, -0.09193552, -0.1642503, 
    -0.1074796, -0.1298754, 0.02212667, 0.129174, 0.2407629, 0.2543534, 
    0.2253169, 0.202335, 0.2328365, 0.2575598, 0.1748774, 0.1199296, 
    0.04276478, 0.03456163, -0.01171088, -0.07797068, -0.176099, -0.2317957, 
    -0.2537683, -0.1459233, 0.03072062, 0.1068925, 0.1390865, 0.1639562, 
    0.1467851, 0.08894002, -0.007560551, -0.04999214, 0.04409952, 0.1508378, 
    0.2670162, 0.3028719, 0.08425236, -0.1911056, -0.3443771, -0.3260665, 
    -0.2453047, -0.08732969, -0.080917, -0.1649827, -0.3416589, -0.6823167, 
    -0.762297, -0.9006434,
  -0.9920497, -0.8209071, -0.6048586, -0.3590256, -0.1735764, -0.08244681, 
    -0.0923264, -0.3394129, -0.6126223, -0.7705325, -0.824276, -0.8707769, 
    -0.7340742, -0.561125, -0.2959884, -0.1236902, 0.03070434, 0.1507076, 
    0.2461666, 0.3038, 0.2456783, 0.1580807, 0.09795702, 0.08122504, 
    0.1075923, 0.1192297, 0.1384355, 0.1288, 0.105981, 0.1313716, 0.1438554, 
    0.1439856, 0.1434157, 0.1522702, 0.1750404, 0.1887284, 0.2374589, 
    0.2667395, 0.2696204, 0.2076411, 0.1961178, 0.1162674, 0.06415153, 
    0.01042461, -0.03347194, -0.07495952, -0.1111412, -0.1495364, -0.1863202, 
    -0.1916589, -0.1723231, -0.1350675, -0.08412409, -0.009514093, 0.0439527, 
    0.1000242, 0.1258049, 0.1386304, 0.1293695, 0.08981872, 0.05974078, 
    0.0709548, 0.103035, -0.1441007, -0.1477137, -0.1503175, -0.1906822, 
    -0.2408777, -0.2937424, -0.2402755, -0.2532963, -0.2069747, -0.1321374, 
    -0.1463464, -0.1138757, -0.08399293, -0.06327349, -0.03633666, 
    0.06856242, 0.1844315, 0.2529701, 0.2305577, 0.201896, 0.009154916, 
    -0.2886968, -0.5774174, -0.7023035, -0.628557, -0.3021245, -0.02723813, 
    0.08109474, 0.03850058, -0.1356856, -0.3852625, -0.6835047, -0.9167402,
  -0.5827883, -0.4023522, -0.2829843, -0.1809497, -0.2507093, -0.3770597, 
    -0.4071541, -0.4296473, -0.5126711, -0.6479739, -0.7055426, -0.6469, 
    -0.4874108, -0.275334, -0.08098185, 0.07014132, 0.1719804, 0.2361732, 
    0.2585364, 0.2685623, 0.2767819, 0.259985, 0.2566156, 0.2432693, 
    0.2174393, 0.1656651, 0.1150793, 0.08363402, 0.03265738, 0.01437938, 
    0.03187609, 0.0442785, 0.07920682, 0.1073155, 0.145548, 0.1569901, 
    0.1421138, 0.1255611, 0.06179154, 0.001375079, -0.05360568, -0.105103, 
    -0.1629481, -0.1675377, -0.1268476, -0.07818222, -0.04170763, 
    0.0004961491, 0.02753067, 0.0432694, 0.06416774, 0.04398549, 0.02342868, 
    -0.02089095, -0.07108617, -0.1181239, -0.184188, -0.2532802, -0.3149825, 
    -0.3796636, -0.4269292, -0.4803306, -0.5240643, -0.5473554, -0.4985601, 
    -0.6371669, -0.6519128, -0.6425541, -0.6388921, -0.6207931, -0.5786544, 
    -0.5255619, -0.4801518, -0.3810633, -0.3396407, -0.2382735, -0.1642501, 
    -0.1169518, -0.05271077, -0.04768133, -0.002010822, -0.04447508, 
    -0.1890546, -0.3929121, -0.5507247, -0.6754155, -0.7385993, -0.6583591, 
    -0.4635668, -0.2577231, -0.087134, 0.005818069, -0.03794798, -0.1337976, 
    -0.2481368, -0.3574306,
  -0.1632409, -0.1862553, -0.1784103, -0.1397711, -0.2276779, -0.2212814, 
    -0.231991, -0.2208907, -0.2103763, -0.1825118, -0.1209396, -0.03309774, 
    0.06447715, 0.1631915, 0.2324784, 0.2837318, 0.3236243, 0.3399491, 
    0.3345942, 0.3037024, 0.2645096, 0.2128819, 0.1540117, 0.1216385, 
    0.1253332, -0.02071178, -0.04475117, -0.003947139, -0.02658725, 
    -0.02989125, -0.0216558, 0.002042055, 0.04842854, 0.09237421, 0.1267492, 
    0.142781, 0.1451085, 0.1532141, 0.1446528, 0.1230056, 0.1069248, 
    0.08306426, 0.06978297, 0.06530702, 0.06201941, 0.06735778, 0.06151474, 
    0.03622174, 0.01501435, -0.02644074, -0.07875198, -0.1438398, -0.2031986, 
    -0.2457118, -0.2942469, -0.33064, -0.3479578, -0.3646895, -0.3586023, 
    -0.3717859, -0.3874109, -0.4112228, -0.4374109, -0.4576095, -0.4783777, 
    -0.4823653, -0.481405, -0.4800053, -0.4587813, -0.4144291, -0.3490645, 
    -0.2586673, -0.1727462, -0.133114, -0.08783412, -0.06358278, -0.06089759, 
    -0.04613495, -0.08887589, -0.1699795, -0.2234136, -0.3336349, -0.4026777, 
    -0.4562261, -0.4966235, -0.5248299, -0.5168552, -0.486012, -0.4314213, 
    -0.3001876, -0.1560469, -0.06151581, -0.0407474, -0.05118042, 
    -0.07826376, -0.1179773,
  -0.09471884, -0.07447144, -0.04392132, -0.01221558, 0.009578019, 
    0.02868611, 0.04146278, 0.04597139, 0.06527478, 0.0857662, 0.1142817, 
    0.1442133, 0.1686438, 0.1824946, 0.1888423, 0.1772374, 0.1558344, 
    0.1325923, 0.1160231, 0.1003654, 0.08895588, 0.07879961, 0.06859457, 
    0.06395614, 0.07116652, 0.08368278, 0.08801222, 0.1160721, 0.1343664, 
    0.1638911, 0.1683507, 0.1685295, 0.1681226, 0.1690506, 0.1729732, 
    0.1614009, 0.1483963, 0.1279211, 0.1072016, 0.07678169, 0.04772902, 
    0.02674931, 0.01507938, -0.0002364218, -0.009464949, -0.01910034, 
    -0.02740115, -0.04177289, -0.06761923, -0.09981323, -0.126685, 
    -0.1541101, -0.1871342, -0.2237065, -0.2522547, -0.2927983, -0.3263106, 
    -0.3491622, -0.3700769, -0.3835535, -0.3961186, -0.4114018, -0.4194747, 
    -0.4269942, -0.4206629, -0.403394, -0.3761967, -0.3374923, -0.2725672, 
    -0.203866, -0.1353438, -0.07152539, -0.04369348, -0.02307177, 0.01380974, 
    0.03221804, 0.05435342, 0.05827595, 0.02425903, 0.003897697, 0.02782351, 
    0.009578109, -0.008813977, -0.04325402, -0.01561737, -0.1000086, 
    -0.1574631, -0.1813725, -0.2040612, -0.2272545, -0.2103114, -0.1949467, 
    -0.1611088, -0.1323979, -0.1188562, -0.1089441,
  -0.1181075, -0.08394408, -0.05718628, -0.0250411, 0.006664604, 0.0366939, 
    0.06525835, 0.09326935, 0.1134843, 0.1350826, 0.1561112, 0.175968, 
    0.1882564, 0.2003658, 0.2124263, 0.2142981, 0.2153073, 0.209106, 
    0.2055741, 0.2060949, 0.2014237, 0.1969153, 0.1913815, 0.1740963, 
    0.160815, 0.1586177, 0.1598384, 0.1503983, 0.140942, 0.1331131, 
    0.1179113, 0.1039789, 0.08815879, 0.07556117, 0.06136841, 0.04151163, 
    0.02989054, 0.01942506, 0.01540485, 0.01426554, 0.002937406, 
    -0.001229256, -0.03371623, -0.04994345, -0.0621993, -0.07053263, 
    -0.090129, -0.1039799, -0.1231694, -0.1396896, -0.1537846, -0.1742111, 
    -0.1948002, -0.212476, -0.232349, -0.2433353, -0.2617435, -0.2777267, 
    -0.2949141, -0.3152104, -0.3261479, -0.3405684, -0.3536381, -0.3544356, 
    -0.3586512, -0.360295, -0.3625248, -0.3591069, -0.3492924, -0.3478926, 
    -0.340422, -0.3284916, -0.329517, -0.3248458, -0.3187585, -0.3179936, 
    -0.318905, -0.3172449, -0.3211186, -0.3233484, -0.3248783, -0.3267176, 
    -0.3320398, -0.334644, -0.3375086, -0.3346765, -0.3285567, -0.3200606, 
    -0.3081303, -0.2878015, -0.2777267, -0.266366, -0.2487227, -0.2198491, 
    -0.190129, -0.1529871,
  -0.5371165, -0.5280833, -0.5187082, -0.5093009, -0.4997635, -0.48964, 
    -0.4781812, -0.4653886, -0.4503657, -0.4330805, -0.4126705, -0.3905514, 
    -0.367179, -0.3423417, -0.3150954, -0.2868564, -0.2574291, -0.2281158, 
    -0.1984284, -0.1682038, -0.1370354, -0.1043363, -0.06984758, -0.03244543, 
    0.00775671, 0.05145741, 0.09839773, 0.147584, 0.1972263, 0.2458262, 
    0.292099, 0.3350677, 0.3740325, 0.4077401, 0.4311616, 0.4499924, 
    0.4623294, 0.4669521, 0.4641525, 0.454517, 0.4388759, 0.4176356, 
    0.3911217, 0.3609133, 0.3275639, 0.2935472, 0.2572031, 0.199358, 
    0.165683, 0.1219816, 0.09162712, 0.05337858, -0.002416134, -0.08955765, 
    -0.04870462, -0.1296291, -0.1681871, -0.1906319, -0.1735253, -0.1297269, 
    -0.1488018, -0.2377186, -0.1752505, -0.188077, -0.1793528, -0.1765857, 
    -0.1720123, -0.1750398, -0.175544, -0.1674223, -0.1675854, -0.1694083, 
    -0.1739655, -0.1623931, -0.1320219, -0.1856194, -0.1250238, -0.311286, 
    -0.2423244, -0.2827215, -0.308845, -0.3385487, -0.3657947, -0.3984609, 
    -0.4284577, -0.4555249, -0.4805732, -0.502286, -0.5210519, -0.5363841, 
    -0.5474358, -0.5542555, -0.5552154, -0.5545635, -0.5517802, -0.5455313,
  -0.2477454, -0.2452226, -0.2453852, -0.2442947, -0.2407466, -0.2348221, 
    -0.2300044, -0.2277583, -0.2289464, -0.2327225, -0.2376866, -0.2425857, 
    -0.2466708, -0.2496984, -0.2502846, -0.2480874, -0.2445065, -0.2415116, 
    -0.2375565, -0.2421625, -0.2467031, -0.2546134, -0.2576406, -0.2516022, 
    -0.2286687, -0.188776, -0.1352611, -0.0740633, -0.008779049, 0.05814791, 
    0.1237888, 0.1837826, 0.2335711, 0.2716079, 0.2966242, 0.3085217, 
    0.308815, 0.3003507, 0.2856531, 0.2661874, 0.2405682, 0.2146571, 
    0.1951421, 0.1727786, 0.1615484, 0.1740971, 0.148577, 0.1579843, 
    0.1695242, 0.193352, 0.1900158, 0.2260351, 0.1703866, 0.1713471, 
    0.1249113, 0.1165462, 0.05241871, -0.03869486, -0.1461167, -0.25489, 
    -0.3394923, -0.41752, -0.4493892, -0.4516346, -0.4320714, -0.4047767, 
    -0.3811274, -0.360408, -0.3671952, -0.3754959, -0.3827388, -0.3423581, 
    -0.2780676, -0.2084551, -0.1364987, -0.09053528, -0.04559684, 
    -0.03101349, 0.005640209, 0.004549503, -0.02394938, -0.03973722, 
    -0.02175188, -0.02915764, -0.06166029, -0.07199574, -0.07603216, 
    -0.09977865, -0.130394, -0.160944, -0.1896882, -0.2148023, -0.2314687, 
    -0.240567, -0.2458248, -0.2483311,
  0.01967013, -0.03607534, -0.0581131, -0.05804789, -0.05109817, -0.04925895, 
    -0.04654086, -0.04514104, -0.04304141, -0.03526154, -0.0213618, 
    -0.001700327, 0.01613826, 0.0265547, 0.03259325, 0.03265905, 0.01664352, 
    -0.02642345, -0.09182024, -0.1678133, -0.2376699, -0.2691803, -0.2548254, 
    -0.2448481, -0.2663325, -0.3240151, -0.3816646, -0.4042557, -0.3845456, 
    -0.332999, -0.2696688, -0.2025461, -0.1426344, -0.09282923, -0.06398821, 
    -0.05611038, -0.05178356, -0.03456306, -0.001782417, 0.0426836, 
    0.09401703, 0.1423922, 0.1115327, 0.1309988, 0.08908725, 0.07985878, 
    0.06039286, 0.06234588, 0.06296438, 0.06159717, 0.06369677, 0.07168841, 
    0.09123588, 0.1100998, 0.09650898, 0.0620203, -0.01797652, -0.1547279, 
    -0.3419998, -0.5307693, -0.6999425, -0.8127518, -0.8628818, -0.848429, 
    -0.8066482, -0.7473058, -0.68562, -0.610392, -0.5231848, -0.4236079, 
    -0.3228755, -0.2216549, -0.125756, -0.04658985, 0.01280141, 0.04147995, 
    0.07066298, 0.08951056, 0.0949468, 0.1143153, 0.120012, 0.1186122, 
    0.113127, 0.135295, 0.1692955, 0.2200119, 0.2494066, 0.3164642, 
    0.3272395, 0.2151136, 0.29498, 0.2367277, 0.2112398, 0.1886482, 
    0.1416759, 0.08496952,
  0.2850518, 0.2492278, 0.1798105, 0.1132739, 0.04790902, -0.02043414, 
    -0.08475721, -0.1123123, -0.08351994, -0.03161561, 0.01812387, 
    0.04838105, 0.06032759, 0.05288959, 0.02300656, -0.01602328, -0.08127391, 
    -0.1708899, -0.2431059, -0.2925687, -0.2885652, -0.3246002, -0.3486719, 
    -0.3875725, -0.4257564, -0.4358962, -0.4890378, -0.5278071, -0.5132893, 
    -0.4932208, -0.487345, -0.4856035, -0.483569, -0.4802002, -0.4842362, 
    -0.5179272, -0.5824776, -0.6559973, -0.7283278, -0.7276936, -0.6218357, 
    -0.4210052, -0.2060308, 0.002059937, 0.1261163, 0.0724051, -0.09610128, 
    -0.2027423, -0.2864658, -0.3636632, -0.3809484, -0.3562902, -0.2845617, 
    -0.1758865, -0.05091912, 0.02391791, -0.05996895, 0.05581999, 
    -0.09486389, -0.2888417, -0.4715569, -0.6879308, -0.8024485, -0.9159744, 
    -0.9572504, -0.9245353, -0.8384023, -0.7065175, -0.5829334, -0.4703848, 
    -0.3644114, -0.2758052, -0.2065506, -0.1320879, -0.1168209, -0.1093501, 
    -0.1060785, -0.08916771, -0.05277456, 0.007853699, 0.145663, 0.2695236, 
    0.3671636, 0.4568608, 0.4962977, 0.4860438, 0.408163, 0.3239018, 
    0.2008874, 0.1985281, 0.187737, 0.289104, 0.2938085, 0.3322682, 
    0.3654065, 0.3299246,
  0.00494051, 0.09431267, 0.07577324, 0.1525159, 0.1047292, 0.1075611, 
    0.04333591, -0.01699877, -0.1599836, -0.1682196, -0.2198639, -0.1996174, 
    -0.1286368, -0.05881262, -0.02741647, 0.03303266, 0.0878346, 0.0873301, 
    0.09878793, 0.0562911, 0.03052711, -0.1258049, -0.3047943, -0.4079657, 
    -0.4520898, -0.429955, -0.3837805, -0.3520255, -0.3486404, -0.3719149, 
    -0.4178455, -0.4650953, -0.4616125, -0.4258217, -0.4101474, -0.4419346, 
    -0.5240473, -0.6401117, -0.783048, -0.9088132, -0.9501542, -0.8918369, 
    -0.7037342, -0.4818268, -0.2453034, -0.05427194, -0.1182858, -0.1311438, 
    -0.2827066, -0.4228594, -0.5195715, -0.5587477, -0.5436763, -0.4902744, 
    -0.4181066, -0.318188, -0.2003494, -0.1358474, -0.1227779, -0.1731685, 
    -0.2489332, -0.3836176, -0.5447991, -0.6679438, -0.7718501, -0.8124588, 
    -0.8286861, -0.8069575, -0.7253656, -0.6832922, -0.7399001, -0.5142982, 
    -0.3254148, -0.1156491, 0.09455585, 0.2813239, 0.3430753, 0.4857834, 
    0.4315679, 0.40328, 0.435116, 0.5608484, 0.6995692, 0.8901128, 1.039641, 
    1.133358, 1.135165, 1.073918, 0.942961, 0.767782, 0.6232188, 0.2208261, 
    0.2797947, 0.2635026, 0.194427, 0.06563425,
  -0.06415081, -0.02907562, -0.2733626, -0.4121809, -0.339118, -0.2782617, 
    -0.2144113, -0.2722237, -0.3889394, -0.4782948, -0.5284905, -0.4838281, 
    -0.2812572, -0.09338284, 0.003834724, 0.04305887, 0.1559657, 0.146965, 
    0.1706629, 0.1026613, 0.0207448, 0.001815796, 0.1577077, 0.1500893, 
    0.1485424, 0.1368723, 0.1034584, 0.07883358, 0.09343338, 0.1368408, 
    0.1549406, 0.1043224, -0.01599026, -0.09629536, -0.168366, -0.2164135, 
    -0.252758, -0.2816477, -0.2690012, -0.2650464, -0.2359445, -0.1993237, 
    -0.148982, -0.06826949, -0.03631955, 0.02834523, 0.04494679, 0.06109279, 
    0.01475453, -0.05993629, -0.106209, -0.147241, -0.203019, -0.2185953, 
    -0.1870358, -0.1526119, -0.09024215, 0.03129113, 0.1892501, 0.2474205, 
    0.2873131, 0.2672449, 0.22592, 0.1470789, 0.03225124, -0.04724085, 
    -0.09767997, -0.07980889, -0.02504009, 0.05336159, 0.1449957, 0.202027, 
    0.1975185, 0.2241786, 0.3146896, 0.4450933, 0.6020594, 0.6828048, 
    0.5736089, 0.6901128, 0.5947841, 0.5670985, 0.6597255, 0.8526454, 
    1.052173, 1.157919, 1.207724, 1.204891, 1.198349, 1.17802, 1.120679, 
    0.9780032, 0.8153732, 0.5903571, 0.3760996, 0.1599863,
  0.994133, 0.7690026, 0.5086675, 0.308814, 0.1656504, 0.04611921, 
    -0.03281951, -0.0222733, 0.1191978, 0.3842206, 0.7404871, 1.024194, 
    0.9233971, 0.526669, 0.08500266, -0.2913971, -0.5046458, -0.6469479, 
    -0.6371822, -0.5011142, -0.2915602, -0.06389129, 0.1055748, 0.1793056, 
    0.246412, 0.2507091, 0.2566009, 0.2512784, 0.3489509, 0.4683197, 
    0.5187428, 0.6751561, 0.8124604, 0.8245211, 0.7597585, 0.6071222, 
    0.2157316, -0.01250696, -0.2142975, -0.2503326, -0.1158111, -0.0829339, 
    -0.050138, 0.1642663, 0.3342045, 0.5521408, 0.6662847, 0.7489831, 
    0.7930424, 0.8102629, 0.8349049, 0.922828, 1.026408, 1.16705, 1.254583, 
    1.323918, 1.427255, 1.494752, 1.579159, 1.61246, 1.569345, 1.481405, 
    1.395972, 1.339202, 1.30621, 1.336728, 1.348463, 1.28899, 1.164104, 
    1.079973, 1.096102, 1.177808, 1.249976, 1.298203, 1.311858, 1.386191, 
    1.549228, 1.81954, 1.946949, 1.936207, 1.268498, 0.9081465, 0.859807, 
    0.9867601, 1.234156, 1.425465, 1.520143, 1.511923, 1.519947, 1.511418, 
    1.470142, 1.375285, 1.282951, 1.221998, 1.231454, 1.162639,
  2.217652, 2.151392, 2.063909, 2.03287, 1.99384, 2.011939, 2.009025, 
    1.987476, 1.972518, 1.97981, 2.088762, 2.239234, 2.348593, 2.291822, 
    2.0733, 1.765536, 1.498235, 1.309563, 1.170484, 1.089348, 1.078167, 
    1.151702, 1.176734, 1.06124, 0.9889088, 0.9753668, 0.984953, 1.028817, 
    1.015487, 1.042342, 1.121721, 1.277629, 1.560686, 1.867164, 2.113062, 
    2.213029, 2.165862, 2.014657, 1.868905, 1.695989, 1.536956, 1.424146, 
    1.350986, 1.35538, 1.433668, 1.59555, 1.780869, 2.001343, 2.155396, 
    2.233668, 2.236142, 2.194361, 2.189674, 2.222974, 2.326506, 2.471054, 
    2.62317, 2.797779, 2.920142, 2.979745, 3.044035, 3.06954, 2.973983, 
    2.764185, 2.559286, 2.405038, 2.236044, 1.998805, 1.702548, 1.427385, 
    1.193596, 1.052157, 1.029989, 1.027401, 1.015813, 1.04078, 1.198577, 
    1.488941, 1.781471, 1.930184, 1.919068, 1.8983, 2.008277, 1.921184, 
    1.975676, 2.218564, 2.462851, 2.624163, 2.651197, 2.591138, 2.532023, 
    2.455298, 2.348381, 2.192945, 2.16941, 2.210149,
  1.721885, 1.678818, 1.684466, 1.722096, 1.734108, 1.754177, 1.835118, 
    1.950547, 1.963616, 1.830478, 1.616985, 1.459319, 1.436532, 1.493123, 
    1.525888, 1.506795, 1.468009, 1.421883, 1.336418, 1.24524, 1.224715, 
    1.292457, 1.372014, 1.428314, 1.436646, 1.404989, 1.357463, 1.267718, 
    1.114593, 0.9941015, 0.9494562, 0.9828219, 1.060133, 1.179485, 1.380413, 
    1.662038, 1.914968, 2.128412, 2.266612, 2.297325, 2.276133, 2.221332, 
    2.167344, 2.17278, 2.193011, 2.199896, 2.229046, 2.288193, 2.407497, 
    2.57553, 2.730723, 2.848578, 2.981358, 3.200123, 3.418304, 3.539283, 
    3.595533, 3.657855, 3.712135, 3.724619, 3.768596, 3.806862, 3.758831, 
    3.571331, 3.311566, 3.025026, 2.686369, 2.314576, 1.981861, 1.703915, 
    1.490781, 1.298674, 1.117424, 0.9414644, 0.8297133, 0.7958918, 0.7863379, 
    0.7660904, 0.8264747, 1.040928, 1.320078, 1.519379, 1.562542, 1.506569, 
    1.548171, 1.692636, 1.895176, 2.079503, 2.168499, 2.196364, 2.209304, 
    2.220127, 2.189919, 2.100498, 1.962787, 1.816986,
  1.624668, 1.550546, 1.55551, 1.600872, 1.610751, 1.586728, 1.583179, 
    1.57784, 1.56915, 1.563535, 1.539444, 1.499146, 1.473249, 1.449697, 
    1.387815, 1.285391, 1.220156, 1.213548, 1.212767, 1.197743, 1.165339, 
    1.131159, 1.131533, 1.161465, 1.198021, 1.217715, 1.253148, 1.256567, 
    1.208471, 1.159303, 1.157707, 1.192295, 1.242978, 1.321738, 1.425644, 
    1.539169, 1.652369, 1.790894, 1.929093, 2.040439, 2.088665, 2.092652, 
    2.109742, 2.166659, 2.226995, 2.216969, 2.164494, 2.109839, 2.104404, 
    2.246558, 2.505039, 2.672372, 2.720225, 2.82322, 3.025758, 3.178395, 
    3.249505, 3.318938, 3.412314, 3.458457, 3.508994, 3.6025, 3.650123, 
    3.52579, 3.36067, 3.173024, 2.876523, 2.42942, 1.994264, 1.645159, 
    1.328346, 1.069638, 0.9101334, 0.832448, 0.832171, 0.8434176, 0.76194, 
    0.5550222, 0.3323984, 0.3106537, 0.4774995, 0.6571217, 0.7678151, 
    0.8016529, 0.8651457, 0.9720469, 1.087769, 1.242831, 1.439185, 1.629224, 
    1.784173, 1.905559, 1.978881, 1.990975, 1.902548, 1.755706,
  1.463826, 1.433764, 1.408587, 1.340487, 1.220418, 1.100514, 1.068532, 
    1.053785, 0.9915438, 0.9505301, 0.9423571, 0.9419832, 0.9670811, 1.0156, 
    1.103408, 1.252154, 1.38194, 1.400022, 1.306565, 1.213303, 1.162473, 
    1.105507, 0.9933643, 0.8787975, 0.8582573, 0.9250059, 1.040485, 1.117112, 
    1.051261, 0.89042, 0.7941322, 0.7783279, 0.8183661, 0.915225, 0.9751205, 
    0.9312572, 0.8972073, 0.9658442, 1.10559, 1.318498, 1.540145, 1.624959, 
    1.639462, 1.743969, 1.812899, 1.765568, 1.71845, 1.704844, 1.622715, 
    1.606097, 1.758668, 1.862721, 1.764267, 1.631195, 1.673089, 1.852565, 
    2.021348, 2.153802, 2.325058, 2.467392, 2.540049, 2.598431, 2.621738, 
    2.532122, 2.467929, 2.503753, 2.409726, 2.099456, 1.674489, 1.305202, 
    1.009694, 0.7746191, 0.5758886, 0.4294534, 0.3584409, 0.3259535, 
    0.1638274, 0.09128571, 0.06187439, -0.018888, -0.09981203, -0.04611731, 
    0.04654264, 0.09900045, 0.1753826, 0.3404703, 0.4867096, 0.5678959, 
    0.6886969, 0.8859615, 1.103832, 1.305363, 1.447159, 1.500886, 1.506552, 
    1.498495,
  0.9211826, 0.8786211, 0.7871819, 0.6989508, 0.6672935, 0.6144948, 
    0.5711846, 0.55831, 0.5254645, 0.5183358, 0.5287366, 0.5202403, 
    0.5750093, 0.6682062, 0.6960707, 0.774601, 0.9370184, 1.00323, 0.9690666, 
    0.9341869, 0.9211655, 0.8477106, 0.6865463, 0.569129, 0.5627327, 
    0.5846567, 0.5893459, 0.6267967, 0.677659, 0.6582575, 0.6584368, 
    0.6705799, 0.6532297, 0.6004133, 0.519474, 0.4701729, 0.4777098, 
    0.4240303, 0.3373613, 0.3503981, 0.4839916, 0.5887785, 0.7314382, 
    0.9947352, 1.179762, 1.133994, 1.067441, 1.039186, 0.9077897, 0.7925715, 
    0.7881284, 0.7390232, 0.5496845, 0.3067641, 0.2340593, 0.3962989, 
    0.5900159, 0.7106543, 0.8590102, 1.017914, 1.070078, 1.031781, 1.041091, 
    1.068777, 1.17169, 1.340911, 1.449115, 1.438975, 1.351491, 1.205788, 
    1.041514, 0.8323832, 0.5398698, 0.2624445, 0.1199155, -0.03573275, 
    -0.1880281, -0.1603911, -0.227839, -0.5236564, -0.742764, -0.6399975, 
    -0.5312572, -0.4916415, -0.341918, -0.1060624, 0.06582928, 0.1310949, 
    0.1207914, 0.1117907, 0.1673908, 0.313386, 0.4616117, 0.6498928, 
    0.845108, 0.9313231,
  0.2121506, 0.2874918, 0.2876554, 0.3120861, 0.4298759, 0.5044847, 
    0.4773855, 0.3513117, 0.1233983, 0.02583933, 0.061728, 0.07636023, 
    0.1629162, 0.3242769, 0.4393163, 0.5661879, 0.7430267, 0.8794198, 
    0.8870859, 0.8080983, 0.6838779, 0.4743395, 0.2486238, 0.07077503, 
    0.02575493, 0.1055889, 0.1518135, 0.2022696, 0.2552805, 0.1722078, 
    0.06987953, 0.03581429, 0.02129555, 0.04450798, 0.03257751, -0.02468204, 
    -0.135684, -0.2978754, -0.3506432, -0.2611561, -0.2161531, -0.268692, 
    -0.2971253, -0.144733, -0.003050327, -0.01538754, -0.01452541, 0.1487727, 
    0.05595016, -0.05339241, -0.05124378, -0.1286206, -0.2735419, -0.3966379, 
    -0.5615797, -0.5912833, -0.5203848, -0.4870348, -0.4598379, -0.3913321, 
    -0.2925854, -0.2171946, -0.1933665, -0.109138, -0.008242607, 0.0492115, 
    0.207058, 0.4196553, 0.5878358, 0.6176367, 0.5051208, 0.383018, 
    0.1202083, -0.2394271, -0.43155, -0.6514554, -0.8333731, -0.7078362, 
    -0.6812735, -0.888484, -0.9482818, -0.8895254, -1.005346, -1.1177, 
    -1.025056, -0.8923249, -0.7780833, -0.6507888, -0.6055093, -0.6069579, 
    -0.5011969, -0.3403721, -0.2326097, -0.1247311, 0.00747776, 0.109334,
  -0.4225006, -0.3326569, -0.1484447, -0.04308987, -0.1184311, -0.2829337, 
    -0.366478, -0.2797599, -0.2164624, -0.1337636, 0.04556561, 0.2410736, 
    0.4029715, 0.4332449, 0.4177175, 0.4031506, 0.274277, 0.1801853, 
    0.1293874, 0.03890896, -0.0006575584, -0.08024788, -0.2237864, 
    -0.3990469, -0.5859609, -0.5193758, -0.3750076, -0.2728591, -0.1665435, 
    -0.24405, -0.3395252, -0.3948965, -0.4900136, -0.4401436, -0.4216213, 
    -0.5942779, -0.7688866, -0.8698635, -0.9443755, -0.9769764, -0.9128165, 
    -0.9856839, -1.204483, -1.225707, -1.053197, -0.9214585, -0.8198152, 
    -0.7033601, -0.8249581, -0.9743557, -0.9502025, -1.022924, -1.132152, 
    -1.170254, -1.288109, -1.42141, -1.495417, -1.516039, -1.51459, 
    -1.549909, -1.530996, -1.403376, -1.348184, -1.352156, -1.305785, 
    -1.17128, -0.8983307, -0.6742091, -0.4908757, -0.3693423, -0.3723211, 
    -0.2947502, -0.2981029, -0.5145903, -0.6967192, -0.9574776, -1.190812, 
    -1.081893, -1.016234, -0.9767487, -1.141251, -1.304076, -1.52364, 
    -1.695189, -1.768757, -1.703669, -1.485424, -1.165209, -0.9726806, 
    -0.9425201, -0.9031811, -0.8560615, -0.792748, -0.7147207, -0.6238194, 
    -0.5075264,
  -0.6863189, -0.8093162, -0.8015368, -0.8577058, -0.9598222, -0.9918208, 
    -1.028588, -0.8799232, -0.5810137, -0.3666255, -0.2592365, -0.2267169, 
    -0.2134519, -0.3145258, -0.4569411, -0.563468, -0.7905027, -0.912573, 
    -0.8809974, -0.9538325, -0.9260979, -0.9833407, -1.013647, -0.8644116, 
    -0.8669829, -0.842813, -0.8208239, -0.8138742, -0.6749742, -0.7989655, 
    -0.9677639, -1.018431, -1.169701, -1.162686, -1.134952, -1.264265, 
    -1.166007, -0.8400469, -0.8413491, -1.007837, -0.9965568, -1.296996, 
    -1.593725, -1.713761, -1.580591, -1.414542, -1.419604, -1.477563, 
    -1.59366, -1.731372, -1.708097, -1.713175, -1.774894, -1.858097, 
    -2.088289, -2.248673, -2.353409, -2.447452, -2.34724, -2.291755, 
    -2.291251, -2.110115, -1.90445, -1.716169, -1.536482, -1.3031, 
    -0.9823639, -0.7809968, -0.7434313, -0.8169017, -0.9482002, -0.955476, 
    -0.8762116, -0.903995, -0.9728752, -0.9606199, -0.7952875, -0.6232825, 
    -0.8972406, -0.7335526, -0.5629471, -0.8987057, -1.242406, -1.501684, 
    -1.682966, -1.661238, -1.618839, -1.477383, -1.244098, -1.088337, 
    -1.067276, -1.124486, -1.099275, -0.928051, -0.7679758, -0.660017,
  -0.9092852, -1.039901, -1.120971, -1.063956, -0.7385818, -0.3105382, 
    -0.2958573, -0.3885984, -0.4575433, -0.5465083, -0.5050694, -0.720548, 
    -0.955753, -0.9585363, -1.079516, -1.295288, -1.475838, -1.599828, 
    -1.537035, -1.503149, -1.339575, -1.174763, -1.227156, -1.115926, 
    -1.13256, -1.234334, -1.306811, -1.443871, -1.466788, -1.59838, -1.49213, 
    -1.077416, -1.034887, -0.8972081, -0.8166904, -0.754337, -0.7662835, 
    -0.6643794, -0.6250238, -0.7913487, -1.021866, -1.549047, -1.631111, 
    -1.626033, -1.687377, -1.565633, -1.540502, -1.596313, -1.648494, 
    -1.776928, -1.867097, -1.89768, -1.887182, -1.933487, -2.21573, 
    -2.422078, -2.481941, -2.656193, -2.573673, -2.331241, -2.250936, 
    -2.09213, -1.903963, -1.598201, -1.273478, -1.128279, -1.036336, 
    -0.9757401, -1.052774, -1.26241, -1.328523, -1.362247, -1.351717, 
    -1.161157, -1.09768, -0.9268304, -0.2865474, -0.04553175, -0.5849198, 
    -0.4953689, -0.2558181, -0.5345129, -0.7438065, -1.10017, -1.328979, 
    -1.196118, -1.109253, -1.175284, -1.200415, -1.154793, -1.111775, 
    -0.9981849, -0.9978591, -1.023299, -0.9916741, -0.9441643,
  -1.009757, -1.035554, -0.9966546, -0.6874914, -0.2404863, -0.02048302, 
    0.09398645, -0.07129669, -0.3984614, -0.6896398, -0.817537, -0.9520254, 
    -1.134903, -1.225447, -1.113045, -1.097175, -1.113484, -1.228816, 
    -1.177953, -1.203555, -1.304581, -1.16835, -1.162263, -1.181762, 
    -1.267341, -1.400382, -1.425951, -1.438614, -1.464591, -1.493757, 
    -1.197305, -0.8918207, -0.927742, -0.9463779, -0.9145583, -0.6485428, 
    -0.5253657, -0.5854567, -0.6778723, -0.7589922, -0.9732171, -1.484399, 
    -1.624226, -1.727709, -1.812605, -1.655541, -1.45808, -1.220336, 
    -1.063109, -1.024698, -1.080671, -1.287068, -1.467553, -1.575724, 
    -1.703002, -1.828132, -1.820857, -1.884708, -1.878735, -1.71215, 
    -1.599129, -1.43767, -1.372631, -1.394506, -1.387215, -1.374568, 
    -1.387052, -1.331876, -1.106486, -1.071053, -1.00476, -0.9785558, 
    -1.04353, -0.8846267, -0.6713619, -0.4055413, 0.009204507, 0.3098882, 
    -0.07899526, -0.3777096, -0.1941484, -0.1836015, -0.2725335, -0.4001378, 
    -0.7028721, -0.7674394, -0.5924717, -0.6711826, -0.8784906, -0.8349847, 
    -0.8767003, -0.7968338, -0.7563878, -0.8921301, -0.9366613, -0.9826576,
  -0.6469474, -0.5135486, -0.3241446, -0.05314875, -0.02504009, -0.157804, 
    -0.1247637, -0.3378495, -0.4383376, -0.4901932, -1.017651, -0.8908441, 
    -0.7489655, -0.8813553, -0.8265696, -0.7645569, -0.7049708, -0.7273669, 
    -0.7631903, -0.8346906, -1.041788, -1.021735, -0.8910065, -0.9306707, 
    -1.037067, -1.097451, -1.135016, -1.102676, -0.9180408, -0.7108307, 
    -0.3891997, -0.2648509, -0.4046946, -0.5424876, -0.6653395, -0.5495842, 
    -0.3541253, -0.3214922, -0.4505441, -0.5780833, -0.7871332, -0.926537, 
    -1.014704, -1.35686, -1.459202, -1.222208, -1.078018, -0.8783927, 
    -0.7584705, -0.6672273, -0.7520418, -0.9279208, -1.009154, -1.091218, 
    -1.031843, -1.008926, -0.902009, -0.8907785, -1.065339, -1.119393, 
    -1.096492, -1.018611, -0.9963619, -1.126489, -1.329435, -1.382738, 
    -1.26075, -1.180053, -0.8645256, -0.7081292, -0.6699452, -0.6821523, 
    -0.6975169, -0.5603588, -0.2141676, 0.3025149, 0.31814, 0.2510338, 
    -0.1079996, -0.3436764, -0.1212969, 0.07051647, -0.07637477, -0.07375455, 
    -0.1749427, -0.4453528, -0.432071, -0.4279861, -0.5627027, -0.4495354, 
    -0.5269279, -0.5419021, -0.4603424, -0.5429759, -0.6288319, -0.671345,
  0.02483082, 0.06597567, 0.186028, 0.258, -0.06686974, -0.2382727, 
    -0.2378006, -0.5073152, -0.391593, -0.1305742, -0.3673418, -0.376261, 
    -0.1430739, -0.2136471, -0.3038645, -0.4548407, -0.5051498, -0.4425855, 
    -0.5081453, -0.5789785, -0.5867581, -0.5857983, -0.4419017, -0.4428296, 
    -0.6045485, -0.6478586, -0.5614491, -0.5417547, -0.3459539, -0.1006904, 
    0.03060818, 0.03500271, -0.2358789, -0.2856846, -0.3264718, -0.1992421, 
    -0.1146231, -0.1522045, -0.2552156, -0.382494, -0.5163474, -0.4394927, 
    -0.4194727, -0.8455305, -1.143415, -1.01153, -0.7060127, -0.5145416, 
    -0.4946523, -0.2823801, -0.2405019, -0.3422756, -0.3408113, -0.2970285, 
    -0.1890373, -0.1867747, -0.2044671, -0.2757721, -0.3280182, -0.3757234, 
    -0.4763417, -0.6155019, -0.7204335, -0.8155184, -0.8866446, -0.8513579, 
    -0.6544666, -0.5218329, -0.4617257, -0.4516182, -0.3881259, -0.4023671, 
    -0.3205638, -0.1113839, 0.01307869, 0.4225183, 0.4265873, 0.1769125, 
    -0.2205968, -0.3031815, -0.1245844, -0.1071198, -0.1503162, 0.01718044, 
    -0.04011154, -0.2926022, -0.2930899, -0.1555567, -0.1424708, -0.1764226, 
    -0.1450262, -0.1399317, -0.1157293, -0.07502317, -0.1064196, -0.05420637,
  0.436923, 0.4066496, 0.313143, 0.2371503, -0.1608799, -0.1858799, 
    -0.01590967, -0.2590077, -0.3494539, -0.07686317, 0.1967534, 0.3745041, 
    0.01428258, -0.2725661, -0.2422597, -0.314671, -0.4611235, -0.5943432, 
    -0.4578199, -0.4508533, -0.5013256, -0.4722075, -0.3211007, -0.1880608, 
    -0.1790924, -0.1424389, -0.02772522, -0.0480051, -0.007949352, 0.208375, 
    0.3013277, 0.3294697, 0.2992115, 0.1751068, -0.02012396, -0.04556417, 
    -0.0115633, 0.1071224, 0.06897068, 0.0410738, -0.06047249, -0.01141644, 
    -0.08884192, -0.2871485, -0.5544662, -0.7227287, -0.6087475, -0.3255606, 
    -0.116446, 0.1510997, 0.2423272, 0.2435155, 0.2682714, 0.3179288, 
    0.3982353, 0.3218517, 0.1274018, -0.0651927, -0.0363512, -0.172842, 
    -0.3131256, -0.4197659, -0.4426503, -0.4224834, -0.3624907, -0.3202538, 
    -0.3234277, -0.2434964, -0.2534571, -0.234056, -0.2521715, -0.2866116, 
    -0.2158918, -0.08286762, -0.02163792, 0.3042239, 0.2955002, 0.08492082, 
    -0.158227, -0.1625401, -0.1164953, -0.2425852, -0.05806422, 0.06221628, 
    -0.0308013, -0.1456614, -0.05962563, -0.05441809, 0.1019297, 0.1684499, 
    0.1147876, 0.09515905, 0.1847095, 0.2625251, 0.2912035, 0.3583751,
  0.4611421, 0.358391, 0.200334, 0.3168055, 0.1392826, -0.02886486, 
    0.1034753, 0.008163452, -0.007201672, 0.06228077, 0.1085861, 0.5935308, 
    0.2774835, -0.1028061, 0.1007576, 0.08643532, 0.04908133, -0.1935458, 
    -0.08954096, -0.1452055, -0.3415599, -0.2977772, -0.109951, -0.03806019, 
    0.03650045, 0.4403577, 0.6773038, 0.6921968, 0.6069589, 0.6067476, 
    0.5913177, 0.5987072, 0.7426686, 0.7265878, 0.385963, 0.2624605, 
    0.1880624, 0.185019, 0.2521415, 0.3296967, 0.2339125, 0.2217059, 
    0.09351587, -0.02723694, -0.1616607, -0.293334, -0.3635654, -0.3668857, 
    -0.1043205, 0.3261158, 0.4026461, 0.3522882, 0.2616625, 0.1013441, 
    0.07738543, 0.1586356, 0.2288179, 0.1091242, 0.16959, 0.1140714, 
    0.09750271, -0.008698463, -0.1524, -0.1752515, -0.1486888, -0.1268463, 
    -0.1644115, -0.1165109, -0.1238842, -0.09527111, -0.1996975, -0.1456447, 
    -0.05777025, -0.1629629, -0.1173251, 0.08145396, 0.1320721, -0.1432369, 
    -0.06291443, 0.02222544, 0.04198456, -0.08548951, 0.03519738, 0.0342865, 
    0.08013606, 0.01537371, 0.2022715, 0.1039968, 0.07753181, 0.2687917, 
    0.291904, 0.2519946, 0.3452892, 0.3033295, 0.4073668, 0.4698496,
  0.3161712, 0.2388108, 0.2060794, 0.3683191, 0.4373457, 0.1657803, 0.19314, 
    0.2360117, 0.1236417, 0.127857, -0.1001215, 0.3817466, 0.4267187, 
    0.1842051, 0.5306406, 0.4825938, 0.7227144, 0.7535248, 0.7514091, 
    0.6658456, 0.5440848, 0.3067634, 0.449244, 0.5754807, 0.4686778, 
    0.7862394, 0.953167, 0.9365489, 0.6695893, 0.6707287, 0.810312, 
    0.7530694, 0.7825613, 0.7197032, 0.6716399, 0.8315682, 0.7097259, 
    0.4762955, 0.2266687, 0.08369994, 0.1090424, 0.2258554, 0.1355071, 
    -0.06517673, -0.2988682, -0.3579178, -0.2914302, -0.4571528, -0.6669505, 
    -0.2602937, 0.06333923, 0.09174156, 0.09968376, -0.1305084, -0.3395252, 
    -0.347012, -0.1046453, -0.1101632, -0.04440832, 0.04878855, 0.1416273, 
    0.1051521, -0.09797239, -0.1924715, -0.1969471, -0.1575103, -0.09094143, 
    -0.04667044, -0.1006742, -0.08887386, -0.09722376, -0.1687403, 
    -0.1666412, -0.1407623, -0.05720162, 0.07684784, 0.01434779, -0.1439204, 
    -0.0513097, 0.004191577, -0.08765399, -0.01258904, 0.0364182, 0.06701732, 
    0.06018186, 0.0967052, 0.08273959, 0.1473403, 0.1331959, 0.3529229, 
    0.624505, 0.495029, 0.463861, 0.5336032, 0.4657154, 0.3750257,
  0.3872485, 0.2421958, 0.3021083, 0.2918217, 0.6926355, 0.4747481, 
    0.2428473, 0.6123295, 0.498821, 0.2655365, 0.2183516, 0.4194259, 
    0.6305751, 0.4886158, 0.4977298, 0.4541427, 0.6050377, 0.8135988, 
    0.991724, 0.9094163, 0.8531662, 0.6476161, 0.5013596, 0.4550054, 
    0.4586349, 0.6029872, 0.6260012, 0.6084723, 0.1474861, 0.2751713, 
    0.5964444, 0.7005787, 0.5869396, 0.6194263, 0.7871667, 0.6040289, 
    0.2126875, 0.06244354, 0.06416881, 0.12815, 0.2031335, 0.04294479, 
    -0.22408, -0.2105709, -0.2842688, -0.7032955, -0.7238846, -0.4822178, 
    -0.6908766, -0.5810947, -0.251863, -0.2167065, -0.08005261, -0.05728245, 
    -0.1633534, -0.2675691, -0.189167, -0.1678782, -0.1894927, -0.1928287, 
    -0.07474661, 0.01379538, -0.007607937, -0.007639885, 0.03392887, 
    0.04992819, -0.01429701, -0.07884789, -0.05265999, -0.08889055, 
    -0.03472424, -0.003587961, 0.09934139, 0.19856, 0.1463792, 0.1153081, 
    -0.09745252, 0.08005422, 0.02455291, 0.006991148, -0.0391677, 
    -0.09468532, -0.09621543, 0.06228089, 0.1361088, 0.03303266, -0.04613411, 
    0.08949494, 0.2268972, 0.2986095, 0.6884859, 0.6282644, 0.5134695, 
    0.672291, 0.5400319, 0.450253,
  0.2749923, 0.1815842, 0.3004156, 0.1829351, 0.2008876, 0.1801519, 
    0.0177007, 0.1462651, 0.3562421, 0.4186934, 0.5384686, 0.03872935, 
    0.251148, 0.5800054, 0.4791102, 0.3361089, 0.2629807, 0.4035568, 
    0.5749433, 0.5985925, 0.6005945, 0.4471605, 0.06026244, -0.2896883, 
    -0.3413165, -0.1426344, 0.005233049, 0.08498579, -0.1328364, 0.1610763, 
    0.08659719, 0.01846568, -0.04486442, 0.08028185, 0.2757899, 0.09499568, 
    -0.01058705, -0.02383575, 0.2100019, 0.6945072, 0.160116, -0.4547603, 
    -0.8548906, -0.8365964, -0.6882077, -0.7726803, -0.6706945, -0.4352615, 
    -0.369164, -0.2753978, -0.02909255, 0.09128523, 0.171803, 0.3441176, 
    0.4644628, 0.4680271, 0.4046159, 0.3833747, 0.3799739, 0.2983975, 
    0.3623137, 0.3370209, 0.317945, 0.2611909, 0.1899343, 0.2157972, 
    0.2640228, 0.256129, 0.212265, 0.114413, 0.07185102, -0.02207792, 
    0.009969592, 0.009334818, 0.1660404, 0.2166428, -0.04160917, 0.009578943, 
    -0.009008259, 0.01680553, 0.01646376, -0.1051507, -0.239884, -0.07482862, 
    0.001700997, -0.008520365, 0.2026289, 0.3175379, 0.1471929, 0.00293833, 
    0.5563075, 0.777694, 0.5592698, 0.5250572, 0.4870201, 0.4303472,
  0.03659749, 0.08329296, 0.253443, 0.2392826, 0.05321503, 0.07740128, 
    0.04649301, 0.04494682, 0.2614507, 0.5779709, 1.009888, 0.0607509, 
    -0.1230219, 0.3562098, 0.4870853, 0.4477627, 0.3833747, 0.3576419, 
    0.2145112, 0.313746, 0.1078539, -0.3191152, -0.6431389, -0.7999909, 
    -0.9874911, -0.5600176, -0.2685623, -0.229744, -0.4015214, -0.195971, 
    -0.1357661, -0.02385203, -0.06719513, -0.2737219, -0.16241, -0.01698345, 
    0.1800542, 0.3520591, 0.3603599, 0.1411054, -0.3314859, -0.3733151, 
    -0.4624588, -0.577384, -0.5296459, -0.4262929, -0.2430897, -0.1714263, 
    -0.08649731, -0.05785131, 0.002271652, 0.1868744, 0.1962004, 0.2372327, 
    0.2785087, 0.3061776, 0.3213148, 0.3616138, 0.4356542, 0.4494076, 
    0.4659433, 0.4386487, 0.3919852, 0.3114676, 0.2855394, 0.2588303, 
    0.1927168, 0.1582603, 0.1575608, 0.1694585, 0.1360765, 0.03605998, 
    0.02774358, -0.1109772, -0.08955812, -0.0043208, -0.1378496, -0.05570424, 
    0.0173589, 0.0559494, 0.1093022, 0.05953002, -0.2455807, 0.1181569, 
    0.4921155, 0.5383875, 0.8374596, 0.8593348, 0.5086839, 0.2182703, 
    0.3353926, 0.3937747, 0.3860437, 0.4066654, 0.3938726, 0.2791591,
  -0.05944788, -0.02954865, 0.04198462, 0.1655034, 0.2922774, 0.1703212, 
    0.2187098, 0.4470463, 0.4123296, 0.3950121, 0.5478439, 0.2753342, 
    -0.1580318, 0.07548094, 0.5830495, 0.6523361, 0.462769, 0.3327727, 
    0.3561289, 0.2311945, -0.3550854, -0.7966375, -1.303768, -1.491999, 
    -1.395499, -0.6828041, -0.1720132, -0.1325923, -0.6088943, -1.212068, 
    -1.141154, -0.2712967, 0.1436774, 0.01509672, -0.2511634, 0.06361508, 
    0.3498135, 0.5571053, 0.4074311, 0.1602631, 0.1065845, 0.09245706, 
    0.03347301, 0.1267509, 0.2005138, 0.08550739, 0.1616464, 0.2143483, 
    0.2196708, 0.2292571, 0.2117438, 0.2640228, 0.2554617, 0.2354908, 
    0.1864185, 0.1165128, 0.02518845, -0.05265999, -0.09089279, -0.09601879, 
    -0.1350493, -0.112735, -0.08451223, -0.07894659, -0.007397056, 0.0295496, 
    0.02756399, 0.04903208, 0.07735246, 0.0208416, -0.04619908, -0.1977129, 
    -0.317081, -0.3289626, -0.2106357, 0.025383, 0.1471928, 0.08765519, 
    -0.07621205, -0.1022376, 0.1685958, 0.01519465, -0.01574564, 0.3373299, 
    0.7495704, 0.7365327, 0.803443, 0.683472, 0.4856531, 0.3373785, 0.207284, 
    -0.03197384, 0.05176687, 0.1008394, 0.0630458, -0.003506899,
  -0.1437901, 0.04940605, 0.3321052, 0.6147386, 0.5701749, 0.3468024, 
    0.5779384, 0.7027266, 0.4308355, 0.3615971, 0.4714442, 0.3824142, 
    -0.05949657, 0.2132573, 0.9658132, 0.9295502, 0.7678151, 0.6315522, 
    0.5730557, 0.1315689, -0.3883219, -0.7728262, -1.491463, -1.899959, 
    -1.927465, -1.520091, -1.437621, -0.8863356, -1.110212, -1.820027, 
    -2.206046, -1.48881, -0.2502681, -0.06799266, -0.5267, 0.04652548, 
    0.4855556, 0.4585052, 0.2901626, 0.23982, 0.08399343, -0.01751995, 
    0.07810163, 0.1767993, 0.2345796, 0.2286224, 0.3135338, 0.2744713, 
    0.189332, 0.1253672, 0.1364498, 0.1246338, 0.1910238, 0.1644135, 
    0.1566982, 0.157105, 0.03174686, 0.02069569, -0.02103567, -0.03900433, 
    -0.143024, -0.2591705, -0.2814689, -0.2571685, -0.3067131, -0.2775306, 
    -0.2093827, -0.3021398, -0.398445, -0.4845128, -0.4178624, -0.4411209, 
    -0.7059971, -0.5676185, -0.1324295, 0.08308157, -0.05025184, -0.3705316, 
    -0.3772533, -0.04714298, 0.1989508, -0.006501198, 0.1590261, 0.5413666, 
    0.6203218, 0.6233006, 0.7463636, 0.5588634, 0.4913659, 0.4093023, 
    0.3201259, 0.087672, -0.02848959, 0.1986582, -0.07105291, -0.2283931,
  0.4941168, 0.5789475, 0.7122809, 0.5076585, 0.06737518, -0.09639436, 
    0.1671962, -0.07118279, 0.1075933, 0.5187587, 0.3973883, 0.4627365, 
    -0.05715287, 0.0475018, 0.6885504, 0.7639571, 0.8116138, 0.524879, 
    0.3411713, 0.1823983, -0.1067615, -0.8763583, -1.32032, -1.495629, 
    -1.617944, -0.9771068, -0.5647526, -0.5648999, -0.7318276, -0.9332432, 
    -1.665144, -1.632088, -1.003263, -0.9162836, -0.7153716, -0.07025504, 
    0.1078706, -0.09751701, -0.1259017, -0.190567, -0.3070703, 0.01172829, 
    0.1923757, 0.1300545, 0.1319261, 0.1263113, 0.09849453, -0.04851151, 
    -0.06919765, -0.194768, -0.2032146, -0.2495537, -0.1902761, -0.135231, 
    -0.1075773, -0.03260899, -0.07915783, -0.08810997, -0.1136141, -0.116755, 
    -0.1844473, -0.2187405, -0.2405019, -0.3496652, -0.4097726, -0.4277091, 
    -0.5354245, -0.5276769, -0.3813065, -0.3688878, -0.2534907, 0.05974174, 
    -0.09440875, -0.531322, -0.9974189, -1.432283, -1.419509, -0.973155, 
    -0.2400341, 0.08745766, 0.01706505, -0.01333714, 0.2610121, 0.3761487, 
    0.4164481, 0.5040779, 0.5014091, 0.4445729, 0.5601001, 0.534986, 
    0.5756106, 0.700774, 0.9684012, 0.6557378, 0.2130132, 0.1973231,
  0.8398687, 0.820663, 0.7000901, 0.182886, -0.2049882, -0.302774, 
    -0.1480865, -0.2411046, 0.03719938, 0.1932216, 0.3573003, 0.6474696, 
    -0.03509891, -0.2260332, -0.001374811, 0.158993, 0.382431, 0.2537851, 
    0.368124, 0.4056573, -0.0134511, -1.26254, -1.489412, -1.045695, 
    -0.6673744, -0.0475657, 0.0007898808, -0.6221921, -0.7659256, -0.679695, 
    -0.6729081, -0.345711, -0.5383216, -0.8021719, -0.4942615, -0.3219147, 
    -0.5538158, -0.6379952, -0.6082258, -0.697793, -0.4826074, -0.1612377, 
    -0.1685781, -0.1560621, -0.1133699, -0.2792883, -0.3437581, -0.4348221, 
    -0.505558, -0.5467196, -0.5086994, -0.4629965, -0.3279047, -0.2259026, 
    -0.2893796, -0.2950759, -0.2322016, -0.206811, -0.1841545, -0.1994863, 
    -0.3165112, -0.3766017, -0.4124255, -0.4216218, -0.3317456, -0.2518957, 
    -0.2508866, -0.005427599, 0.07155824, 0.03802948, 0.1534266, 0.238534, 
    -0.3987544, -0.8705144, -1.10528, -1.134953, -0.8342552, -0.6341228, 
    -0.3529062, -0.2192454, -0.1097565, 0.05995369, 0.296298, 0.30901, 
    0.3979421, 0.3676195, 0.3135834, 0.3363862, 0.3290291, 0.4154878, 
    0.5226166, 0.8942957, 1.003671, 0.5606368, 0.2636316, 0.5980392,
  0.4726162, 0.3839114, 0.289852, -0.07915819, -0.2417395, -0.3426509, 
    -0.2989497, -0.1249917, 0.1456792, 0.3414314, 0.8749762, 0.614771, 
    -0.2849848, -0.3595779, -0.3290765, -0.3128169, 0.06415236, 0.1976328, 
    0.01950788, 0.0498147, -0.01498079, -1.208601, -1.346557, -0.04942191, 
    0.4557378, 0.3028407, -0.01286566, -0.316772, -0.2316156, -0.1532466, 
    0.4476163, 0.4266367, -0.3445385, -0.4748445, -0.6202707, -0.6948638, 
    -0.7781811, -0.8454177, -0.855232, -0.7648835, -0.4320869, -0.4690337, 
    -0.5276437, -0.5908594, -0.7029853, -0.907413, -1.000674, -1.018822, 
    -1.131713, -1.114737, -1.11101, -0.9991932, -0.8131089, -0.6496329, 
    -0.5929108, -0.6596103, -0.5758862, -0.5322175, -0.5070057, -0.4760323, 
    -0.446084, -0.439362, -0.414444, -0.3181062, -0.2546461, -0.08692163, 
    0.107935, 0.42343, 0.4520433, 0.08137244, 0.3066654, -0.04346478, 
    -0.8776929, -0.9912992, -0.9516344, -0.9234443, -0.8513083, -0.7646551, 
    -0.5356998, -0.4141994, -0.1622467, 0.03859949, 0.2129169, 0.2561617, 
    0.2816334, 0.1855235, 0.1558847, 0.131259, 0.09092712, 0.2515063, 
    0.2138929, 0.3368412, 0.3890873, 0.2623131, 0.2729253, 0.4794684,
  0.2638268, 0.07743382, -0.2912837, -0.8491774, -1.156534, -0.7648515, 
    -0.3899654, -0.4257239, -0.02652133, 0.4097581, 0.4094485, -0.06949002, 
    -0.4190831, -0.02743274, 0.04283094, -0.1619379, -0.07839322, 0.05168533, 
    0.0524025, 0.1045499, -0.4199452, -1.375024, -0.8968501, 0.2084233, 
    0.4023848, 0.1156825, 0.06127155, -0.06520891, 0.0007736236, 0.1118249, 
    0.4093833, 0.08695507, -0.06359828, 0.2076094, -0.1876867, -0.4549878, 
    -0.7563714, -0.9439688, -0.9016838, -0.7155836, -0.5239656, -0.7649648, 
    -0.7683663, -0.9828527, -1.15935, -1.271655, -1.505492, -1.645222, 
    -1.827351, -1.777058, -1.694782, -1.650625, -1.666966, -1.51529, 
    -1.26472, -1.188027, -0.9482489, -0.7835021, -0.6517158, -0.5340075, 
    -0.4199452, -0.3254626, -0.2428131, -0.1664791, -0.01568146, 0.2679291, 
    0.1008718, 0.2373953, 0.2488042, -0.06223094, -0.06159616, -0.4612374, 
    -0.9068589, -0.6065502, -0.8251209, -1.017064, -0.9302812, -0.6991768, 
    -0.3933177, -0.4163809, -0.2184803, 0.001360416, 0.1725674, 0.2738214, 
    0.2435646, 0.1147065, -0.06533909, -0.233243, -0.3534083, -0.3507071, 
    -0.2311921, 0.100286, 0.2415773, 0.3494878, 0.3460535, 0.267424,
  -0.5717036, -0.9078365, -1.183666, -1.31591, -1.232576, -0.5535394, 
    -0.3902095, -0.7743403, -0.2862869, 0.2366622, -0.2776121, -0.6030511, 
    -0.235701, 0.2209232, 0.1424565, -0.1978269, -0.1351801, 0.1016198, 
    -0.02144289, -0.4037348, -0.760115, -0.5688553, -0.04100728, 0.2111418, 
    0.1487228, 0.008586228, -0.1720129, 0.1143154, 0.3938565, 0.3580488, 
    0.4466882, 0.2498622, 0.1361741, 0.3178631, 0.0981369, -0.1648514, 
    -0.5258866, -0.6641189, -0.7578363, -0.8345942, -0.7782466, -0.8939366, 
    -0.9659581, -1.241495, -1.422859, -1.56005, -1.766593, -1.871687, 
    -2.048835, -2.127172, -2.188207, -2.198787, -2.111059, -1.862931, 
    -1.62989, -1.477546, -1.1857, -1.045971, -0.8905997, -0.6528556, 
    -0.4423087, -0.2936113, -0.1592037, 0.04426324, 0.3173919, 0.2545829, 
    -0.07746482, -0.1041907, -0.05051218, -0.1986403, -0.05578518, 
    -0.4522047, -0.6708732, -0.2961991, -0.4011469, -0.4638098, -0.5522213, 
    -0.477791, -0.3852452, -0.3857499, -0.1767169, -0.08319473, -0.04245567, 
    -0.03503382, -0.1612055, -0.2903879, -0.4370351, -0.5935454, -0.6966383, 
    -0.7415276, -0.6650138, -0.445173, -0.1528723, 0.2135341, 0.2239017, 
    -0.2328852,
  -0.8863683, -1.191495, -1.485847, -1.596704, -1.163435, -0.5582597, 
    -0.4935626, -0.4395584, 0.01903534, 0.1723392, -0.183341, -0.1749914, 
    0.2686771, 0.1290126, -0.3484941, -0.5046788, -0.198966, 0.04340041, 
    -0.1373122, -0.2665767, 0.1878017, 0.8059175, 0.4836354, -0.006045341, 
    0.1855559, -0.0927639, -0.1929426, 0.3741297, 0.4921962, 0.1937425, 
    0.08656454, 0.02912658, 0.007039964, 0.1727952, 0.1793055, 0.02313691, 
    -0.2013098, -0.2647051, -0.4401281, -0.7865477, -1.022974, -1.265177, 
    -1.445434, -1.533732, -1.519848, -1.624275, -1.78396, -1.930558, 
    -2.07281, -2.054467, -2.120955, -2.131486, -2.009464, -1.834041, 
    -1.596948, -1.321655, -1.155004, -1.094018, -0.9730382, -0.8349848, 
    -0.6021234, -0.3445389, -0.06485164, 0.3956635, 0.3848886, 0.06748962, 
    0.0661056, 0.2556726, 0.1604904, -0.1281488, -0.09362721, -0.2696041, 
    -0.3617263, -0.2154699, -0.1934972, -0.03622183, 0.1650476, 0.188306, 
    0.02948451, -0.06223083, 0.009204626, -0.1104244, -0.2207923, -0.3191158, 
    -0.5007889, -0.6403397, -0.7675695, -0.9152257, -1.010603, -1.048152, 
    -1.109187, -1.015193, -0.7191159, -0.4473709, -0.2891515, -0.566007,
  -1.433374, -1.580379, -1.601033, -1.528182, -0.9532301, -0.3612707, 
    0.1096115, 0.3539802, 0.2038336, 0.08010364, 0.1532152, 0.2255783, 
    0.2125409, -0.2279211, -0.497143, -0.4278234, -0.3444575, -0.1517492, 
    0.09274954, 0.2662032, 0.419394, 0.3180916, 0.04252172, 0.293401, 
    0.5515881, 0.2880132, 0.5712816, 0.708049, 0.2272711, -0.1365473, 
    -0.2225173, -0.2114171, -0.0748449, 0.03316294, 0.1420171, 0.1034429, 
    0.01838422, -0.08172977, -0.1336503, -0.3224516, -0.5587149, -0.6458404, 
    -0.6674874, -0.7980864, -0.9630115, -1.15336, -1.287572, -1.451308, 
    -1.572956, -1.535553, -1.599078, -1.603343, -1.461123, -1.3142, 
    -1.104516, -0.9354403, -0.876554, -0.7207757, -0.542244, -0.5048907, 
    -0.3981525, -0.201082, 0.06856346, 0.3071382, 0.3605723, 0.2518803, 
    0.3852462, 0.4498949, 0.03000546, -0.2841873, -0.2496495, -0.2823644, 
    -0.3037186, -0.2450763, -0.2418211, 0.04961789, 0.3858817, 0.4352951, 
    0.1335702, 0.006063938, 0.07316971, 0.06524372, -0.04017615, -0.3046947, 
    -0.588419, -0.7503817, -0.7938389, -0.8681068, -0.9772049, -1.08129, 
    -1.233048, -1.252042, -1.242309, -1.13046, -0.784155, -0.9207923,
  -2.098168, -1.994132, -1.189688, -0.5481193, -0.1424553, 0.03243113, 
    0.1335372, 0.06784713, -0.0945065, 0.02059782, 0.02639198, -0.08605909, 
    -0.1996006, -0.3002518, -0.1841222, -0.05329531, -0.2744704, -0.2445878, 
    0.06372935, 0.1177331, -0.05987096, -0.1048416, 0.2913824, 0.3587325, 
    0.1054286, 0.03970599, 0.6256759, 0.4735437, 0.04865772, -0.0707922, 
    -0.1778072, -0.2906003, -0.2399977, -0.1629798, -0.01755333, -0.02515435, 
    -0.09206462, -0.131762, -0.1744375, 0.0844655, 0.2407317, 0.2999601, 
    0.3252048, 0.2695079, 0.1655045, -0.01441145, -0.1635652, -0.2796297, 
    -0.377172, -0.4437408, -0.5430412, -0.5602288, -0.4335847, -0.3707428, 
    -0.3296456, -0.2603259, -0.1565828, -0.04448938, 0.0429616, 0.1164317, 
    0.220696, 0.2333751, 0.2184658, 0.228166, 0.1426029, 0.1156174, 
    0.1322027, 0.102043, -0.127677, -0.3119054, -0.1630122, 0.01561737, 
    0.1353438, 0.1852298, 0.1375897, 0.09751844, 0.1746993, 0.2783296, 
    0.4471283, 0.4212332, 0.2950935, 0.2620373, 0.1654391, -0.1105051, 
    -0.3465562, -0.4693754, -0.5307035, -0.6518135, -0.7857001, -0.7819242, 
    -0.8098869, -0.9391026, -0.9608634, -0.7231195, -0.58199, -1.256062,
  -0.8001869, -0.3809973, 0.03780222, 0.1654707, 0.113534, 0.2475674, 
    0.3957117, 0.2365647, 0.1238204, 0.2445398, 0.1313237, 0.03225148, 
    0.136581, 0.2323166, 0.477092, 0.4489017, 0.1621341, 0.2334396, 
    0.3619878, 0.153329, 0.05577037, 0.2656336, 0.4559656, 0.372844, 
    0.1500413, 0.2275966, 0.5302334, 0.3429284, 0.05651909, 0.09314013, 
    0.06385934, 0.02251816, 0.1236906, 0.2332611, 0.1863532, 0.08799696, 
    -0.03654647, 0.04291272, 0.293905, 0.5533614, 0.8428478, 0.890341, 
    0.8994558, 0.9459891, 0.9994559, 1.019818, 1.04192, 1.049489, 1.017067, 
    0.9269791, 0.8177991, 0.7166429, 0.6446867, 0.5674901, 0.5323176, 
    0.5919042, 0.6958914, 0.7548919, 0.8627858, 0.9800384, 0.886663, 
    0.5961518, 0.2204514, 0.04125202, -0.003539562, -0.033162, -0.05046332, 
    0.0403893, 0.1524987, 0.1454513, 0.2855393, 0.4811448, 0.5412847, 
    0.5386804, 0.4659917, 0.3871348, 0.144556, 0.08119345, 0.2453704, 
    0.2982514, 0.2488046, 0.3483002, 0.364804, 0.2677827, 0.206243, 
    0.1968026, 0.09390545, -0.1280012, -0.2625551, -0.1960683, -0.2684803, 
    -0.4868069, -0.5807199, -0.578409, -0.7163486, -0.8419182,
  -0.003262997, 0.2049727, 0.4674568, 0.5103439, 0.5434819, 0.6797938, 
    0.8236578, 0.6490647, 0.4177821, 0.5204514, 0.7811285, 1.033944, 1.29423, 
    1.333863, 1.261141, 0.886809, 0.6445072, 0.7043052, 0.7362226, 0.5200605, 
    0.4203374, 0.380982, 0.2269292, 0.05821179, -0.01662546, -0.006290317, 
    0.04235876, 0.0857178, 0.08804572, 0.02012563, -0.03918421, -0.03448009, 
    0.12483, 0.2735443, 0.2543056, 0.1294357, 0.2296799, 0.5897386, 0.929859, 
    1.190308, 1.561923, 1.769752, 1.960263, 2.020321, 1.925611, 1.898951, 
    1.999716, 2.026214, 1.915554, 1.802076, 1.708668, 1.621251, 1.600791, 
    1.596982, 1.595127, 1.624098, 1.647225, 1.644443, 1.539902, 1.320761, 
    0.9459727, 0.4911714, 0.2051518, 0.187541, 0.1958096, 0.3801192, 
    0.5931886, 0.707642, 0.6819912, 0.5382898, 0.4339768, 0.3323329, 
    0.1284918, -0.002628028, 0.08729684, 0.1274173, 0.01358271, -0.08322716, 
    -0.09768057, 0.01029468, 0.04906452, 0.09685111, 0.117815, 0.1313078, 
    0.1820896, 0.2359142, 0.2214284, 0.1250906, 0.08119392, 0.1185312, 
    0.1667409, 0.1540456, 0.1026621, -0.02336311, -0.1216218, -0.1230867,
  0.5785568, 0.7464931, 1.120044, 1.17688, 0.9912847, 0.9064539, 1.053785, 
    1.040813, 0.9757246, 1.082788, 1.338143, 1.465585, 1.345353, 1.052206, 
    0.8048912, 0.6079022, 0.5612877, 0.6432863, 0.6838464, 0.5590256, 
    0.3646083, 0.1487391, 0.001929283, -0.02240348, 0.03278875, 0.07691264, 
    0.160702, 0.2549572, 0.214771, 0.01530802, -0.09027433, 0.03750896, 
    0.1841067, 0.2589279, 0.2162684, 0.2109949, 0.3183029, 0.5082768, 
    0.9048752, 1.457138, 1.689706, 1.785816, 2.0469, 2.298462, 2.323381, 
    2.148609, 1.938453, 1.776555, 1.742392, 1.863192, 1.992554, 2.047437, 
    2.082691, 2.084254, 2.09721, 2.092685, 2.011793, 1.743157, 1.349146, 
    0.951653, 0.5561609, 0.2162846, 0.1427333, 0.2311772, 0.4511155, 
    0.5205652, 0.6209558, 0.5691817, 0.3781821, 0.1841882, 0.01766825, 
    -0.1325597, -0.2315993, -0.2292719, -0.1790439, -0.1665764, -0.1988523, 
    -0.1355059, -0.01825297, 0.06931204, -0.004450977, 0.1264898, 
    -0.08654726, -0.1280026, -0.08636856, -0.08975363, -0.1704338, 
    -0.2716703, -0.2403066, 0.01097918, 0.3794038, 0.5846281, 0.6314869, 
    0.6204189, 0.6335053, 0.5927333,
  1.213567, 1.171949, 1.211565, 0.9472743, 0.8270269, 0.9886807, 1.201831, 
    1.12426, 0.9830817, 0.9391526, 0.9357669, 0.8829677, 0.6815355, 
    0.4221767, 0.3085698, 0.2207769, 0.1918706, 0.1597254, 0.1312588, 
    0.05344272, -0.0890379, -0.1886473, -0.1394773, 0.03669453, 0.1751227, 
    0.1226645, 0.01818895, 0.07432508, 0.1041588, 0.08758986, 0.2092862, 
    0.3595461, 0.3703211, 0.2155522, 0.178101, 0.3151454, 0.4307541, 
    0.4937098, 0.6325445, 0.85577, 0.8224692, 0.7333746, 0.7504644, 
    0.8107343, 0.8436445, 0.802222, 0.8327724, 0.9738693, 1.181552, 1.426294, 
    1.608603, 1.746819, 1.845012, 1.910214, 1.931308, 1.917457, 1.712736, 
    1.342522, 0.9263107, 0.6686773, 0.41329, 0.2564866, 0.1567632, 0.3611253, 
    0.4668708, 0.4222254, 0.2831303, 0.04178894, -0.1233149, -0.1473384, 
    -0.1317947, -0.2512121, -0.4255936, -0.4566646, -0.3641841, -0.2180741, 
    -0.05230236, 0.04893446, 0.1269944, 0.130982, 0.08765513, 0.005949393, 
    -0.09872182, -0.06439567, 0.04969937, 0.04514182, -0.04732239, 
    -0.04348111, 0.2270756, 0.6273034, 0.9605883, 1.100936, 1.127336, 
    1.053915, 1.043043, 1.085197,
  0.9587653, 0.8736416, 0.688648, 0.613827, 0.816724, 0.9551192, 0.9469, 
    0.7817632, 0.4807215, 0.3212489, 0.2048915, 0.1075119, 0.03405813, 
    -0.05181426, -0.1831294, -0.2578037, -0.2821368, -0.2094318, -0.1751704, 
    -0.2489009, -0.3630123, -0.4050045, -0.3406487, -0.2646725, -0.2320225, 
    -0.2038488, -0.1945879, -0.1487545, -0.08713341, 0.1062748, 0.2518964, 
    0.4649665, 0.4734461, 0.3245691, 0.2863043, 0.3751063, 0.4822026, 
    0.4120038, 0.1087976, 0.1052175, 0.06822205, 0.04126835, 0.004370451, 
    -0.0700922, -0.1273835, -0.1453521, -0.08644915, 0.08077073, 0.3742599, 
    0.6358972, 0.8219485, 0.9805912, 1.082365, 1.120061, 1.281454, 1.048691, 
    0.934335, 0.774667, 0.6056893, 0.4304612, 0.124227, 0.02821505, 
    0.1591884, 0.3177984, 0.4256759, 0.3569098, 0.2146246, 0.1459234, 
    0.1037684, 0.08941296, 0.03394419, -0.07884878, -0.1729894, -0.08801219, 
    0.03454643, 0.2037848, 0.4314865, 0.5429124, 0.4545009, 0.2753505, 
    0.1823003, 0.2501226, 0.4583582, 0.7389573, 0.9130293, 0.7431566, 
    0.4458745, 0.4128993, 0.6114345, 0.8028896, 0.9766363, 1.178378, 
    1.377971, 1.406552, 1.220517, 1.136711,
  0.7133061, 0.5323979, 0.2825282, 0.3346766, 0.3708908, 0.4489019, 
    0.3641688, 0.2028732, 0.09172414, -0.03833771, -0.1630447, -0.2393468, 
    -0.2439041, -0.2031326, -0.2336177, -0.2864332, -0.2266192, -0.1042072, 
    -0.09203255, -0.1556718, -0.2352779, -0.2987708, -0.2555742, -0.1786376, 
    -0.136043, -0.07687932, -0.01594192, 0.04642785, 0.1470627, 0.3217695, 
    0.5017177, 0.5524011, 0.3941655, 0.1568609, 0.124797, 0.2851486, 
    0.4222419, 0.2875901, 0.2286054, 0.1169518, 0.04379129, -0.1431556, 
    -0.2556715, -0.2724361, -0.3487053, -0.4191639, -0.4919343, -0.9457099, 
    -0.7814524, -0.5767159, -0.3557854, -0.2227128, 0.09720922, 0.0645268, 
    -0.04434371, -0.1639237, -0.1551021, -0.06706512, -0.02919066, 
    -0.0381586, 0.04982961, 0.1751063, 0.3480068, 0.4647385, 0.4541265, 
    0.3684983, 0.3639735, 0.3913824, 0.3943934, 0.3576423, 0.2389246, 
    0.09712778, 0.08693899, 0.1617925, 0.2852788, 0.4599208, 0.7401779, 
    0.766008, 0.524618, 0.3679774, 0.311467, 0.3793381, 0.5774499, 0.7128174, 
    0.7816654, 0.7167895, 0.6324308, 0.6500248, 0.8054609, 0.8997155, 
    0.9841067, 1.083326, 1.215796, 1.226864, 1.07159, 0.8763267,
  0.4811123, 0.4080002, 0.3751877, 0.2984136, 0.2961675, 0.205982, 
    0.08693898, -0.1794835, -0.3312088, -0.4516515, -0.5070063, -0.4651606, 
    -0.3524653, -0.233634, -0.1135005, -0.0584386, -0.06610489, -0.06390762, 
    -0.1247963, -0.2006589, -0.2107502, -0.1775146, -0.1607664, -0.1437576, 
    -0.1003169, -0.06926221, 0.008293152, 0.08682506, 0.1179774, 0.1599045, 
    0.1441818, -0.003262838, -0.1908768, -0.2687413, -0.1961828, -0.02193141, 
    0.06319231, 0.08796442, 0.01866108, -0.01869243, -0.08389425, -0.1943762, 
    -0.2890863, -0.364347, -0.3877192, -0.3610265, -0.3495681, -0.323103, 
    -0.2416899, -0.1470778, -0.1440504, -0.05803192, -0.2571853, -0.2236243, 
    -0.1941484, -0.1585364, -0.09518999, -0.0755772, 0.04105687, 0.1736579, 
    0.2901292, 0.3999112, 0.4719648, 0.4443606, 0.3561773, 0.3132083, 
    0.3014733, 0.3223716, 0.323674, 0.2403895, 0.1554123, 0.09737193, 
    0.1115321, 0.2335861, 0.3562098, 0.5759038, 0.7186447, 0.7537358, 
    0.4764572, 0.3027267, 0.22037, 0.2811937, 0.4558517, 0.3317795, 
    0.08422136, -0.07215929, -0.03714967, 0.2304289, 0.5036225, 0.6515553, 
    0.6345468, 0.6105391, 0.5621502, 0.59397, 0.6133059, 0.5885988,
  0.1027918, 0.0498457, 0.02956599, 0.05324763, 0.03137258, -0.1085037, 
    -0.2456131, -0.3863846, -0.4529862, -0.4079015, -0.3194738, -0.1823481, 
    -0.02224071, 0.1065028, 0.2059006, 0.2936284, 0.3258387, 0.2839278, 
    0.1811447, 0.08125871, 0.03036338, 0.02227426, 0.03718313, 0.0683029, 
    0.1271083, 0.1999435, 0.2633224, 0.2459071, 0.1567958, 0.02435756, 
    -0.08314574, -0.1310298, -0.1357987, -0.03845173, 0.03842008, 0.1152918, 
    0.2533941, 0.1937587, 0.2761968, 0.2823492, 0.2928146, 0.2360764, 
    0.139771, 0.04825068, -0.03073692, -0.08804488, -0.04385543, 0.03742707, 
    0.1378342, 0.2252036, 0.259302, 0.2927818, 0.3181076, 0.2233815, 
    0.2704682, 0.317538, 0.3300707, 0.3101809, 0.2186121, 0.3844161, 
    0.3146734, 0.2316496, 0.1169357, 0.03020048, -0.01854622, 0.05469596, 
    0.100269, 0.06537318, -0.03978634, -0.04095814, -0.04304149, 0.05632376, 
    0.249439, 0.3858973, 0.5224533, 0.4526779, 0.3436285, 0.1561935, 
    0.04580942, -0.00752716, 0.04738823, 0.1384364, 0.04025912, -0.1922929, 
    -0.5194414, -0.6510493, -0.5247473, -0.2943598, -0.03944439, 0.1771083, 
    0.3227297, 0.341496, 0.229289, 0.1644289, 0.18313, 0.1767174,
  -0.4457923, -0.4104568, -0.3350338, -0.259936, -0.1792558, -0.1159909, 
    -0.03625441, 0.02458537, 0.1142502, 0.203557, 0.2824631, 0.3524338, 
    0.4230881, 0.422079, 0.4417892, 0.4781336, 0.3191493, 0.2541916, 
    0.2061936, 0.2019129, 0.233342, 0.2861089, 0.3633878, 0.448218, 
    0.4914471, 0.4909102, 0.42286, 0.3465093, 0.2723394, 0.2525966, 
    0.2111415, 0.2225995, 0.2470138, 0.2683842, 0.3294194, 0.3472905, 
    0.3384361, 0.3164799, 0.2684491, 0.2382898, 0.2589442, 0.2247318, 
    0.1922612, 0.1819909, 0.2231531, 0.3132247, 0.4188234, 0.476343, 
    0.530705, 0.541317, 0.5253015, 0.5127201, 0.4865649, 0.4840908, 
    0.5017996, 0.5029385, 0.452255, 0.3643312, 0.2844164, 0.2398036, 
    0.2046797, 0.1573329, 0.08212113, -0.162231, -0.1246496, -0.1785722, 
    -0.2046302, -0.2307693, -0.2493566, -0.2024328, -0.1646886, -0.03081818, 
    0.08794811, 0.2028407, 0.1634038, 0.06753795, -0.03352, -0.05568799, 
    0.02163959, 0.1146245, 0.2153732, 0.09883666, 0.003426433, -0.2301672, 
    -0.4409419, -0.5204828, -0.4670001, -0.2517169, -0.009073317, 0.1529058, 
    0.189006, 0.1178472, -0.01848093, -0.1434971, -0.3854893, -0.4671625,
  -0.3817295, -0.2304602, -0.05586696, 0.0745362, 0.1600832, 0.1588626, 
    0.1270269, 0.2223233, 0.2485278, 0.322258, 0.3372645, 0.3276779, 
    0.3380132, 0.3450933, 0.3260503, 0.2756923, 0.2204513, 0.1682867, 
    0.1309983, 0.1237392, 0.1446539, 0.1737388, 0.229354, 0.2817469, 
    0.3094649, 0.1935794, 0.1379805, 0.1366134, 0.09055209, 0.06345248, 
    0.09058499, 0.1252689, 0.1334395, 0.1247156, 0.1342373, 0.1476488, 
    0.1450117, 0.1604251, 0.153638, 0.1539311, 0.1469649, 0.1592858, 
    0.2127851, 0.2885176, 0.3863039, 0.485604, 0.5282636, 0.531356, 
    0.4986086, 0.4447838, 0.3628503, 0.2557214, 0.1558191, 0.08882689, 
    0.04745317, 0.004305363, -0.03474081, -0.06765079, -0.09942162, 
    -0.1406976, -0.1762445, -0.1951739, -0.202563, -0.192716, -0.1173742, 
    -0.1848709, -0.1423579, -0.09056752, -0.03767039, 0.02458547, 0.0766037, 
    0.1450933, 0.1592534, 0.133993, 0.09071502, 0.05080616, 0.09982967, 
    0.1243086, 0.06024611, 0.1012293, 0.1485111, 0.1035242, 0.008276939, 
    -0.1304764, -0.273266, -0.3756752, -0.4020748, -0.3539791, -0.2537026, 
    -0.192781, -0.1701248, -0.2942297, -0.3509516, -0.4249425, -0.423673, 
    -0.4225173,
  -0.07881622, -0.02032013, 0.0274826, 0.0640223, 0.03749236, 0.06687063, 
    0.1143478, 0.1082606, 0.1543381, 0.1882085, 0.2325607, 0.269605, 
    0.3147059, 0.3380295, 0.3349859, 0.2970464, 0.230803, 0.1478439, 
    0.05892783, -0.02237093, -0.06844831, -0.1043698, -0.1245846, -0.1018145, 
    -0.08700323, -0.2575109, -0.2390051, -0.1109452, -0.07491004, 
    -0.04445767, 0.0119226, 0.0547775, 0.09141481, 0.1239343, 0.1414636, 
    0.1549239, 0.1547936, 0.1542563, 0.1540774, 0.1513107, 0.1519291, 
    0.1447189, 0.1571051, 0.1596441, 0.1656662, 0.1738856, 0.1610113, 
    0.1472744, 0.1201584, 0.08990127, 0.06771702, 0.04107305, 0.006226093, 
    -0.01880646, -0.04452261, -0.08358511, -0.1098384, -0.1366287, -0.167423, 
    -0.1999425, -0.2467362, -0.2714269, -0.2783117, -0.2685623, -0.251977, 
    -0.219604, -0.1631912, -0.1022863, -0.02969513, 0.04128469, 0.09510954, 
    0.1182378, 0.1189052, 0.07762909, 0.04595596, 0.02985901, 0.02054912, 
    0.008618712, -0.005264699, -0.02360788, -0.06071727, -0.1308019, 
    -0.2114658, -0.2883379, -0.3509681, -0.3780025, -0.3856685, -0.376619, 
    -0.3521401, -0.3132889, -0.2638585, -0.21477, -0.2114171, -0.1806391, 
    -0.1545486, -0.1222733,
  -0.03060659, -0.001521301, 0.02707571, 0.06512909, 0.1132736, 0.1552007, 
    0.1924728, 0.2159103, 0.2373947, 0.2564377, 0.2763433, 0.2807866, 
    0.2825282, 0.2795985, 0.2619227, 0.2355555, 0.1935468, 0.1434331, 
    0.1039637, 0.06947482, 0.04628158, 0.01301336, -0.002334952, 
    0.0009850264, 0.01403844, 0.03301632, 0.05100131, 0.07486212, 0.1088626, 
    0.1447513, 0.1780847, 0.2020267, 0.2194259, 0.248641, 0.2656009, 
    0.276636, 0.27994, 0.2912196, 0.2977626, 0.295891, 0.2949468, 0.2885666, 
    0.2837326, 0.2840581, 0.2762457, 0.2505132, 0.2234624, 0.1999761, 
    0.1706304, 0.1323003, 0.1017339, 0.07162323, 0.02878469, -0.02393341, 
    -0.06888784, -0.1202062, -0.1738358, -0.2081456, -0.2397049, -0.2740962, 
    -0.2979569, -0.299324, -0.2965083, -0.2753494, -0.2408442, -0.2081131, 
    -0.1676997, -0.1336176, -0.09183708, -0.05674589, -0.01835066, 
    0.01342016, 0.03142142, 0.03132385, 0.02792209, 0.02430886, 
    -0.0006260872, -0.0358963, -0.05869901, -0.10852, -0.1328527, -0.1718175, 
    -0.1660395, -0.1992589, -0.1941483, -0.2300857, -0.2032954, -0.2120193, 
    -0.2021398, -0.1809972, -0.1715571, -0.1499914, -0.1279048, -0.110229, 
    -0.09685007, -0.06686961,
  0.04899952, 0.06804249, 0.08697155, 0.1116787, 0.1282313, 0.1361253, 
    0.1487718, 0.1601161, 0.1804937, 0.1864833, 0.1829026, 0.1841558, 
    0.1852138, 0.1793868, 0.1712977, 0.1573003, 0.1395919, 0.1302658, 
    0.1168705, 0.1066655, 0.09691614, 0.08467656, 0.07486212, 0.07030481, 
    0.06343627, 0.06825405, 0.06597537, 0.07113492, 0.07020718, 0.06766808, 
    0.06722867, 0.0700444, 0.07198137, 0.08404195, 0.09178931, 0.1018966, 
    0.1210698, 0.1276779, 0.1317958, 0.1369227, 0.140536, 0.1368576, 
    0.1384526, 0.1282801, 0.1117111, 0.1030034, 0.08407441, 0.06146699, 
    0.03749239, 0.01485237, -0.01211703, -0.03680772, -0.06144971, 
    -0.09182078, -0.1020747, -0.1214758, -0.1441483, -0.1586828, -0.1705317, 
    -0.1837804, -0.1956782, -0.1994217, -0.1940994, -0.1927648, -0.184464, 
    -0.1711014, -0.1590408, -0.1546137, -0.1432856, -0.1305578, -0.1163488, 
    -0.1059484, -0.09157665, -0.0764562, -0.05829214, -0.05161895, 
    -0.04491322, -0.03693797, -0.03049266, -0.02852326, -0.0358963, 
    -0.03972117, -0.03838654, -0.03648224, -0.03959096, -0.0436437, 
    -0.04558054, -0.04431102, -0.04304148, -0.03955841, -0.02774201, 
    -0.01548614, -0.01338653, -0.004923001, 0.01197153, 0.02741751,
  0.4246776, 0.3838084, 0.3367219, 0.2848668, 0.2298375, 0.1725127, 
    0.1146516, 0.05677408, 0.0005729049, -0.05297518, -0.1021779, -0.1478647, 
    -0.1899056, -0.2297652, -0.2679334, -0.3047822, -0.3413055, -0.3782685, 
    -0.4157031, -0.4529104, -0.4905405, -0.5271125, -0.5617318, -0.592917, 
    -0.619854, -0.6404433, -0.6543913, -0.6607881, -0.6593723, -0.6491508, 
    -0.6287079, -0.5984344, -0.5589812, -0.5116832, -0.4570117, -0.3970177, 
    -0.3330045, -0.2664841, -0.198988, -0.1325813, -0.06807944, -0.006946623, 
    0.05013335, 0.103242, 0.1522822, 0.1983266, 0.2336295, 0.2801299, 
    0.3101757, 0.3183298, 0.3456082, 0.3395052, 0.3650422, 0.4425974, 
    0.4573765, 0.4839706, 0.5403337, 0.5638852, 0.5480647, 0.5753431, 
    0.6221371, 0.6358738, 0.6637058, 0.6647482, 0.669517, 0.6745148, 
    0.6736522, 0.6749377, 0.6641955, 0.648994, 0.628633, 0.6125193, 
    0.6002798, 0.3357778, 0.4393263, 0.4655304, 0.3889189, 0.2320018, 
    0.4236183, 0.3927584, 0.379169, 0.3747749, 0.3808126, 0.3855653, 
    0.3936868, 0.4102397, 0.4311543, 0.4529967, 0.4738951, 0.4923043, 
    0.5054874, 0.513413, 0.5128107, 0.5030956, 0.4840527, 0.4580107,
  0.4816926, 0.4981965, 0.4924675, 0.4716829, 0.4374056, 0.394567, 0.3484082, 
    0.3041862, 0.2634961, 0.2238151, 0.184834, 0.1481967, 0.1155469, 
    0.08743817, 0.06541657, 0.04930317, 0.0365591, 0.02716792, 0.01336598, 
    -0.004960775, -0.0341115, -0.07475281, -0.1300914, -0.1998014, 
    -0.2825813, -0.374053, -0.4653292, -0.5481267, -0.6147447, -0.6606269, 
    -0.6837378, -0.6798964, -0.6503558, -0.5968242, -0.5238099, -0.4375138, 
    -0.3429184, -0.2457666, -0.1513801, -0.0636363, 0.01839495, 0.05845022, 
    0.0551953, 0.1064973, 0.1131544, 0.06759763, 0.1221874, 0.1288443, 
    0.110729, 0.06645823, 0.0585804, 0.06779289, 0.04871726, 0.1040397, 
    0.1752145, 0.05540609, 0.0451684, 0.01273012, 0.01674938, 0.007994175, 
    0.05148363, 0.1129417, 0.1625681, 0.1769238, 0.2306671, 0.3233271, 
    0.3745962, 0.4151887, 0.474515, 0.5218783, 0.5620638, 0.5732456, 
    0.5675815, 0.5248082, 0.4879426, 0.3992546, 0.3436719, 0.2358919, 
    0.08405268, 0.1389682, -0.00525403, -0.1657197, -0.05020857, -0.1880176, 
    -0.1716275, -0.1796193, -0.1118302, -0.06746149, -0.00997448, 0.06068039, 
    0.1381869, 0.2152371, 0.2795928, 0.3467481, 0.4101596, 0.4547886,
  0.196455, 0.2515332, 0.2868197, 0.3112989, 0.316198, 0.3048373, 0.2885124, 
    0.2701856, 0.2437207, 0.2225618, 0.2059277, 0.1926466, 0.1691273, 
    0.1325555, 0.07510066, -0.01580095, -0.1343393, -0.2621717, -0.3680801, 
    -0.4354467, -0.4689589, -0.4518685, -0.372848, -0.3056607, -0.268112, 
    -0.2550424, -0.257093, -0.2879524, -0.3412075, -0.3985152, -0.4393525, 
    -0.4518523, -0.4443007, -0.414175, -0.3594871, -0.3081512, -0.2496061, 
    -0.188179, -0.1217899, -0.05103874, 0.01670265, 0.1050477, 0.1647811, 
    0.22082, 0.1591669, 0.1790069, 0.1316928, 0.09328124, 0.05625325, 
    0.01230793, -0.03132813, -0.06791668, -0.09503257, -0.1090788, 
    -0.1172168, -0.1284475, -0.1505991, -0.2077768, -0.2526494, -0.3076625, 
    -0.358574, -0.3812956, -0.3497363, -0.2772105, -0.206735, -0.1495247, 
    -0.1059863, -0.06526363, -0.01711929, 0.02759099, 0.06902981, 0.1098014, 
    0.1617708, 0.1988313, 0.2464063, 0.2833856, 0.347692, 0.2731152, 
    0.2868848, 0.2626496, 0.2205108, 0.1337106, 0.1227245, 0.05433273, 
    0.04466486, -0.06313157, -0.1059053, -0.0901823, -0.09797859, -0.1667452, 
    -0.08375406, -0.05880213, 0.00041008, 0.04800129, 0.09249997, 0.1409211,
  0.02863264, 0.1372914, 0.2612822, 0.3345573, 0.3588738, 0.3547562, 
    0.3641311, 0.4147816, 0.5017446, 0.5814322, 0.6252799, 0.6406934, 
    0.63778, 0.6243196, 0.5809602, 0.4725456, 0.3220084, 0.1603062, 
    -0.0372529, -0.3120255, -0.4785795, -0.5666327, -0.5450492, -0.4268684, 
    -0.2847136, -0.2335091, -0.2568166, -0.2918591, -0.3028617, -0.2950003, 
    -0.3004363, -0.3302702, -0.3783823, -0.4246062, -0.4432907, -0.4245574, 
    -0.4050589, -0.3769517, -0.3681288, -0.3865528, -0.3896618, -0.3290987, 
    -0.1990042, -0.03867054, 0.08642912, 0.2323272, 0.05039382, 0.01186812, 
    -0.08318365, -0.1531544, -0.2316537, -0.2884407, -0.2900358, -0.2539681, 
    -0.2177864, -0.1445605, -0.06923509, -0.1186817, -0.1485159, -0.1676562, 
    -0.2490203, -0.3520637, -0.4233365, -0.4127245, -0.3637829, -0.292347, 
    -0.2478323, -0.2159476, -0.1911106, -0.1528127, -0.09884119, -0.05881858, 
    -0.03985667, -0.03453469, 0.00249362, 0.0151726, 0.06634426, 0.132783, 
    0.2031282, 0.2774446, 0.3252962, 0.3932812, 0.3973014, 0.363024, 
    0.2971222, 0.2359733, 0.1673697, 0.06046891, -0.0390594, -0.0983367, 
    -0.01099968, 0.02181244, -0.0487113, -0.07947493, -0.08023834, -0.06101608,
  -0.1303692, -0.07700014, -0.04041147, -0.03505659, -0.004571438, 
    -0.01948071, -0.05382204, -0.08043289, -0.1603656, -0.07940865, 
    -0.02957153, 0.05133724, 0.1993995, 0.2517285, 0.2893261, 0.5678255, 
    0.7179556, 0.6494982, 0.4777376, 0.2682161, 0.3110375, 0.2210636, 
    0.0577507, -0.03842545, -0.08292532, -0.03048229, 0.01860666, 0.01803684, 
    0.0150094, 0.02594709, 0.03398752, 0.04975891, 0.03115582, -0.04818988, 
    -0.1525685, -0.264694, -0.3507617, -0.4052213, -0.4571257, -0.5426238, 
    -0.622051, -0.680824, -0.6031218, -0.392868, -0.2001758, 0.0067904, 
    0.03390622, 0.0821321, 0.03699863, -0.03316772, -0.09773469, -0.1769828, 
    -0.2528615, -0.2885223, -0.2687957, -0.2040984, -0.1732064, -0.1990691, 
    -0.235446, -0.2992969, -0.3411915, -0.4043423, -0.4648077, -0.4868621, 
    -0.4892058, -0.4385065, -0.3221161, -0.1722951, 0.01603484, 0.1916862, 
    0.2373405, 0.3220739, 0.4399123, 0.4624711, 0.540319, 0.5974153, 
    0.4189646, 0.4547722, 0.3722363, 0.3847851, 0.4082552, 0.4906771, 
    0.4824576, 0.5030468, 0.4984894, 0.4755728, 0.4125194, 0.3581249, 
    0.3000846, 0.2417517, 0.1705434, -0.02418327, -0.016078, -0.0734024, 
    -0.1254044, -0.1177559,
  -0.02634788, -0.04329109, -0.3344374, -0.3526011, -0.3947563, -0.365622, 
    -0.3748014, -0.3944306, -0.4217904, -0.451299, -0.4317675, -0.3856583, 
    -0.3029776, -0.1597643, -0.08803415, 0.007164478, 0.32165, 0.4457878, 
    0.5343131, 0.4413606, 0.3037794, 0.2282257, 0.2770529, 0.3025913, 
    0.2247105, 0.1541538, 0.07586575, -0.00190258, -0.08622837, -0.1421843, 
    -0.1741829, -0.2049608, -0.278481, -0.2787747, -0.3160133, -0.3540821, 
    -0.3347464, -0.2328095, -0.1099577, 0.03717756, 0.1339712, 0.1774282, 
    0.213057, 0.2806182, 0.230293, 0.1642448, 0.1451855, 0.1033398, 
    0.08514285, 0.03120458, -0.03787088, -0.1354295, -0.2417772, -0.3522753, 
    -0.4121387, -0.4250453, -0.377161, -0.2936978, -0.2277148, -0.1889451, 
    -0.2288537, -0.2931118, -0.3810511, -0.4851203, -0.5870897, -0.670293, 
    -0.6912239, -0.6664032, -0.5927703, -0.4835094, -0.2942352, -0.113034, 
    0.003616452, 0.1033724, 0.2336296, 0.3776562, 0.5559603, 0.7199576, 
    0.7172722, 0.6923534, 0.5543002, 0.6065137, 0.6576205, 0.7278355, 
    0.8128287, 0.8809764, 0.903584, 0.9588087, 1.022367, 1.092239, 1.114033, 
    1.059395, 0.9707388, 0.7638706, 0.5123897, 0.2564809,
  0.397334, 0.1333367, -0.06103194, -0.1462204, -0.2266078, -0.3278129, 
    -0.3858695, -0.3918912, -0.3282845, -0.2068489, -0.06392905, 0.01579106, 
    -0.03808272, -0.1807907, -0.3479135, -0.4697561, -0.5683889, -0.553317, 
    -0.4660611, -0.3341439, -0.1736133, 0.02189445, 0.1624218, 0.2626824, 
    0.2346873, 0.1881866, 0.1966338, 0.1966834, 0.1631382, 0.06411433, 
    -0.07641315, -0.1012831, -0.03154039, -0.222198, -0.1233211, -0.2725229, 
    -0.2623339, -0.2995412, -0.23473, -0.1001434, -0.002389669, 0.06600285, 
    0.1324087, 0.2173697, 0.2747591, 0.2959669, 0.2506706, 0.115905, 
    0.07295251, 0.1055858, 0.1516144, 0.01297522, -0.1030407, -0.2413218, 
    -0.3501108, -0.4469206, -0.4401662, -0.3429983, -0.2797983, -0.1928356, 
    -0.09802747, 0.01658845, 0.03486633, 0.02615857, -0.05063152, 
    -0.07270193, -0.11834, -0.1541963, -0.1635873, -0.1715457, -0.06042933, 
    0.132165, 0.3074739, 0.4361525, 0.5705601, 0.7214717, 0.915856, 1.093444, 
    1.292191, 1.249873, 0.8806676, 0.7873732, 0.8100452, 0.8902537, 
    0.9859892, 1.025361, 1.010843, 0.9976106, 1.020609, 1.080505, 1.173604, 
    1.201468, 1.165823, 1.037536, 0.861478, 0.6608106,
  1.601435, 1.429723, 1.228225, 1.122269, 1.076126, 1.026777, 0.9831407, 
    0.9618518, 1.014749, 1.101126, 1.217093, 1.31387, 1.342484, 1.315335, 
    1.244681, 1.233124, 1.221732, 1.169209, 1.041002, 0.9121611, 0.8846381, 
    1.011103, 1.18389, 1.369909, 1.414961, 1.324189, 1.19569, 1.23708, 
    1.293265, 1.219567, 1.098311, 0.9996777, 1.028356, 1.203747, 1.363691, 
    1.343102, 1.12598, 0.8643588, 0.7347363, 0.7187365, 0.7342479, 0.7818227, 
    0.7806184, 0.7430043, 0.7552767, 0.697968, 0.5214872, 0.3580594, 
    0.3490424, 0.4654322, 0.6132679, 0.6810412, 0.5949898, 0.3399925, 
    0.1126008, -0.0261035, 0.0004262924, -0.08448601, -0.190443, -0.1523571, 
    -0.04135466, 0.06277943, 0.09316683, 0.110013, 0.1989775, 0.2977242, 
    0.4056668, 0.4841666, 0.535924, 0.5332875, 0.5314322, 0.5611033, 
    0.5520701, 0.4813342, 0.3694367, 0.3067575, 0.3566923, 0.5659208, 
    0.8792839, 1.248457, 1.72528, 1.909004, 1.603323, 1.364049, 1.487829, 
    1.573473, 1.541866, 1.360599, 1.222139, 1.216279, 1.322301, 1.453388, 
    1.572952, 1.692272, 1.709508, 1.671829,
  1.843622, 1.75176, 1.718801, 1.654055, 1.49385, 1.283808, 1.103355, 
    1.063315, 1.08353, 1.068897, 0.9971046, 0.9511085, 0.9607453, 1.0647, 
    1.22912, 1.403226, 1.585907, 1.753925, 1.950296, 2.263186, 2.526825, 
    2.576353, 2.517433, 2.449318, 2.458205, 2.405014, 2.323211, 2.259703, 
    2.233319, 2.185272, 2.01802, 1.768525, 1.526402, 1.439439, 1.533076, 
    1.680634, 1.689618, 1.578063, 1.469485, 1.508775, 1.651662, 1.752525, 
    1.747301, 1.693606, 1.61522, 1.488365, 1.321584, 1.160907, 1.106772, 
    1.175164, 1.264179, 1.302248, 1.325132, 1.309898, 1.149368, 0.9329453, 
    0.7855983, 0.70788, 0.6067734, 0.5468616, 0.5421572, 0.5280786, 
    0.4951854, 0.5643744, 0.7477403, 0.8908229, 0.9342146, 0.9736843, 
    1.057278, 1.123652, 1.175833, 1.23192, 1.206903, 1.037926, 0.7977891, 
    0.6271996, 0.5322456, 0.4877958, 0.5542507, 0.7750835, 1.022805, 
    1.080146, 0.9630075, 0.8456731, 0.6598821, 0.6983261, 0.9050479, 
    1.222968, 1.551858, 1.588349, 1.52427, 1.627314, 1.812226, 1.977004, 
    2.007082, 1.939358,
  1.660971, 1.628695, 1.604884, 1.562453, 1.487095, 1.375995, 1.303778, 
    1.286575, 1.269306, 1.264049, 1.253632, 1.203681, 1.108891, 0.9727421, 
    0.8783236, 0.8980169, 1.005342, 1.094144, 1.122155, 1.175573, 1.289749, 
    1.458565, 1.667011, 1.951142, 2.259932, 2.459721, 2.476665, 2.339034, 
    2.18083, 2.061006, 1.896812, 1.644989, 1.37601, 1.191375, 1.082423, 
    1.076255, 1.145819, 1.196112, 1.214569, 1.306202, 1.517139, 1.729379, 
    1.910614, 2.046143, 2.105372, 2.1105, 2.079494, 1.98983, 1.916115, 
    2.022186, 2.232961, 2.339781, 2.376499, 2.437307, 2.440904, 2.299774, 
    2.142971, 1.995673, 1.851337, 1.733238, 1.705959, 1.640204, 1.512649, 
    1.478225, 1.526744, 1.516002, 1.434834, 1.389895, 1.412112, 1.363528, 
    1.303307, 1.329658, 1.338089, 1.19818, 0.9794774, 0.8079925, 0.6089869, 
    0.3842478, 0.2401719, 0.2408552, 0.3911805, 0.61343, 0.7508159, 
    0.6454124, 0.5499859, 0.5718932, 0.6583843, 0.7433939, 0.8424339, 
    0.9040871, 0.9431496, 1.012275, 1.125181, 1.286655, 1.443915, 1.595363,
  1.541164, 1.566734, 1.559784, 1.580601, 1.593215, 1.586494, 1.564, 
    1.455521, 1.252412, 1.068329, 0.9395046, 0.8241901, 0.7256708, 0.6349974, 
    0.5874214, 0.5979519, 0.6365271, 0.6575232, 0.632719, 0.6104364, 
    0.6523972, 0.7297726, 0.7970095, 0.8942099, 1.066851, 1.261885, 1.390579, 
    1.413854, 1.397676, 1.428243, 1.403048, 1.243641, 1.067419, 0.9698439, 
    0.8521347, 0.7056017, 0.6489611, 0.7174177, 0.8182473, 0.974628, 
    1.176189, 1.312257, 1.456511, 1.766489, 2.030015, 2.013137, 1.980666, 
    2.01426, 2.115383, 2.332782, 2.673733, 2.894745, 2.885403, 2.897398, 
    3.011265, 3.041279, 2.926858, 2.758694, 2.627981, 2.630195, 2.664797, 
    2.585159, 2.327997, 2.102558, 1.948717, 1.819843, 1.6744, 1.559915, 
    1.45609, 1.323896, 1.132067, 0.9646349, 0.8739443, 0.7892103, 0.7101898, 
    0.5927272, 0.3336945, 0.2573276, 0.1964865, 0.06100464, -0.1234841, 
    -0.07161283, 0.1306171, 0.2036643, 0.33008, 0.5560255, 0.6828318, 
    0.603632, 0.5112324, 0.5508652, 0.697073, 0.8811378, 1.01566, 1.096959, 
    1.217157, 1.407229,
  1.052834, 1.098603, 1.175605, 1.23454, 1.239553, 1.139732, 1.072773, 
    1.011168, 0.8469262, 0.6391778, 0.4427104, 0.2785339, 0.1970072, 
    0.1355324, 0.09756088, 0.1113634, 0.1653357, 0.2117062, 0.217452, 
    0.2592974, 0.340662, 0.3393602, 0.2519407, 0.2449265, 0.3459024, 
    0.4485874, 0.5271692, 0.6154823, 0.7034531, 0.7822456, 0.8223829, 
    0.8126822, 0.7422724, 0.6228876, 0.5249386, 0.454154, 0.387291, 
    0.3298206, 0.3170271, 0.4541035, 0.687469, 0.625278, 0.4466972, 
    0.6441417, 1.019989, 1.04927, 1.024612, 1.289374, 1.714765, 2.084915, 
    2.430276, 2.753063, 2.879527, 2.815465, 2.77038, 2.760777, 2.670478, 
    2.565986, 2.506985, 2.505749, 2.544729, 2.559264, 2.509361, 2.405048, 
    2.242954, 2.050979, 1.813349, 1.459605, 1.144338, 1.012275, 0.8619814, 
    0.731627, 0.6726103, 0.5765977, 0.4424009, 0.3200388, 0.1585317, 
    0.1206737, 0.1261244, 0.02339077, -0.2256827, -0.3906064, -0.432713, 
    -0.4735003, -0.4136205, -0.1751938, 0.1135931, 0.3369818, 0.533206, 
    0.6445332, 0.7150087, 0.8619823, 1.025605, 1.093166, 1.070868, 1.046226,
  0.7915711, 0.8695483, 0.8701506, 0.8827486, 0.9995451, 1.097609, 1.090594, 
    0.9794459, 0.7436385, 0.5627794, 0.4897485, 0.4352727, 0.3696475, 
    0.3037457, 0.2538743, 0.2161469, 0.2077169, 0.2101583, 0.09844112, 
    -0.1041155, -0.1908503, -0.2198048, -0.2388315, -0.1236944, 0.07251263, 
    0.1917677, 0.2047882, 0.1898146, 0.1853056, 0.1044788, -0.03354168, 
    -0.07930946, -0.05468464, -0.08009243, -0.08279324, -0.07527351, 
    -0.1254206, -0.1582155, -0.1722136, -0.1224265, -0.01373529, -0.1568017, 
    -0.3997707, -0.2675595, 0.1469588, 0.4005404, 0.3479197, 0.4190462, 
    0.7566109, 1.161201, 1.424352, 1.655895, 1.780553, 1.68874, 1.570055, 
    1.622008, 1.800866, 1.909947, 1.928421, 1.878632, 1.851223, 1.919502, 
    1.993183, 1.994322, 1.909508, 1.738837, 1.470966, 1.050507, 0.6961613, 
    0.4992867, 0.4240909, 0.4179549, 0.457571, 0.3605981, 0.1487818, 
    -0.0143857, -0.08562517, -0.01217103, 0.03721046, -0.06793499, 
    -0.1358223, -0.1868148, -0.2865219, -0.4732404, -0.6137991, -0.5870743, 
    -0.4316225, -0.14505, 0.2455258, 0.5867209, 0.8198748, 0.9260116, 
    0.9303083, 0.8724475, 0.7641463, 0.7134461,
  1.060923, 1.084751, 1.033238, 0.8933783, 0.7550807, 0.658824, 0.5408883, 
    0.5645208, 0.5604029, 0.4244008, 0.4233918, 0.4573598, 0.4182973, 
    0.3461618, 0.2738309, 0.1431508, -0.1160126, -0.3185196, -0.4635553, 
    -0.6648421, -0.7819161, -0.8217592, -0.8152976, -0.7643204, -0.6953106, 
    -0.5913868, -0.5091276, -0.5131645, -0.4386034, -0.3710413, -0.4041147, 
    -0.4510221, -0.506052, -0.4849424, -0.3808899, -0.4045229, -0.466795, 
    -0.4228001, -0.472476, -0.5318823, -0.569953, -0.8164692, -1.164076, 
    -1.251592, -1.069805, -0.7642384, -0.566761, -0.479131, -0.281312, 
    -0.04236341, 0.1782093, 0.3027701, 0.3657582, 0.3877311, 0.3290236, 
    0.3864937, 0.4901233, 0.5397167, 0.6524282, 0.7954946, 0.8934598, 
    0.964293, 0.9578314, 0.9624372, 0.9713244, 0.906383, 0.7870145, 
    0.6362004, 0.4724474, 0.3141141, 0.1773462, 0.02112913, -0.1219378, 
    -0.1808238, -0.126657, -0.1826468, -0.2866013, -0.1571093, -0.01313186, 
    0.01562834, 0.00924778, -0.07004881, -0.1671357, -0.3665333, -0.6193166, 
    -0.6164031, -0.4482718, -0.3473454, -0.2684069, -0.07475471, 0.235548, 
    0.4857922, 0.6272798, 0.7661471, 0.8408051, 0.9326348,
  0.6534204, 0.5053091, 0.4982128, 0.4299676, 0.2875519, 0.1295767, 
    -0.2046516, -0.1963999, 0.06880188, 0.07635403, 0.08389044, 0.2134471, 
    0.2316113, 0.06409836, -0.07418299, -0.1370248, -0.3826952, -0.7167445, 
    -1.003333, -1.236944, -1.360837, -1.423386, -1.433412, -1.400274, 
    -1.450974, -1.438523, -1.369644, -1.230451, -0.9770494, -0.9407372, 
    -0.9272771, -0.7311511, -0.6819639, -0.6618638, -0.5983219, -0.7050762, 
    -0.7066541, -0.4439259, -0.4626269, -0.6194301, -0.6832001, -1.043128, 
    -1.40081, -1.685837, -1.786357, -1.713164, -1.67275, -1.587399, 
    -1.489596, -1.428496, -1.300159, -1.22498, -1.140312, -0.9582975, 
    -0.890166, -0.7995574, -0.5957322, -0.586992, -0.6423309, -0.6907847, 
    -0.7447884, -0.6713998, -0.5789521, -0.4958138, -0.3912566, -0.2767873, 
    -0.1021454, 0.1255889, 0.2335155, 0.137991, -0.01233435, -0.1646452, 
    -0.3253224, -0.386797, -0.3498178, -0.3284636, -0.3419238, -0.2647104, 
    -0.26987, -0.1759083, -0.01596379, -0.1164356, -0.1593719, -0.1759737, 
    -0.3898892, -0.4613414, -0.3770967, -0.3608694, -0.4384413, -0.6042452, 
    -0.6372037, -0.4700165, -0.2093239, 0.1835151, 0.484426, 0.6292019,
  -0.1831999, -0.1043749, -0.05728853, -0.2054492, -0.2105925, 0.006725246, 
    -0.1051562, -0.2699021, -0.1895804, -0.2796192, -0.1711231, -0.2918261, 
    -0.5100554, -0.5788538, -0.7191863, -0.8873179, -1.034437, -1.113831, 
    -1.167363, -1.294593, -1.439678, -1.572913, -1.760039, -1.781312, 
    -1.678854, -1.550078, -1.388961, -1.266956, -1.089401, -1.127698, 
    -1.085609, -0.6269501, -0.4953909, -0.4163704, -0.3918262, -0.5003222, 
    -0.5627571, -0.5125946, -0.4860807, -0.5338346, -0.7747853, -1.20929, 
    -1.145521, -1.203203, -1.530059, -1.820358, -2.171432, -2.41432, 
    -2.536064, -2.568617, -2.420277, -2.259502, -2.039727, -1.793438, 
    -1.664873, -1.68167, -1.579017, -1.423532, -1.452243, -1.645342, 
    -1.847946, -1.851657, -1.730661, -1.494658, -1.172913, -0.9049931, 
    -0.6878383, -0.4802699, -0.3540659, -0.4019659, -0.4258265, -0.4951949, 
    -0.5873339, -0.6113251, -0.7475554, -0.7082001, -0.380661, -0.08202839, 
    -0.2881641, -0.3059538, -0.1686817, -0.2105436, -0.2672494, -0.2435514, 
    -0.4297982, -0.5508107, -0.6267872, -0.8147916, -0.9223435, -0.9596643, 
    -0.9970345, -0.9327605, -0.835218, -0.6413541, -0.459681, -0.3244762,
  -0.7085091, -0.5404589, -0.487969, -0.5047983, -0.1998341, 0.2400099, 
    0.3308949, 0.03777999, -0.2163379, -0.5723438, -0.4361296, -0.4643199, 
    -0.7223926, -0.7821259, -0.6204071, -0.5370085, -0.5665336, -0.663815, 
    -0.7043753, -0.8516731, -1.123207, -1.202471, -1.316761, -1.340101, 
    -1.232354, -1.205091, -1.125306, -1.097979, -1.059762, -1.049492, 
    -0.9088511, -0.5674284, -0.5381803, -0.4742154, -0.50125, -0.4942187, 
    -0.4009733, -0.4199186, -0.399899, -0.3619596, -0.5610156, -0.9805794, 
    -1.022165, -1.079636, -1.426934, -1.775339, -2.125664, -2.419724, 
    -2.623304, -2.663474, -2.575827, -2.308021, -1.911666, -1.746334, 
    -1.616094, -1.649655, -1.779538, -1.764564, -1.81318, -1.957028, 
    -2.089222, -2.038897, -1.871026, -1.619121, -1.481931, -1.397702, 
    -1.383981, -1.385462, -1.210479, -1.186537, -1.030059, -0.9322396, 
    -1.004473, -0.81611, -0.6932909, -0.4730113, -0.07473612, 0.2820344, 
    0.1491569, -0.07895184, -0.1319956, -0.2279266, -0.3059212, -0.2123014, 
    -0.4974577, -0.8183236, -0.7777636, -0.8153776, -1.073874, -1.087074, 
    -1.119658, -1.146335, -1.046367, -0.9776172, -0.8818164, -0.8155404,
  -0.9190886, -0.7340789, -0.540622, -0.2677379, 0.08509439, 0.2034372, 
    0.1624222, -0.1707815, -0.3575162, -0.5604134, -0.7362113, -0.388864, 
    -0.5108042, -0.75125, -0.6660457, -0.5774388, -0.3910146, -0.3961415, 
    -0.4206696, -0.4564281, -0.7632642, -0.9043612, -0.9893212, -1.117153, 
    -1.009292, -0.9360814, -0.9277482, -0.8237767, -0.7047496, -0.7273567, 
    -0.6585255, -0.4920056, -0.4029589, -0.3501108, -0.46541, -0.4852993, 
    -0.333379, -0.2324023, -0.2299938, -0.3780564, -0.4553351, -0.4948213, 
    -0.6864066, -0.9072237, -1.135153, -1.355531, -1.611472, -1.874574, 
    -1.94072, -1.710609, -1.599981, -1.546888, -1.32542, -1.26974, -1.140118, 
    -1.151039, -1.264629, -1.302667, -1.312204, -1.341338, -1.420569, 
    -1.410478, -1.407728, -1.430335, -1.607061, -1.604977, -1.552878, 
    -1.581019, -1.288848, -1.085788, -0.8108206, -0.5776174, -0.5756481, 
    -0.4399548, -0.2945118, 0.1092968, 0.3032587, 0.2206903, 0.05386078, 
    -0.06757489, -0.04747438, -0.006946683, -0.2706509, -0.240101, 
    -0.4423633, -0.8983204, -0.9218397, -0.6792939, -0.8214648, -0.7964485, 
    -0.8197396, -0.9349742, -0.9354627, -1.035674, -1.036618, -0.9487114,
  -0.5522919, -0.3868623, -0.1206186, 0.1984737, 0.2380731, 0.2029495, 
    0.1641312, -0.2235808, -0.2586558, -0.187578, -0.2787893, 0.01155913, 
    -0.04355156, -0.1542777, -0.04171276, -0.2773266, -0.1937003, 0.05029535, 
    0.005486488, -0.1110659, -0.3223124, -0.4559875, -0.5374327, -0.6963196, 
    -0.763947, -0.6301737, -0.6451969, -0.6595531, -0.4565744, -0.2843885, 
    -0.2787085, -0.2460589, -0.1891251, -0.1002898, -0.250371, -0.1897268, 
    -0.1118622, 0.0300324, -0.02136731, -0.2272918, -0.3120737, -0.2509751, 
    -0.3605118, -0.5344863, -0.6905899, -0.8972306, -1.016892, -1.115281, 
    -1.103611, -0.8795872, -0.6563606, -0.5800586, -0.5067675, -0.4350555, 
    -0.3818653, -0.4526174, -0.5706513, -0.5979624, -0.4614227, -0.4594858, 
    -0.6447723, -0.8792777, -1.20169, -1.308119, -1.431149, -1.454115, 
    -1.279131, -1.147669, -0.8983693, -0.5942678, -0.3804173, -0.2906709, 
    -0.2389455, -0.002178192, 0.0815134, 0.4450551, 0.4465857, -0.1196092, 
    -0.1435027, -0.132386, -0.08359063, 0.02202487, -0.2853487, -0.1317515, 
    -0.1121871, -0.2238247, -0.1625781, -0.1965461, -0.4640603, -0.5803523, 
    -0.6913061, -0.8005672, -0.9105768, -0.9172173, -0.8925261, -0.7436495,
  -0.2001758, -0.1804655, -0.08027005, 0.0417676, 0.08431315, 0.02267623, 
    0.1555537, 0.02454734, -0.2219861, -0.1757454, -0.1455534, 0.08791015, 
    0.08055329, -0.06051135, 0.007132053, -0.02766848, -0.0249815, 
    0.09520149, 0.1715355, 0.0347681, -0.05043793, -0.07949066, -0.2225723, 
    -0.2363424, -0.3966446, -0.365818, -0.2669253, -0.3355451, -0.2362132, 
    0.04552555, 0.1065607, 0.1633472, 0.4083023, 0.2475615, 0.0950551, 
    -0.05328465, -0.02253914, 0.1604347, -0.02644539, 0.005714893, 
    0.04054451, 0.05107594, -0.02118969, -0.08626032, -0.1703429, -0.3687472, 
    -0.4649067, -0.4957004, -0.4795709, -0.4404435, -0.2749977, -0.06254578, 
    0.04515266, 0.07597923, 0.1383491, 0.213789, 0.2620797, 0.1734896, 
    0.1629748, -0.04906893, -0.3339486, -0.561748, -0.8432908, -0.9375134, 
    -0.9490857, -0.8681293, -0.6991024, -0.4286432, -0.3358698, -0.1806455, 
    -0.103075, 0.05566692, 0.1412296, 0.2591333, 0.2554717, 0.3904489, 
    0.2682486, -0.01425457, 0.1467969, -0.002275348, -0.1186003, -0.07621765, 
    -0.08632469, 0.03125286, -0.05426145, 0.02267575, 0.4013853, 0.2161307, 
    -0.0276022, -0.1740866, -0.490119, -0.5217438, -0.5949697, -0.479198, 
    -0.4719048, -0.3419247,
  -0.01578474, 0.09067678, 0.1017282, -0.03020509, 0.04245114, 0.1006546, 
    0.2155473, 0.1521189, -0.02340174, 0.003421068, -0.22861, -0.04866195, 
    -0.08163738, -0.2793918, 0.003746033, 0.1394548, 0.2051282, 0.1849132, 
    0.3675961, 0.3098817, 0.2146993, 0.2432151, 0.1346865, 0.2969413, 
    0.3016133, 0.2626157, 0.2759786, 0.3055196, 0.3745303, 0.4803085, 
    0.4252791, 0.4980483, 0.6645522, 0.6650081, 0.509572, 0.1973011, 
    0.02529621, 0.078403, 0.07749319, 0.213397, 0.1757178, 0.2089872, 
    0.1732111, -0.01134157, -0.1249647, -0.2227187, -0.1728163, -0.03619528, 
    0.046422, 0.2526555, 0.4808292, 0.6132193, 0.644567, 0.5782909, 
    0.5704622, 0.4610219, 0.4611683, 0.3098984, 0.1587591, 0.02148724, 
    -0.1104302, -0.2355609, -0.4018693, -0.511651, -0.4642224, -0.3110161, 
    -0.3252273, -0.1738105, -0.1006012, 0.04425573, 0.1084328, 0.3297877, 
    0.2959824, 0.2558784, 0.323441, 0.1496289, 0.09124672, -0.2567024, 
    -0.02507815, -0.01069012, -0.0191862, -0.01801443, 0.01207972, 
    0.05778289, 0.02388, 0.1446483, 0.5819674, 0.4984722, 0.2696633, 
    0.2784848, 0.01147652, -0.02716303, -0.07070208, -0.03701067, 
    -0.04435062, -0.004164219,
  0.1025908, 0.1966345, 0.2252799, 0.3072787, 0.3148466, 0.04977536, 
    0.212568, 0.1790233, 0.04865217, -0.007955551, -0.1870085, -0.1059213, 
    -0.2628388, -0.3438611, 0.04616165, 0.05031252, 0.1556988, 0.2108912, 
    0.3784032, 0.5293474, 0.6495624, 0.5891628, 0.4559269, 0.5025749, 
    0.667695, 0.9206901, 0.9367852, 1.019419, 0.8635936, 0.9928894, 0.904233, 
    0.6436863, 0.5938816, 0.6108904, 0.5308452, 0.4915385, 0.2766123, 
    -0.06943083, -0.05360985, 0.05259109, 0.1285026, 0.1383166, 0.1882029, 
    0.1183462, 0.1997914, 0.1879911, 0.2456737, 0.5079293, 0.4230013, 
    0.2843285, 0.3083687, 0.4314966, 0.4784846, 0.4362321, 0.3979993, 
    0.2702656, 0.2609224, 0.2172542, 0.1115899, 0.05686998, -0.07748938, 
    -0.2340808, -0.2863593, -0.3422189, -0.3623199, -0.3625965, -0.2778797, 
    -0.1043611, 0.004656792, 0.1084652, 0.1298203, 0.1417179, 0.1769562, 
    0.1337922, 0.2611849, 0.4022493, 0.05693674, -0.2302864, -0.06514975, 
    -0.0252409, -0.04260737, 0.003762901, 0.01160789, 0.01352859, 0.1009634, 
    0.1548531, 0.2330437, 0.6743674, 0.5825863, 0.5944839, 0.4619322, 
    0.3667169, 0.270721, 0.2619967, 0.1967311, 0.12012,
  0.4508171, 0.5213578, 0.5181507, 0.6886424, 0.8137402, 0.3067415, 
    0.1576529, 0.3413117, 0.107604, 0.1716175, 0.001565814, -0.1203254, 
    0.02278996, -0.04503274, -0.05784202, 0.0389843, 0.136673, 0.1250846, 
    0.19346, 0.2749052, 0.5034046, 0.4641469, 0.3060741, 0.03524113, 
    0.274385, 0.8210812, 1.051517, 0.9468291, 0.4936556, 1.078079, 1.156839, 
    0.8616714, 0.6525092, 0.6103873, 0.7814324, 0.6144891, 0.3508661, 
    0.02220376, -0.05634433, 0.03159499, 0.116556, -0.005579472, -0.04503298, 
    -0.09695339, 0.08657503, 0.1475942, 0.08615208, 0.2989128, 0.4063344, 
    0.2657583, -0.01630545, 0.002607346, 0.14639, 0.302526, 0.3153186, 
    0.2264352, 0.1040878, 0.0517602, 0.02869654, 0.003273964, -0.007469177, 
    -0.08328295, -0.1521306, -0.264256, -0.209065, -0.2018051, -0.1287584, 
    -0.09070396, 0.05869389, 0.05071878, 0.1693878, 0.2279816, 0.3479033, 
    0.1790233, 0.3497754, 0.5715363, -0.2378063, 0.01725585, -0.0330534, 
    -0.04651368, -0.07017899, -0.05719078, -0.08121419, 0.0932976, 0.3093946, 
    0.1796744, 0.3231641, 0.8717155, 0.8247428, 0.8026562, 0.63026, 
    0.5509634, 0.3505077, 0.3605337, 0.4098988, 0.3322134,
  0.5355176, 0.5605824, 0.4695508, 0.310078, 0.3083692, 0.200166, 0.03262044, 
    0.1334505, 0.1088734, 0.2704785, 0.4064809, -0.2516569, -0.1034636, 
    0.1928581, 0.1312044, 0.1150261, 0.09629226, 0.06460261, -0.02454066, 
    -0.07944012, 0.1381379, 0.2378126, 0.09087238, -0.3432097, -0.4939746, 
    -0.1611621, 0.3041049, 0.2734897, -0.02268559, 0.5915557, 0.234069, 
    0.05081703, -0.005498052, 0.05307961, 0.3282422, 0.06172201, -0.02485028, 
    -0.04819012, -0.02707994, 0.3408072, 0.04787159, -0.3026336, -0.2669889, 
    -0.2059538, -0.1262826, -0.03665066, 3.457069e-006, 0.1238315, 0.4237177, 
    0.7004588, 0.689033, 0.7155793, 0.7357941, 0.8708525, 0.8589387, 
    0.7128448, 0.5659523, 0.382587, 0.2246118, 0.02965784, -0.07110739, 
    -0.1829562, -0.196775, -0.2191381, -0.1605439, -0.2180963, -0.0867157, 
    -0.002015114, 0.170397, 0.1708851, 0.298229, 0.2756543, 0.2998406, 
    0.1709017, 0.5267286, 0.6485059, -0.1291962, 0.025166, -0.03066084, 
    -0.05769527, -0.06894195, -0.05619788, -0.1893196, -0.1637499, 
    -0.0440886, 0.1418655, 0.6436884, 0.9920772, 0.7960643, 0.7320184, 
    0.5399938, 0.6929071, 0.4984252, 0.4552119, 0.5898149, 0.5815628,
  0.5419793, 0.4938184, 0.4411005, 0.1492221, 0.04979166, 0.09676439, 
    0.09243488, 0.132653, 0.02853514, 0.2167838, 0.609118, 0.09472981, 
    -0.2671195, -0.07706404, 0.2587597, 0.1677444, 0.0340364, -0.1301237, 
    -0.33792, -0.3098926, -0.142184, -0.1638477, -0.2969043, -0.3204236, 
    -0.5449839, -0.483086, -0.1650844, -0.09062177, -0.2062306, 0.1567741, 
    0.08032554, 0.008710925, -0.02146487, -0.2966766, -0.3230436, -0.3571419, 
    -0.3419561, -0.2280245, -0.02851272, -0.003317118, -0.253773, -0.3143685, 
    -0.2153124, -0.1327608, -0.163229, -0.2376435, -0.2647758, -0.2631481, 
    -0.2658985, -0.1877737, -0.09656286, 0.1079297, 0.2509308, 0.3661981, 
    0.4140654, 0.3689804, 0.3387074, 0.2971215, 0.3194532, 0.2501984, 
    0.193574, 0.1291208, -0.02515936, -0.09247732, -0.09169626, -0.186667, 
    -0.1205862, -0.1406538, -0.03458309, 0.08133435, 0.2117219, 0.3007519, 
    0.4547232, 0.2222852, 0.09907579, 0.1038444, 0.01956689, -0.009567052, 
    -0.0005013123, 0.00926432, 0.1771516, 0.04533213, -0.4440396, -0.5354297, 
    -0.2265592, 0.08841467, 0.6662956, 1.028991, 0.8740104, 0.5962758, 
    0.2004913, 0.3053255, 0.472334, 0.5615104, 0.5603549, 0.6517286,
  -0.00741899, 0.1254265, 0.08179027, 0.08388996, 0.1323435, 0.1577344, 
    0.2258008, 0.08454072, 0.08828449, 0.4230664, 0.2949577, 0.2126008, 
    -0.1066701, -0.4002085, -0.04137182, 0.1178255, -0.05470085, -0.4776988, 
    -0.5734339, -0.5271616, -0.4558415, -0.2597642, -0.2346168, -0.3644676, 
    -0.6645823, -0.5202434, -0.112025, -0.1624479, -0.2242481, -0.2692516, 
    -0.3245735, -0.09395835, -0.001510382, -0.2661263, -0.7476041, 
    -0.3877735, -0.2843719, -0.3419569, -0.2226532, -0.4745897, -0.5488249, 
    -0.4079555, -0.2288866, -0.192461, -0.3263316, -0.3258433, -0.3003716, 
    -0.2438288, -0.2974095, -0.3267226, -0.3446264, -0.3248186, -0.2239885, 
    -0.2796197, -0.2675433, -0.2572889, -0.2046356, -0.1756477, -0.07486677, 
    -0.0905242, -0.1704721, -0.1836724, -0.2338673, -0.1102668, -0.0287239, 
    -0.06054364, -0.08499023, -0.05621421, -0.09158212, -0.07987988, 
    0.1762241, 0.1605337, -0.1339488, -0.3973112, -0.1951792, 0.02316405, 
    0.2896194, 0.201761, 0.2149935, -0.04731131, 0.001386881, -0.3336232, 
    -0.4426074, 0.1162953, 0.611201, 0.7337439, 0.8853872, 0.8874381, 
    0.7737012, 0.5316762, 0.149971, 0.05871105, 0.3018584, 0.3935902, 
    0.1200391, 0.06868821,
  -0.1795052, 0.03956997, 0.07225251, 0.344111, 0.475329, 0.2917349, 
    0.303617, 0.2725616, 0.1233594, 0.2619825, 0.2164909, 0.1243846, 
    0.3001823, -0.02631545, -0.1304502, -0.1830711, -0.2675276, -0.5258121, 
    -0.6640124, -0.4614725, -0.2224102, -0.2439108, -0.3505659, -0.6277962, 
    -0.8783512, -0.7328596, -0.628058, -0.3831182, -0.372653, -0.6236625, 
    -1.216697, -1.125468, -0.1479948, 0.005895168, -0.6165655, -0.3077931, 
    -0.1640915, -0.10304, -0.02732372, -0.3118134, -0.2926726, -0.05828142, 
    0.1409698, 0.07265854, 0.02203941, 0.1739597, 0.2164087, 0.1713233, 
    0.08860874, 0.0312686, 0.04726744, 0.06910992, 0.166018, 0.1018577, 
    0.1543965, 0.08857536, 0.04762506, 0.009003162, -0.07625103, -0.1460252, 
    -0.285023, -0.3756154, -0.3964159, -0.3582486, -0.6026823, -0.836146, 
    -0.8321095, -0.6273564, -1.004326, -1.089173, -0.7117156, -0.996644, 
    -1.465068, -1.163555, -0.1400195, 0.0909701, 0.06639338, 0.01771188, 
    0.02907205, -0.2858057, -0.3102045, -0.3065257, -0.003968716, 0.5841012, 
    0.6097198, 0.5371449, 0.6289744, 0.488529, 0.4929881, 0.3958855, 
    0.2530305, 0.05900383, -0.02878952, 0.1985545, 0.04751289, -0.05308926,
  0.2310414, 0.4214391, 0.6465034, 0.814147, 0.5202669, 0.1256379, 0.2496775, 
    0.3360222, -0.02895176, 0.2294629, 0.4508979, 0.2578647, 0.4352082, 
    0.09538066, -0.08459997, -0.07831812, -0.1368132, -0.2230444, -0.2553186, 
    -0.06438589, -0.07288218, -0.4353328, -0.5183249, -0.680727, -0.8666487, 
    -0.7670393, -0.4141245, -0.199964, -0.4421678, -0.886894, -1.837138, 
    -1.945634, -1.158753, -0.6214812, -0.4737436, -0.1651499, -0.09280252, 
    -0.08015609, -0.1529751, -0.4134085, -0.4562793, -0.1359186, 0.0560236, 
    0.08878851, 0.3520532, 0.414732, 0.3310409, 0.1296411, 0.1156597, 
    0.1229506, 0.1215515, 0.06105423, -0.02804089, -0.08427525, -0.04299927, 
    -0.04897213, -0.1179829, -0.1989889, -0.2768707, -0.2839494, -0.2610817, 
    -0.2146454, -0.3273568, -0.5632131, -0.8516244, -1.015736, -1.132907, 
    -1.140589, -1.289629, -0.8568978, -0.7130339, -1.116891, -0.8236949, 
    -0.5406055, -0.3218079, -0.2723265, -0.1670208, -0.1442347, -0.09617233, 
    -0.1044741, -0.001935005, 0.1711936, 0.4285822, 0.4601426, 0.4497089, 
    0.5381374, 0.5078969, 0.4109893, 0.4565787, 0.3726108, 0.3481966, 
    0.405895, 0.7959666, 0.6098992, 0.003893137, 0.06162429,
  0.6003939, 0.6523147, 0.6393264, 0.4094759, 0.01593745, -0.01977193, 
    0.2074251, 0.2516797, 0.285306, 0.5723991, 0.3536327, 0.5217155, 
    0.7502147, 0.07980454, -0.2347787, -0.006230354, 0.2043962, 0.1864443, 
    0.2499704, 0.2200861, 0.03068256, -0.3198066, -0.7673469, -0.8956189, 
    -0.6740692, -0.289222, 0.132197, -0.1373177, -0.8086233, -1.485983, 
    -1.653903, -1.173581, -1.198206, -0.8837205, -0.2051725, 0.0103873, 
    -0.1643038, -0.400306, -0.5239062, -0.6860161, -0.5240045, -0.1077785, 
    0.1387396, 0.3137064, 0.5614443, 0.47715, 0.4256368, 0.3237162, 0.266685, 
    0.1975117, 0.1866555, 0.1135111, 0.03984594, 0.07848549, -0.02880621, 
    -0.1242166, -0.1799784, -0.2131162, -0.249413, -0.2756987, -0.3481092, 
    -0.4221487, -0.5415497, -0.6625619, -0.6988416, -0.6041797, -0.5559376, 
    -0.5185188, -0.5033659, -0.05385417, 0.1452506, -0.1463671, -0.4162238, 
    -0.2193832, -0.08876705, 0.06974697, 0.1265345, 0.05394363, -0.01977253, 
    0.03864193, 0.1757832, 0.2454772, 0.3566427, 0.3459654, 0.46701, 
    0.4112821, 0.3491879, 0.3741064, 0.3700876, 0.365921, 0.4622266, 
    0.8181343, 1.305097, 0.6625846, 0.07134113, 0.3178907,
  0.1399284, -0.0004037023, -0.1873013, -0.2028286, -0.1765432, -0.02008128, 
    0.09901023, 0.2489128, 0.5347688, 0.4908886, 0.5355825, 0.8179557, 
    0.8815135, 0.2626333, -0.3242648, -0.2985644, 0.1985872, 0.264894, 
    0.2435732, 0.2799826, 0.0833683, -0.6147757, -0.7826792, 0.07207346, 
    0.4121941, 0.1719108, 0.01699543, -0.2094858, -0.148011, -0.4384409, 
    0.02785134, 0.4539092, -0.2407687, -0.1532845, 0.007392883, -0.3225882, 
    -0.8299286, -0.9835906, -0.8511851, -0.8179169, -0.2586889, 0.202867, 
    0.4706721, 0.512485, 0.4198909, 0.335907, 0.310565, 0.3185244, 0.2526388, 
    0.1477885, 0.1252136, 0.110043, 0.1818051, 0.2125177, 0.07068825, 
    -0.03513765, -0.05680132, -0.05673742, -0.1497064, -0.1468735, -0.176755, 
    -0.2480278, -0.2851369, -0.3902316, -0.4652801, -0.4050912, -0.1455207, 
    0.0994339, 0.06613278, -0.04473954, 0.225801, -0.349427, -0.8143849, 
    -0.05299282, 0.3021998, 0.213006, 0.0308938, -0.02584457, 0.03131723, 
    0.01406479, 0.2038431, 0.3177428, 0.4035172, 0.4501805, 0.4143248, 
    0.3475933, 0.3989935, 0.3985205, 0.3866878, 0.4528837, 0.4091177, 
    0.4563507, 0.4035514, 0.04943383, -0.02330422, 0.1341341,
  -0.2152963, -0.1107228, -0.2734344, -0.371335, -0.497246, -0.2637501, 
    -0.1088673, 0.005341768, 0.3895052, 0.392028, 0.4513542, 0.7868683, 
    0.3714876, 0.2157906, -0.03879881, -0.2131804, -0.05854166, 0.0519886, 
    0.144094, 0.3818059, -0.3459601, -1.150094, -0.6791309, 0.1720248, 
    0.3289908, 0.04987311, -0.1495086, 0.3273633, 0.788561, 0.2981315, 
    0.4652704, 0.5247594, 0.196764, 0.7282425, 0.5764683, 0.01754904, 
    -0.5422335, -0.5822396, -0.4990368, -0.5504525, -0.02807331, 0.2872586, 
    0.4394722, 0.324954, 0.2720566, 0.2929554, 0.1559596, 0.1283879, 
    0.08274984, 0.07168198, -0.0449357, -0.1805477, -0.157517, -0.2522111, 
    -0.2744274, -0.241128, -0.1569972, -0.003807068, 0.09186363, 0.1377301, 
    0.1128612, 0.1436877, 0.1038933, -0.04900384, -0.1241504, 0.002948999, 
    0.06012678, 0.2093129, 0.09495771, -0.05632794, -0.1780405, -0.902699, 
    -0.6807108, 0.3367381, -0.04329109, -0.4055476, -0.2555313, -0.1639948, 
    0.02169895, 0.05765295, 0.2248893, 0.3549023, 0.4534206, 0.4896665, 
    0.4116879, 0.3105807, 0.1503921, 0.1154151, 0.1484556, 0.185288, 
    0.2799993, 0.3308136, 0.2416537, 0.1374707, -0.02629884, -0.3106412,
  -0.009502053, -0.09348643, -0.4069631, -0.5024544, -0.6911917, -0.4675421, 
    -0.3357878, -0.3344533, 0.2169141, 0.3663282, 0.03852844, 0.0669629, 
    0.2656771, 0.3162794, 0.1585319, 0.07207358, 0.1589876, 0.1583853, 
    0.01160789, -0.06015298, -0.5924773, -0.5493132, 0.3087437, 0.4387889, 
    0.2448763, 0.04632485, -0.2176726, 0.4021842, 0.5816925, 0.2026073, 
    0.6572461, 0.842386, 0.8576853, 1.235485, 1.03485, 0.4914094, 0.08817041, 
    0.03642881, 0.01733708, 0.02135766, 0.2592642, 0.2660191, 0.1244826, 
    -0.1305301, -0.2032359, -0.2942839, -0.3624644, -0.2403615, -0.2671843, 
    -0.329294, -0.4364228, -0.4863739, -0.4985971, -0.5816216, -0.5733204, 
    -0.4870572, -0.3114715, -0.1998506, -0.09928083, 0.07184553, 0.2091827, 
    0.3600786, 0.3220084, 0.2007682, -0.008444309, 0.007099152, 0.3112335, 
    0.008125067, -0.232305, -0.005319357, -0.1213837, -0.3987117, 0.1467481, 
    0.5247589, 0.083125, -0.1668423, -0.2281871, -0.3217416, -0.3121876, 
    -0.2350228, -0.02091146, 0.1309111, 0.2126007, 0.229707, 0.1698437, 
    0.07685852, -0.02668953, -0.05878639, -0.1848121, -0.2496071, -0.1494441, 
    -0.01609373, 0.1852574, 0.2331901, 0.09202814, -0.01762371,
  0.1202995, -0.2567024, -0.7626598, -0.8615692, -0.6996388, -0.2827441, 
    -0.02970049, 0.205651, 0.3066601, 0.1749547, -0.1387825, 0.1363801, 
    0.5426302, 0.2470574, -0.04366538, -0.09226596, 0.1150094, 0.08678699, 
    -0.2605599, -0.1888151, 0.003942251, 0.07070637, 0.07435203, -0.4965787, 
    -0.5064418, -0.5038707, -0.4654911, 0.2253121, 0.2493198, -0.08398104, 
    0.2514192, 0.3651073, 0.3659211, 0.6909862, 0.8010774, 0.6643425, 
    0.5763704, 0.6127638, 0.6004752, 0.6556672, 0.5140007, 0.2109731, 
    -0.09918296, -0.4042937, -0.5804819, -0.7710905, -0.8340951, -0.723776, 
    -0.7363737, -0.7986132, -0.8823047, -0.8656217, -0.8295701, -0.784681, 
    -0.6412404, -0.4943813, -0.3435349, -0.2900193, -0.1827276, -0.03201175, 
    0.09529972, 0.2574576, 0.3003614, 0.3126335, 0.05810785, -0.03962898, 
    0.2082067, 0.0273633, -0.1481901, 0.1824899, 0.1051462, 0.03548515, 
    0.1776562, 0.127754, -0.1026009, -0.2560188, -0.2184048, -0.1298143, 
    -0.1619107, -0.1786914, -0.1458625, -0.2532683, -0.3144987, -0.3089323, 
    -0.3673471, -0.440752, -0.5138476, -0.6627088, -0.7785943, -0.7597139, 
    -0.7174125, -0.460674, -0.06834006, 0.007197142, 0.1216829, 0.1782096,
  -0.7433235, -0.7489225, -0.6300749, -0.4095507, -0.1462696, 0.2532583, 
    0.7320831, 0.6841992, 0.276094, 0.009605885, 0.3925164, 0.6745634, 
    0.4586133, -0.2105436, -0.3865529, -0.3068978, -0.2386526, -0.07991219, 
    -0.04239583, 0.2358756, 0.4721544, 0.1956087, -0.02455723, -0.01594746, 
    0.07117832, 0.1545606, 0.3246614, 0.4545767, 0.1846875, -0.218356, 
    -0.3354294, -0.4232878, -0.4304817, -0.2637174, -0.3021778, -0.2520965, 
    -0.03012395, 0.13638, 0.2050817, 0.3208365, 0.2979529, 0.118037, 
    -0.1134243, -0.4011359, -0.6778452, -0.874948, -0.9160125, -0.8908498, 
    -0.9191532, -0.9710736, -1.048824, -0.9854133, -0.9246057, -0.8524055, 
    -0.6654755, -0.5127409, -0.4284961, -0.377308, -0.1915658, -0.04667645, 
    -0.009664722, 0.1486686, 0.2725942, 0.01914358, -0.05328465, -0.08422518, 
    -0.03321588, -0.09994781, -0.07900059, -0.01544273, -0.09612298, 
    -0.05683269, -0.1207486, -0.3132781, -0.3715625, -0.2590461, -0.2177703, 
    -0.3217907, -0.5441537, -0.6190076, -0.6655407, -0.6556933, -0.6444628, 
    -0.7269988, -0.908541, -1.080774, -1.111992, -1.145489, -1.234111, 
    -1.291842, -1.286553, -1.014466, -0.5965136, -0.1636686, 0.1181023, 
    -0.2001595,
  -1.483053, -0.9274871, -0.116875, 0.03148103, -0.01000619, 0.1369662, 
    0.3240266, -0.03368855, -0.1331513, 0.2182162, 0.3241568, 0.1627473, 
    -0.1616992, -0.7043915, -0.4698698, -0.2341276, -0.2228483, -0.08446932, 
    0.1536491, 0.2288442, -0.07657553, -0.1784799, 0.277705, 0.3633659, 
    0.3483917, 0.3266959, 0.5477247, 0.2532097, -0.1129525, -0.3224903, 
    -0.5041799, -0.5426564, -0.495993, -0.5182261, -0.5311166, -0.5190883, 
    -0.3888803, -0.1223115, -0.07061887, 0.09359026, 0.3255563, 0.2434926, 
    -0.08027029, -0.3931286, -0.6857066, -0.9206836, -0.9443493, -0.8967905, 
    -0.9281869, -0.9130015, -0.8369274, -0.7555633, -0.6685843, -0.5569305, 
    -0.4776175, -0.4332488, -0.3526821, -0.2839808, -0.1684864, -0.02403641, 
    0.06561184, 0.164717, 0.1714873, 0.1326041, -0.1193981, -0.2043425, 
    -0.120358, -0.03787148, -0.0487597, -0.2121549, -0.1938769, 0.04679686, 
    0.05340499, -0.1655082, -0.2173307, -0.2447069, -0.4578743, -0.7300913, 
    -0.7018523, -0.5733371, -0.4997687, -0.4517221, -0.6301079, -0.936553, 
    -1.094609, -1.251364, -1.251266, -1.229147, -1.394349, -1.415736, 
    -1.304716, -1.330253, -1.225892, -0.5333951, -0.05611634, -0.794886,
  -0.6863737, -0.2878223, -0.1455863, -0.1000785, -0.09418619, 0.04507148, 
    0.1535838, -0.01103181, 0.1336293, 0.3754101, 0.05680668, -0.2748177, 
    -0.1843555, -0.0005338788, 0.1737012, 0.3297396, 0.07710284, -0.03477866, 
    0.1188835, 0.03986327, -0.2295541, -0.306361, -0.1150521, -0.03398103, 
    -0.03588539, 0.2078316, 0.4040394, 0.06346363, -0.3538704, -0.4239712, 
    -0.3230112, -0.158623, 0.02838874, 0.1605825, 0.1101758, 0.006985545, 
    0.09746385, 0.2364615, 0.1442904, -0.03134441, -0.1459439, -0.3287888, 
    -0.5489714, -0.6916635, -0.8028941, -0.9101694, -0.969821, -1.060218, 
    -1.185723, -1.156003, -0.9109998, -0.5873342, -0.271872, 0.02861643, 
    0.111917, 0.009686947, -0.04153347, -0.01632214, 0.08693337, 0.2432485, 
    0.1848176, 0.02570295, -0.1119432, -0.1286099, -0.2496063, -0.3000619, 
    -0.2176237, -0.1580859, -0.1510547, -0.2643196, -0.2154427, 0.00854817, 
    0.06837888, -0.09649742, -0.3347945, -0.3264942, -0.3680468, -0.3141408, 
    -0.1706512, -0.1045871, -0.07965183, -0.03482771, -0.2435193, -0.5581188, 
    -0.6925588, -0.8116341, -0.9210744, -1.08556, -1.294007, -1.267982, 
    -1.133688, -1.200567, -1.208428, -0.9282843, -0.7363575, -0.6826629,
  0.07698905, 0.03830075, 0.107718, 0.2857454, 0.3877474, 0.4882846, 
    0.6863151, 0.6445346, 0.4961132, 0.4167839, 0.3795928, 0.6448761, 
    1.039164, 1.049027, 0.636429, 0.2294467, -0.1182259, -0.1914356, 
    -0.1912728, -0.1930143, -0.05741864, 0.06146166, 0.0636263, 0.1527376, 
    0.1889027, 0.1625681, -0.04654616, -0.2822233, -0.2450004, 0.03104162, 
    0.284443, 0.4165075, 0.5117378, 0.4465039, 0.3410512, 0.327168, 
    0.3758171, 0.3572624, 0.3590365, 0.2029654, -0.02065146, -0.1741016, 
    -0.3537891, -0.5642381, -0.7127404, -0.780303, -0.8759735, -1.014255, 
    -1.079977, -1.025664, -0.8362598, -0.4809537, -0.05396795, 0.2919626, 
    0.4645209, 0.5551949, 0.6267447, 0.6947782, 0.7043974, 0.5897491, 
    0.2866569, -0.03243518, -0.1766891, -0.196237, -0.266794, -0.1942186, 
    0.0413121, 0.2385123, 0.336966, 0.3288119, 0.1762403, 0.004039705, 
    -0.1098763, -0.1448861, -0.09563482, -0.1260056, -0.2048795, -0.213994, 
    -0.06829083, 0.1163607, 0.1648955, 0.1009796, 0.05456066, 0.0300808, 
    -0.1409311, -0.3550425, -0.593389, -0.7859993, -0.8270965, -0.6679168, 
    -0.5275035, -0.5345182, -0.5846488, -0.7207162, -0.5985484, -0.1816375,
  0.5083363, 0.5225778, 0.9728868, 1.420413, 1.273457, 0.9397002, 0.871683, 
    0.8369987, 0.7452182, 0.6769727, 0.6643587, 0.6905631, 0.6811391, 
    0.4629099, 0.01606762, -0.388034, -0.4399869, -0.3880016, -0.4765755, 
    -0.4716114, -0.2407359, -0.06418946, -0.07125336, -0.037871, 0.02674484, 
    0.0113802, 0.01396775, 0.1380074, 0.2083042, 0.1648955, 0.09269524, 
    0.2324579, 0.3154331, 0.2590853, 0.3088086, 0.4884634, 0.4249217, 
    0.3492383, 0.5059928, 0.9544467, 0.8356315, 0.3378125, 0.01208007, 
    -0.07955402, -0.0630666, -0.1100225, -0.2707489, -0.3416307, -0.2699997, 
    -0.2155406, -0.1352997, 0.06020832, 0.3859081, 0.6496127, 0.7141471, 
    0.672708, 0.6928415, 0.7719595, 0.7616076, 0.5622752, 0.1264842, 
    -0.1615038, -0.1490042, -0.04605806, 0.01763022, 0.2164254, 0.5500846, 
    0.7850131, 0.8791701, 0.7711782, 0.4749544, 0.133125, -0.0109179, 
    -0.03508794, -0.0833627, -0.1546682, -0.09477222, 0.1328322, 0.4418004, 
    0.5823599, 0.4170118, 0.5535351, 0.470348, 0.7400746, 0.6790233, 
    0.4005075, 0.06579089, -0.1801405, -0.1959443, -0.03674841, 0.1007357, 
    0.2134147, 0.4077992, 0.4625683, 0.4503453, 0.5002472,
  0.8565464, 0.8466179, 1.316311, 1.374222, 1.175427, 0.9514843, 0.8022818, 
    0.6648308, 0.5314813, 0.5158235, 0.4875194, 0.3045604, 0.128291, 
    -0.03933591, -0.2838022, -0.4768687, -0.6245738, -0.7404592, -0.7145151, 
    -0.5402802, -0.3213347, -0.2098113, -0.1604137, -0.06454766, 0.002867818, 
    0.08751965, 0.1464715, 0.1919954, 0.118444, -0.05129886, 0.06175447, 
    0.3568715, 0.405765, 0.2317904, 0.2171582, 0.4417186, 0.5107778, 
    0.4875844, 0.636917, 0.8346715, 0.5092317, 0.02565438, -0.0310514, 
    0.1678906, 0.4129915, 0.4637239, 0.4345084, 0.423099, 0.458597, 
    0.5642937, 0.6996453, 0.9060255, 0.9861035, 0.85653, 0.5481316, 
    0.3971224, 0.3930535, 0.4998566, 0.4500358, 0.2028841, 0.02926761, 
    -0.03695965, 0.156709, 0.4078972, 0.5171256, 0.5692739, 0.7495313, 
    0.7967807, 0.6982455, 0.4980013, 0.2581901, 0.05910155, -0.05266604, 
    -0.1683724, -0.2285938, -0.05035496, 0.3307649, 0.787129, 1.010713, 
    1.140921, 1.293591, 1.25627, 1.357686, 1.203405, 0.9199087, 0.6419953, 
    0.4718133, 0.4133983, 0.5181184, 0.6480174, 0.701061, 0.8564157, 
    1.084752, 1.09888, 1.040318, 0.872529,
  1.165807, 1.310176, 1.205228, 1.099971, 0.7939161, 0.6915723, 0.5109246, 
    0.3451691, 0.129707, 0.03890306, -0.009957612, -0.1012175, -0.2340626, 
    -0.4391569, -0.6401498, -0.7834767, -0.8155568, -0.8021616, -0.733558, 
    -0.5921192, -0.4799448, -0.4562956, -0.4866667, -0.4197071, -0.2984833, 
    -0.1579396, -0.05068052, 0.03898442, 0.03369474, 0.0003614426, 0.1498567, 
    0.3810906, 0.3809441, 0.355586, 0.3816276, 0.458483, 0.4076201, 
    0.1977895, 0.02319646, -0.2169406, -0.5351205, -0.5358363, -0.4855925, 
    -0.1287404, 0.1519563, 0.2836618, 0.3856152, 0.5093457, 0.6820507, 
    0.9414909, 1.258304, 1.478486, 1.416344, 1.09486, 1.028243, 0.8000364, 
    0.8080766, 0.6968946, 0.409427, 0.1748077, 0.1043001, 0.364782, 
    0.6631217, 0.6894724, 0.4655306, 0.3820834, 0.4803093, 0.5365105, 
    0.4016145, 0.08509439, -0.2464812, -0.5451628, -0.4366667, -0.545472, 
    -0.3964649, 0.00566709, 0.6990104, 1.269958, 1.618851, 1.746455, 
    1.460859, 1.459248, 1.100882, 0.8170278, 0.7128125, 0.6605664, 0.6242057, 
    0.7637727, 1.013122, 1.260094, 1.452526, 1.563659, 1.602005, 1.477445, 
    1.205293, 1.270739,
  1.106807, 0.866198, 0.700703, 0.4284375, 0.1583528, 0.06032225, 
    -0.01124352, 0.02830738, -0.01396161, -0.09513022, -0.1817839, 
    -0.2558399, -0.3931283, -0.5354297, -0.6887338, -0.7599089, -0.7256966, 
    -0.6821257, -0.6222135, -0.573711, -0.4978646, -0.4251107, -0.3465462, 
    -0.2371061, -0.1387175, -0.08982423, -0.06619142, -0.09788087, 
    -0.1520638, -0.1405403, -0.05367523, 0.08854496, 0.276989, 0.3994987, 
    0.3791862, 0.1797721, -0.07504553, -0.2696419, -0.3970996, -0.4448048, 
    -0.4221649, -0.3506151, -0.1917285, 0.02018535, 0.1799345, 0.3482782, 
    0.612373, 0.7336463, 0.9363809, 1.122139, 1.218411, 1.191263, 1.39473, 
    1.104333, 0.7693883, 0.3922881, 0.2473012, 0.1564811, 0.1402539, 
    0.1875846, 0.3237175, 0.4888541, 0.5824413, 0.5406771, 0.4522982, 
    0.4345573, 0.4358919, 0.4203157, 0.1848991, -0.1388477, -0.3925098, 
    -0.3119597, -0.3213997, -0.2061166, 0.08097655, 0.4002311, 1.116263, 
    1.391556, 1.071601, 0.8307811, 0.4263378, 0.06401694, -0.1599412, 
    -0.1637826, 0.0349319, 0.3909705, 0.5644729, 0.7312696, 0.9593779, 
    1.189131, 1.36042, 1.516279, 1.621113, 1.609102, 1.485859, 1.280521,
  0.6529492, 0.4721712, 0.2794466, 0.08861001, -0.1594694, -0.3012012, 
    -0.2246224, -0.4090625, -0.423304, -0.4568326, -0.4893521, -0.5453255, 
    -0.6058073, -0.6795215, -0.7447397, -0.7261849, -0.6302702, -0.554554, 
    -0.5195606, -0.4945768, -0.4274056, -0.2850716, -0.1450163, -0.07288087, 
    -0.1201628, -0.2181934, -0.281849, -0.3029427, -0.2366016, -0.07239259, 
    0.04238605, 0.1150586, 0.119095, 0.03774738, -0.08694333, -0.2331022, 
    -0.2830209, -0.2107389, -0.08873373, -0.004440129, 0.08032551, 0.1218131, 
    0.2261751, 0.3236524, 0.4477896, 0.5693878, 0.8374219, 0.980114, 
    0.8327509, 0.9810419, 0.968428, 0.370039, 0.7393585, 0.5298859, 
    0.3165886, 0.1367709, 0.03587565, 0.06811848, 0.20347, 0.3792838, 
    0.4786816, 0.4719922, 0.4028841, 0.3255892, 0.2370638, 0.1865104, 
    0.09263021, -0.09434903, -0.2398404, -0.2224577, -0.005514354, 0.3412631, 
    0.7309115, 1.061706, 0.9121126, 0.9634798, 0.8609896, 1.206237, 
    0.8785189, 0.5034048, -0.08095372, -0.3399221, -0.2665169, -0.1949673, 
    -0.1465628, -0.01682591, 0.1903355, 0.4882848, 0.674206, 0.7506871, 
    0.7155797, 0.8239291, 0.7601756, 0.8338408, 0.872171, 0.8236848,
  0.4371775, 0.3655142, 0.2668815, 0.1641146, 0.03052086, -0.1342741, 
    -0.2317839, -0.3553353, -0.4793098, -0.606735, -0.675306, -0.6196256, 
    -0.6060026, -0.5602669, -0.6688932, -0.5325976, -0.3631803, -0.2118783, 
    -0.1044889, -0.03180014, 0.04788736, 0.1204134, 0.1654329, 0.1671745, 
    0.05737633, -0.1327278, -0.1145638, -0.001103461, 0.04752934, 0.07313156, 
    0.01502609, -0.09911776, -0.2341927, -0.3227018, -0.3410611, -0.3556281, 
    -0.1829718, -0.01637053, 0.106025, 0.2030791, 0.2345084, 0.2693063, 
    0.3640003, 0.486087, 0.5678741, 0.6110056, 0.58555, 0.461087, 0.3304393, 
    0.2662305, 0.2104851, 0.1757682, 0.117386, 0.432637, 0.4207392, 
    0.3439326, 0.26112, 0.1953319, 0.2421418, 0.3551952, 0.3943392, 
    0.2779977, 0.1386913, -0.02581048, -0.1543912, -0.2325488, -0.3067838, 
    -0.3281542, -0.2198535, 0.01196613, 0.3353873, 0.6063184, 0.7656119, 
    0.6207389, 0.7431022, 0.3883333, 0.5973666, 0.4982943, 0.4158398, 
    0.1874544, 0.05687177, -0.1336393, -0.1173795, -0.1329719, -0.1290169, 
    -0.1101855, -0.05391929, 0.04163736, 0.162308, 0.2448762, 0.3003775, 
    0.2688509, 0.3124055, 0.3687532, 0.3967154, 0.4404002,
  0.06144524, 0.05399072, 0.04337883, 0.0274446, 0.01019204, -0.04841805, 
    -0.1281868, -0.2219694, -0.2973274, -0.3408333, -0.3538704, -0.3519824, 
    -0.2858691, -0.167819, -0.1007129, -0.0542936, 0.05122393, 0.1070345, 
    0.1524609, 0.2127474, 0.3469758, 0.4468619, 0.478893, 0.412324, 
    0.2940136, 0.1743845, 0.1159211, 0.08909833, 0.1208527, 0.1736519, 
    0.1497265, 0.1281279, 0.08485043, 0.05765319, 0.05918264, 0.08139968, 
    0.1124218, 0.0988636, 0.1731312, 0.2156444, 0.2307165, 0.2393262, 
    0.2447788, 0.2574253, 0.2506542, 0.2399446, 0.201175, 0.1223173, 
    0.04214168, -0.02146506, -0.00517261, 0.1028352, 0.243786, 0.377705, 
    0.4381866, 0.4091501, 0.3338573, 0.2686558, 0.2531608, 0.2500517, 
    0.2212921, 0.110078, -0.02665687, 0.01769495, -0.02502936, -0.06311518, 
    -0.0630013, -0.04174481, -0.022181, -0.02893556, 0.08927733, 0.1141471, 
    0.083597, 0.04909179, 0.03758463, 0.04988931, 0.1106315, 0.214196, 
    0.2752308, 0.2460644, 0.1348338, -0.06251311, -0.1360156, -0.1269336, 
    -0.1175749, -0.1004037, -0.03752929, 0.01520506, 0.02420574, 0.06221028, 
    0.05319335, 0.07327797, 0.08657551, 0.01792315, 0.06094077, 0.08242512,
  -0.1120247, -0.1346158, -0.1593066, -0.1932585, -0.2504524, -0.2534146, 
    -0.2919563, -0.2785611, -0.2406706, -0.1889779, -0.04875977, 0.0861686, 
    0.2024935, 0.3001335, 0.337487, 0.3550488, 0.3666211, 0.3597201, 
    0.3591341, 0.3647004, 0.3771842, 0.4199739, 0.4445994, 0.4330759, 
    0.4128773, 0.2630405, 0.2668328, 0.3912308, 0.4376335, 0.5097203, 
    0.5284867, 0.4108433, 0.3703809, 0.3226273, 0.2740922, 0.2556188, 
    0.2468457, 0.2387726, 0.2616729, 0.2793652, 0.3039743, 0.3023797, 
    0.2443551, 0.2074251, 0.1547395, 0.09899402, 0.07121086, 0.0624218, 
    0.0519076, 0.07418936, 0.1149609, 0.1624382, 0.1952018, 0.2206901, 
    0.2143261, 0.1834018, 0.1451693, 0.1362663, 0.1439811, 0.1638216, 
    0.2092643, 0.239554, 0.2362825, 0.2267448, 0.1897168, 0.2549187, 
    0.2965854, 0.3235547, 0.3195508, 0.3329459, 0.3360384, 0.3527051, 
    0.3372591, 0.3162467, 0.3004915, 0.2894238, 0.2589063, 0.2137402, 
    0.04108357, -0.01824236, -0.07037431, -0.0582324, -0.01707033, 
    0.02057615, 0.04324874, 0.05241215, 0.05714852, 0.04341149, -0.01060873, 
    -0.03905925, -0.08018881, -0.212627, -0.1476855, -0.1136361, -0.09444663, 
    -0.1646777,
  0.02010415, 0.04069334, 0.02807942, 0.02710285, 0.09376952, 0.1168815, 
    0.15347, 0.1098502, 0.1691927, 0.2036979, 0.2549186, 0.2995801, 
    0.3510937, 0.3761263, 0.4022005, 0.4232617, 0.433239, 0.4373568, 
    0.4440299, 0.4475619, 0.4385124, 0.4375357, 0.4598014, 0.4577341, 
    0.4642446, 0.5474153, 0.5587597, 0.547236, 0.5579619, 0.5476754, 
    0.5250683, 0.5383333, 0.5163443, 0.4752636, 0.4470732, 0.4230498, 
    0.403535, 0.3882842, 0.3718293, 0.3440787, 0.3089061, 0.2541863, 
    0.1862826, 0.1260287, 0.06585616, 0.008776069, -0.02086258, -0.03134441, 
    -0.02369469, -0.009567052, 0.02028319, 0.07329426, 0.1126497, 0.1438346, 
    0.1576205, 0.1579949, 0.1601595, 0.1598015, 0.1550489, 0.1714063, 
    0.1918165, 0.2059441, 0.2250358, 0.263545, 0.2894727, 0.3064324, 
    0.3065951, 0.3022169, 0.2948764, 0.293916, 0.2910677, 0.3067253, 
    0.2729687, 0.1791862, 0.1250032, 0.07265949, 0.01710933, -0.02493167, 
    -0.05444014, -0.0694629, -0.06798179, -0.05753256, -0.05219403, 
    -0.04415366, -0.02113932, -0.009599626, -0.003300816, -0.01516601, 
    -0.04830405, -0.08105145, -0.1149544, -0.1195931, -0.09303061, 
    -0.07472007, -0.0464974, -0.01850262,
  0.08279948, 0.1274772, 0.1710807, 0.1885286, 0.2001172, 0.2143262, 
    0.2230338, 0.2131868, 0.2103711, 0.2030957, 0.1865104, 0.1810091, 
    0.1830762, 0.1853223, 0.1893424, 0.1976107, 0.2199414, 0.242207, 
    0.2780469, 0.3276726, 0.3710482, 0.4209995, 0.4621776, 0.4962923, 
    0.5223826, 0.5323924, 0.5379425, 0.5339061, 0.5339549, 0.5288604, 
    0.517272, 0.5045116, 0.4850128, 0.4600129, 0.4293001, 0.3947948, 
    0.3631381, 0.3293165, 0.2876824, 0.2547233, 0.2294303, 0.2006217, 
    0.1806836, 0.1616243, 0.1454297, 0.1371777, 0.1248568, 0.1287955, 
    0.1375684, 0.142793, 0.1560742, 0.1590365, 0.159834, 0.154235, 0.1444695, 
    0.126875, 0.1130078, 0.1086622, 0.1037956, 0.1055697, 0.1079786, 
    0.1254265, 0.1391635, 0.1409213, 0.147334, 0.1553743, 0.1488314, 
    0.1444531, 0.1355664, 0.1243196, 0.09468099, 0.07575193, 0.06024089, 
    0.03115559, 0.01969725, -0.021709, -0.05751628, -0.1019824, -0.143763, 
    -0.1666634, -0.1889616, -0.2393522, -0.2296192, -0.2537728, -0.2541797, 
    -0.2677214, -0.2742806, -0.2603646, -0.2488249, -0.2327116, -0.1933236, 
    -0.1524056, -0.1086882, -0.05969727, -0.01163414, 0.03099284,
  -0.2447233, -0.2378548, -0.2318002, -0.2266732, -0.2219206, -0.219821, 
    -0.2200814, -0.2167448, -0.2074512, -0.1997689, -0.2013477, -0.1967741, 
    -0.1832487, -0.1708138, -0.1533334, -0.1331348, -0.110918, -0.08263022, 
    -0.05191734, -0.01991865, 0.01610026, 0.05277017, 0.08747071, 0.1254915, 
    0.1608756, 0.19403, 0.2251823, 0.2543164, 0.2794629, 0.301875, 0.3244499, 
    0.3462435, 0.3668164, 0.3839551, 0.3974805, 0.4074251, 0.418737, 
    0.4324414, 0.4422884, 0.4474967, 0.4535026, 0.4560742, 0.4575879, 
    0.446569, 0.4385775, 0.4308463, 0.4106315, 0.3883333, 0.3645377, 
    0.3377962, 0.3093457, 0.2804557, 0.2467643, 0.2090853, 0.1663444, 
    0.1366081, 0.1034375, 0.06826496, 0.03574544, 0.007392555, -0.01835611, 
    -0.04672527, -0.06147137, -0.07724285, -0.0860482, -0.0958301, 
    -0.1098926, -0.1187468, -0.1272754, -0.1350553, -0.1477832, -0.1613249, 
    -0.174541, -0.1883268, -0.2005339, -0.2156218, -0.2302051, -0.2432096, 
    -0.2564421, -0.2716602, -0.2869759, -0.2994922, -0.3083138, -0.3134245, 
    -0.3140267, -0.3187305, -0.3223275, -0.3283008, -0.328903, -0.3211719, 
    -0.3115365, -0.3003711, -0.2899544, -0.2780404, -0.2634082, -0.2530241,
  -0.217917, -0.2344537, -0.2509246, -0.2669082, -0.2826797, -0.2985487, 
    -0.3143038, -0.3304333, -0.346807, -0.3633271, -0.3798148, -0.3968071, 
    -0.4138649, -0.43154, -0.4498668, -0.4688773, -0.4884086, -0.5086071, 
    -0.5291963, -0.5489717, -0.56847, -0.5873013, -0.6035938, -0.6168427, 
    -0.6256638, -0.6298628, -0.6291142, -0.6230111, -0.6110811, -0.5925426, 
    -0.5679336, -0.5380669, -0.5032196, -0.4635551, -0.4182587, -0.3694468, 
    -0.3168914, -0.2614229, -0.2034966, -0.1440728, -0.08386743, -0.02387409, 
    0.03486615, 0.09186471, 0.1462756, 0.1986518, 0.2600291, 0.293134, 
    0.3300159, 0.3779492, 0.3887239, 0.4178581, 0.48874, 0.4590364, 
    0.4841018, 0.4909539, 0.4943724, 0.4853878, 0.5329623, 0.5492225, 
    0.5578651, 0.5260453, 0.5503941, 0.5529332, 0.5610061, 0.5678906, 
    0.5748572, 0.58498, 0.5860219, 0.5821486, 0.563952, 0.5545115, 0.5654979, 
    0.4022653, 0.4066434, 0.4125361, 0.3765497, 0.2689815, 0.3389845, 
    0.2825556, 0.2408566, 0.2005572, 0.1648803, 0.1235228, 0.08571386, 
    0.05145264, 0.01990986, -0.01028252, -0.03944874, -0.06690645, 
    -0.09263945, -0.1168098, -0.1417603, -0.1627083, -0.1817021, -0.2002902,
  0.1301786, 0.1155465, 0.09593379, 0.07791626, 0.06251913, 0.0517444, 
    0.04292279, 0.03188764, 0.01662068, -0.0008923411, -0.01856813, -0.03849, 
    -0.06220406, -0.09049195, -0.1202121, -0.1474907, -0.1709445, -0.189597, 
    -0.2089169, -0.2227674, -0.24417, -0.2742646, -0.3169727, -0.3754363, 
    -0.4486785, -0.528089, -0.6052537, -0.6752081, -0.7313113, -0.7694459, 
    -0.7887497, -0.790637, -0.7779751, -0.7493954, -0.7035446, -0.6392536, 
    -0.5569625, -0.4601688, -0.3528781, -0.2440727, -0.1251271, -0.05419636, 
    -0.008802533, 0.03177387, 0.03045535, -0.008444786, -0.03053069, 
    -0.07828522, -0.1188447, -0.1507461, -0.2022755, -0.2843881, -0.1425588, 
    -0.2125945, 0.02371716, -0.2774053, -0.201673, -0.1571417, -0.07585907, 
    0.007279396, 0.07890987, 0.1615267, 0.2485542, 0.3259144, 0.4025581, 
    0.4621124, 0.5165066, 0.5636421, 0.5705432, 0.5679391, 0.5618681, 
    0.5299996, 0.4843777, 0.474124, 0.3956572, 0.4092477, 0.3740263, 
    0.3345243, 0.2526232, 0.1886253, 0.1582549, 0.1948924, 0.08170891, 
    0.1060414, 0.06951857, 0.05091524, 0.07062531, 0.07977247, 0.08662462, 
    0.09326506, 0.1010942, 0.1109567, 0.127363, 0.1337759, 0.13638, 0.1350611,
  0.1309272, 0.1352406, 0.1344104, 0.1540231, 0.1796578, 0.2023792, 
    0.2221057, 0.2456572, 0.2770048, 0.3140816, 0.3417997, 0.3574411, 
    0.3558296, 0.3361676, 0.2970896, 0.2393095, 0.1613145, 0.07186222, 
    -0.0118289, -0.08894539, -0.1570606, -0.2221487, -0.2738905, -0.2806123, 
    -0.2673149, -0.2776013, -0.3282686, -0.4043597, -0.4923797, -0.5964975, 
    -0.7159474, -0.8500781, -0.9765105, -1.074801, -1.138278, -1.174575, 
    -1.167739, -1.110058, -0.9856272, -0.7942686, -0.5491524, -0.3089156, 
    0.05127335, 0.2025905, 0.1968938, 0.1551948, 0.07928342, -0.014906, 
    -0.1173311, -0.2276827, -0.3366833, -0.4207003, -0.4704887, -0.4795381, 
    -0.4442842, -0.3878716, -0.3239719, -0.2549614, -0.170505, -0.0943656, 
    -0.01477587, 0.06455362, 0.1450061, 0.2209827, 0.2802112, 0.3212106, 
    0.3506539, 0.3804228, 0.4079292, 0.4209175, 0.4175644, 0.4001817, 
    0.3739934, 0.3300159, 0.3209664, 0.3111845, 0.3022165, 0.2578316, 
    0.2789254, 0.2754423, 0.2580595, 0.2179227, 0.2209661, 0.2005403, 
    0.279788, 0.3146839, 0.3118684, 0.3027377, 0.2768745, 0.2619987, 
    0.2339878, 0.2188349, 0.1811557, 0.1675649, 0.1600616, 0.1522164,
  0.3524451, 0.3407745, 0.3191435, 0.28791, 0.266572, 0.252054, 0.2573918, 
    0.2690618, 0.2872099, 0.317288, 0.3462268, 0.3554716, 0.3429879, 
    0.3226916, 0.2921741, 0.252135, 0.2308459, 0.2336457, 0.2569366, 
    0.3140984, 0.3783245, 0.4240928, 0.3807817, 0.2511909, 0.1175158, 
    0.1024605, 0.06471652, -0.04037809, -0.1589652, -0.2415824, -0.2989229, 
    -0.352048, -0.4114718, -0.5039848, -0.6639621, -0.9077606, -1.165964, 
    -1.386585, -1.515818, -1.505402, -1.337156, -1.055076, -0.596612, 
    -0.08616209, 0.2053905, 0.3368351, 0.2013535, 0.1445177, 0.03844702, 
    -0.0628714, -0.1763318, -0.2401175, -0.292038, -0.3109347, -0.3261364, 
    -0.3201957, -0.2430799, -0.2893364, -0.2776501, -0.2543914, -0.2540498, 
    -0.2390599, -0.2265432, -0.1670868, -0.140264, -0.07857752, -0.03508806, 
    -0.007825851, 0.006790161, 0.04415989, 0.08789372, 0.1268744, 0.1471221, 
    0.1432648, 0.1636255, 0.1395208, 0.09186482, 0.0462268, 0.03340131, 
    0.0145862, 0.06325155, 0.0776884, 0.1258492, 0.1633168, 0.2071644, 
    0.2608916, 0.3125679, 0.3406768, 0.3404648, 0.4473014, 0.4434114, 
    0.3581743, 0.3981476, 0.3628778, 0.3371611, 0.3206735,
  0.06644249, 0.1049681, 0.09435558, 0.1066284, 0.03493261, 0.03139973, 
    0.0224967, 0.03325558, -0.05606747, 0.1060424, 0.1876163, 0.2556019, 
    0.2986693, 0.2911487, 0.2612659, 0.2643421, 0.2656281, 0.237112, 
    0.1854358, 0.1430852, 0.2723179, 0.4284525, 0.499774, 0.5147333, 
    0.4643593, 0.4104691, 0.415628, 0.3910189, 0.3193064, 0.232523, 
    0.1630888, 0.1286001, 0.1100452, 0.07241511, -0.03128004, -0.2337542, 
    -0.4917618, -0.7186332, -0.9547823, -1.211944, -1.348825, -1.278562, 
    -1.006426, -0.6262991, -0.2544239, 0.03839779, 0.1097522, 0.1669787, 
    0.1624213, 0.1327339, 0.01504183, -0.09731162, -0.2198865, -0.2937145, 
    -0.3157686, -0.3098279, -0.3158988, -0.3227673, -0.3192191, -0.3812797, 
    -0.4731092, -0.5752413, -0.6273408, -0.6395155, -0.591322, -0.5363902, 
    -0.4645153, -0.4111137, -0.3303519, -0.2020968, -0.2062311, -0.2277316, 
    -0.1478651, -0.1166149, -0.09324265, -0.1428682, -0.2681449, -0.3606254, 
    -0.3959769, -0.4198702, -0.4178357, -0.32835, -0.2909314, -0.2568168, 
    -0.1752738, -0.06653357, 0.05625284, 0.2008981, 0.3340523, 0.4624867, 
    0.5316112, 0.5758982, 0.5621777, 0.4539094, 0.3346553, 0.1386919,
  0.03875637, 0.03672218, -0.2492485, -0.3739066, -0.4856415, -0.451592, 
    -0.4014459, -0.3436329, -0.2781544, -0.2235489, -0.1824028, -0.05411434, 
    0.01789093, 0.07536173, 0.04692745, 0.02353811, 0.1519233, 0.1532418, 
    0.1648793, 0.1202339, 0.1352732, 0.2200227, 0.354073, 0.3930368, 
    0.3608255, 0.2906933, 0.250246, 0.2811699, 0.3694677, 0.5135117, 
    0.6444693, 0.8239288, 0.9374208, 0.9236689, 0.8670607, 0.7663288, 
    0.6332064, 0.4458528, 0.2463574, 0.05335569, -0.09324217, -0.1964819, 
    -0.1556935, -0.06047893, 0.04022098, 0.1376656, 0.1809924, 0.1999703, 
    0.2409372, 0.2693062, 0.2479845, 0.1969429, 0.1306828, 0.09184813, 
    0.1034043, 0.1948917, 0.2941756, 0.3419464, 0.3301463, 0.2511263, 
    0.140449, 0.02794886, -0.08419275, -0.2320125, -0.3901663, -0.5120738, 
    -0.5918915, -0.623174, -0.6386039, -0.6543432, -0.6647111, -0.5949683, 
    -0.478464, -0.3315076, -0.1781384, -0.08048224, -0.07131889, -0.07079792, 
    -0.1360486, -0.1994438, -0.2827772, -0.219268, -0.1716118, -0.1422335, 
    -0.1497205, -0.1681938, -0.161195, -0.09941131, 0.01419558, 0.1419137, 
    0.3038278, 0.4409208, 0.5471543, 0.5680368, 0.4637401, 0.2743683,
  0.6614612, 0.5059599, 0.310208, 0.1249377, -0.0116508, -0.1040339, 
    -0.1640437, -0.2304983, -0.3089978, -0.3790662, -0.3642712, -0.3331839, 
    -0.3225396, -0.3247044, -0.4104466, -0.4676242, -0.4962213, -0.4478813, 
    -0.3606091, -0.2296358, -0.1004691, 0.03012976, 0.1480497, 0.2160022, 
    0.2590845, 0.1829615, 0.06657159, 0.06028903, 0.1300156, 0.250133, 
    0.4312036, 0.6408231, 0.9524121, 1.25601, 1.316165, 1.391312, 1.147611, 
    1.032116, 0.9242055, 0.8086782, 0.7209177, 0.6869655, 0.6419301, 
    0.5793159, 0.4885935, 0.4115914, 0.3161324, 0.2713895, 0.2619817, 
    0.3153346, 0.3990586, 0.5021183, 0.5994008, 0.6464875, 0.6706574, 
    0.7301626, 0.9232454, 1.032506, 1.079463, 1.105618, 1.075475, 1.05002, 
    1.103307, 1.072366, 1.039131, 0.9040389, 0.8690298, 0.7343616, 0.715205, 
    0.5367057, 0.4050159, 0.3952017, 0.3604848, 0.3406606, 0.2782094, 
    0.1403835, -0.01853585, -0.07224691, -0.1124487, -0.1041968, -0.1381974, 
    -0.1907847, -0.1671357, -0.09565187, -0.01570368, 0.08491445, 0.1423531, 
    0.1363144, 0.09748018, 0.09866822, 0.1684924, 0.3299508, 0.4827015, 
    0.6080594, 0.714456, 0.7321481,
  0.6528509, 0.6132188, 0.6012397, 0.6034532, 0.502558, 0.4803574, 0.5074244, 
    0.5661163, 0.5535023, 0.5026236, 0.6150908, 0.7335317, 0.8132517, 
    0.7203965, 0.532213, 0.3022976, 0.06178641, -0.05896568, -0.1344044, 
    -0.2133434, -0.2325327, -0.1832325, -0.0591929, 0.1112173, 0.2978702, 
    0.4314315, 0.4333849, 0.3526721, 0.3124703, 0.3712106, 0.5988797, 
    0.7628121, 0.9411325, 1.249661, 1.425426, 1.449905, 1.464586, 1.515009, 
    1.368004, 1.195966, 1.088121, 1.121308, 1.165302, 1.201924, 1.149873, 
    0.9858916, 0.691751, 0.4333687, 0.3238635, 0.3809276, 0.4094758, 
    0.4831414, 0.535892, 0.6067572, 0.9124861, 1.109395, 1.383614, 1.800736, 
    2.148408, 2.350785, 2.202201, 2.140221, 2.031253, 1.935176, 1.769795, 
    1.570511, 1.324287, 1.116557, 0.9185743, 0.7598181, 0.6485224, 0.5693069, 
    0.448441, 0.2730832, 0.140873, 0.08493185, 0.1834183, 0.3636265, 
    0.6535354, 0.9544635, 1.121683, 0.7556834, 0.325182, 0.1746938, 
    0.1748891, 0.245348, 0.3406608, 0.4029164, 0.4288278, 0.4700062, 
    0.5090201, 0.5093131, 0.5170765, 0.5769231, 0.6590357, 0.6971867,
  0.9471223, 0.8531117, 0.8904333, 1.03612, 1.080586, 1.007344, 1.066524, 
    0.9939165, 0.8214231, 0.7355666, 0.7504272, 0.7659059, 0.8779988, 
    0.9218626, 1.058208, 1.12795, 1.231303, 1.377999, 1.589946, 1.729122, 
    1.486853, 1.41628, 1.526436, 1.594502, 1.621472, 1.686332, 1.694421, 
    1.591296, 1.352689, 1.153715, 0.9187531, 0.7594762, 0.7507687, 0.7360554, 
    0.711885, 0.7603059, 0.9106321, 1.144926, 1.328291, 1.420772, 1.415807, 
    1.436755, 1.494144, 1.555961, 1.54683, 1.447953, 1.25295, 1.009753, 
    0.8751502, 0.9324903, 1.009834, 0.9621615, 0.9596062, 1.121943, 1.312373, 
    1.474156, 1.665465, 1.893964, 2.15163, 2.333613, 2.316833, 2.153731, 
    2.072969, 2.126223, 2.11151, 2.021308, 1.913285, 1.818574, 1.663203, 
    1.493981, 1.371781, 1.28477, 1.108874, 0.9092975, 0.8558459, 0.8935905, 
    0.8311067, 0.7303581, 0.7228551, 0.8362832, 0.9820518, 1.091117, 
    1.460941, 1.704935, 1.616817, 1.654073, 1.807963, 1.976387, 1.779366, 
    1.744242, 1.712113, 1.445153, 1.154675, 1.034362, 1.042516, 1.084329,
  0.9498415, 0.8196983, 0.7662964, 0.7822795, 0.8005571, 0.8430381, 
    0.8573122, 0.7391644, 0.5633502, 0.3723993, 0.1665239, -0.04916668, 
    -0.20086, -0.2404766, -0.2067842, -0.07527447, 0.1565113, 0.3780451, 
    0.4651375, 0.5035334, 0.6576996, 0.6612158, 0.7221527, 0.8660326, 
    1.004542, 1.136347, 1.24826, 1.311052, 1.310143, 1.232264, 1.091265, 
    0.9735718, 0.9815793, 1.005961, 0.914392, 0.7290893, 0.5898967, 
    0.6106157, 0.7368526, 0.8637085, 0.9447794, 1.027966, 1.144584, 1.222595, 
    1.238904, 1.265499, 1.236608, 1.01335, 0.744307, 0.7062535, 0.7690792, 
    0.7089229, 0.5846553, 0.6702018, 0.8994331, 1.098017, 1.306595, 1.579235, 
    1.90002, 2.238268, 2.408044, 2.333076, 2.21265, 2.293216, 2.374238, 
    2.331058, 2.28879, 2.302819, 2.209281, 2.071308, 1.993948, 1.84639, 
    1.504902, 1.185078, 1.133223, 1.160778, 0.9673696, 0.6574254, 0.6498733, 
    0.9097538, 1.180001, 1.393428, 1.532458, 1.45448, 1.246439, 1.150867, 
    1.133402, 1.132572, 1.172578, 1.234102, 1.191882, 1.126794, 1.036625, 
    0.9914265, 1.01864, 1.064538,
  1.187292, 1.26016, 1.317517, 1.255522, 1.070431, 0.9083538, 0.7639036, 
    0.5979047, 0.4121623, 0.2672567, 0.1477566, 0.01128101, -0.06028461, 
    -0.03897858, 0.01609898, 0.1252289, 0.322917, 0.5120783, 0.5617847, 
    0.5326509, 0.4874201, 0.3792334, 0.2539244, 0.2719898, 0.4475117, 
    0.6581879, 0.8113785, 0.8818531, 0.9118176, 0.9169445, 0.8532896, 
    0.736248, 0.7113609, 0.8209333, 0.9119816, 0.8710155, 0.7324753, 
    0.621911, 0.6160841, 0.718884, 0.8660684, 0.9208698, 0.927299, 1.002755, 
    1.059216, 1.042126, 1.043949, 0.929821, 0.5947785, 0.3548536, 0.3832879, 
    0.2716022, -0.03035164, -0.1239223, 0.0009961128, 0.196568, 0.4681504, 
    0.7840357, 1.149124, 1.584524, 1.979642, 2.030423, 1.941116, 1.964423, 
    2.016914, 2.011901, 2.03013, 2.078893, 2.084297, 2.105179, 2.17191, 
    2.15111, 1.925735, 1.666881, 1.515335, 1.337747, 0.9144232, 0.6861854, 
    0.8105187, 0.8822794, 0.7397504, 0.7440639, 0.9286003, 0.9380088, 
    0.8681526, 0.8770065, 0.8863811, 0.829155, 0.8238316, 0.8839884, 
    0.9615431, 1.05894, 1.137537, 1.11838, 1.082979, 1.12043,
  1.186365, 1.14242, 1.14185, 1.060063, 0.9404497, 0.8749228, 0.8428917, 
    0.7714233, 0.6734738, 0.6183796, 0.6022177, 0.5647016, 0.5198612, 
    0.4931359, 0.4855185, 0.4472694, 0.4312191, 0.4793005, 0.5377464, 
    0.5838394, 0.6910334, 0.6724949, 0.4601898, 0.2956228, 0.3022795, 
    0.3780613, 0.4598484, 0.5076342, 0.4936047, 0.4600601, 0.4442234, 
    0.4274912, 0.3794451, 0.3606129, 0.4434748, 0.5456886, 0.5248556, 
    0.4653015, 0.4425802, 0.5066118, 0.6722364, 0.6958051, 0.5535522, 
    0.622921, 0.7897334, 0.6858759, 0.6332717, 0.8213248, 0.8314977, 
    0.6270049, 0.6043489, 0.5056016, 0.08283138, -0.2416475, -0.3281546, 
    -0.4474092, -0.4725556, -0.2457325, 0.04015565, 0.3494818, 0.6834662, 
    0.883466, 0.9973984, 1.089846, 1.145251, 1.228909, 1.427689, 1.648164, 
    1.777021, 1.876761, 1.930212, 1.868509, 1.727835, 1.554104, 1.383776, 
    1.153258, 0.7145698, 0.5583527, 0.7101102, 0.6892781, 0.2813678, 
    0.01968145, 0.05138779, 0.122107, 0.2165403, 0.3727245, 0.5061884, 
    0.5200729, 0.4677286, 0.44102, 0.4924679, 0.7076864, 0.9322958, 1.041475, 
    1.112227, 1.197188,
  1.024336, 1.043396, 1.110746, 1.163611, 1.231986, 1.350411, 1.417891, 
    1.385128, 1.268493, 1.17349, 1.176973, 1.227869, 1.254692, 1.199597, 
    1.159819, 1.1363, 1.055359, 1.046912, 1.073702, 1.094095, 1.0932, 
    0.9903345, 0.7782402, 0.5741386, 0.4165697, 0.3144865, 0.2746429, 
    0.2798185, 0.257309, 0.1430998, 0.017416, 0.01217556, 0.05633259, 
    0.0976572, 0.2242699, 0.3386412, 0.2760925, 0.2014675, 0.2230501, 
    0.3101425, 0.5282764, 0.6267943, 0.4214392, 0.3902869, 0.5831256, 
    0.5463734, 0.3369823, 0.6016796, 0.9038768, 0.9916697, 1.019241, 
    0.9327993, 0.4984894, -0.02509451, -0.4421036, -0.8990531, -1.203089, 
    -1.185609, -1.054863, -0.8802216, -0.7290173, -0.6381154, -0.5429821, 
    -0.3285778, -0.1146948, 0.06681585, 0.3102238, 0.550019, 0.7069201, 
    0.9079289, 1.164147, 1.375003, 1.406367, 1.197382, 0.9460001, 0.7743521, 
    0.5474803, 0.2450876, 0.3404651, 0.3611522, 0.2555375, 0.1273961, 
    -0.0675745, -0.229033, -0.2967582, -0.3050742, -0.1564412, 0.02908945, 
    0.1132689, 0.142745, 0.1849651, 0.3399458, 0.5631876, 0.7019739, 
    0.8002644, 0.9377642,
  0.9060755, 0.9836793, 1.176274, 1.33031, 1.392436, 1.398441, 1.324369, 
    1.334688, 1.378177, 1.39185, 1.408824, 1.449693, 1.544534, 1.534655, 
    1.446341, 1.346243, 1.149727, 0.9316931, 0.8000522, 0.7864947, 0.7921753, 
    0.6264524, 0.3913774, 0.1257524, -0.1345015, -0.2770653, -0.4106255, 
    -0.5392075, -0.5316553, -0.5081367, -0.5107079, -0.4341278, -0.3818007, 
    -0.3402481, -0.1790333, -0.04512978, -0.07996082, -0.08987236, 
    -0.09040928, -0.06246424, 0.1624064, 0.317029, 0.1987181, 0.07607794, 
    0.2153192, 0.3901072, 0.3192902, 0.2478709, 0.5314808, 0.8015003, 
    0.8864613, 0.6988802, 0.2065296, -0.3022106, -0.7056608, -1.110609, 
    -1.460218, -1.665297, -1.78792, -1.734584, -1.544024, -1.47765, 
    -1.536683, -1.438571, -1.187041, -0.9615202, -0.774297, -0.574297, 
    -0.3468232, -0.08197927, 0.2081575, 0.4197135, 0.5654655, 0.4718132, 
    0.1773467, -0.02542019, -0.1886199, -0.2961562, -0.05688167, 
    -0.002747536, -0.08206081, -0.09791374, -0.2138476, -0.3426237, 
    -0.3769665, -0.4485159, -0.3326464, -0.1346321, 0.01461983, 0.128129, 
    0.1892457, 0.1943889, 0.2691612, 0.4513221, 0.5782428, 0.7531128,
  0.3867388, 0.3943391, 0.5150099, 0.6099648, 0.6444361, 0.7049999, 
    0.7057481, 0.7274771, 0.6997428, 0.7551301, 0.8551946, 0.8095405, 
    0.88511, 0.9762884, 0.9194363, 0.8155462, 0.6814643, 0.4703476, 
    0.1144562, -0.1706188, -0.3466446, -0.6051564, -0.827064, -0.9942679, 
    -1.161308, -1.205465, -1.226868, -1.214238, -1.067737, -1.101787, 
    -1.162382, -0.9518847, -0.8108525, -0.7562299, -0.6024218, -0.546351, 
    -0.4873176, -0.2438772, -0.1778779, -0.3072565, -0.2203422, 0.0152216, 
    0.06940413, -0.07304382, -0.1256804, -0.04374695, -0.09233093, 
    -0.2021291, -0.2199676, -0.1906545, -0.0793426, -0.06054378, -0.312269, 
    -0.7141733, -1.088067, -1.423695, -1.765736, -1.999606, -2.126804, 
    -2.187253, -1.998353, -1.717787, -1.604587, -1.630091, -1.636797, 
    -1.534746, -1.336227, -1.103643, -0.7936492, -0.4960585, -0.3296847, 
    -0.2963996, -0.2620249, -0.2178519, -0.3098772, -0.3275523, -0.1606905, 
    -0.0486787, -0.2067517, -0.02880585, -0.05320358, -0.2050591, -0.4287732, 
    -0.4775524, -0.3113582, -0.1116831, 0.08071613, 0.1998401, 0.2828326, 
    0.2553582, 0.184525, 0.1300983, 0.02192783, 0.09129572, 0.159802, 
    0.2404656,
  -0.2655411, -0.2781219, -0.1767066, -0.1259573, -0.06384805, 0.1285673, 
    0.2471384, 0.2064154, -0.06209028, -0.1943169, 0.03641237, -0.03477901, 
    -0.06184614, 0.1420764, 0.2143583, 0.08501256, -0.06077194, -0.1663384, 
    -0.4429171, -0.7769504, -0.9692842, -1.103204, -1.241713, -1.330433, 
    -1.424346, -1.500729, -1.529294, -1.529668, -1.42625, -1.39155, 
    -1.235169, -0.7432426, -0.5266081, -0.4484835, -0.3753712, -0.3611948, 
    -0.4093559, -0.3206841, -0.244805, -0.2990694, -0.3080211, -0.209877, 
    0.0303086, 0.0006375313, -0.2449516, -0.4991997, -0.8098933, -1.038132, 
    -1.265785, -1.360983, -1.098239, -0.8397917, -0.7826465, -0.9660776, 
    -1.295146, -1.561065, -1.833086, -2.058428, -2.151071, -2.253431, 
    -2.211195, -2.031394, -1.893405, -1.878219, -1.93416, -1.919593, 
    -1.842185, -1.768975, -1.650062, -1.484486, -1.212611, -0.9794898, 
    -0.9157685, -0.8027316, -0.7717419, -0.6524385, -0.1824027, -0.01300168, 
    -0.3152803, -0.1900362, -0.03015664, -0.1054984, -0.3348441, -0.5147107, 
    -0.3960584, -0.1702609, -0.07473683, -0.1262832, -0.06394601, 
    -0.06052804, -0.1052547, -0.01228571, -0.1252899, -0.1637828, -0.2237926, 
    -0.3367972,
  -0.6225069, -0.7127413, -0.6322725, -0.4613255, -0.08767629, 0.2508655, 
    0.3206573, 0.2738636, -0.08586955, -0.5334444, -0.5546361, -0.6046355, 
    -0.88989, -0.746628, -0.1824677, -0.09504914, -0.1956186, -0.2659311, 
    -0.4477673, -0.7056937, -0.8583956, -0.8105767, -0.8004529, -0.8467255, 
    -0.9627581, -1.127406, -1.126967, -1.162758, -1.247898, -1.212709, 
    -0.986423, -0.6835911, -0.5525523, -0.4480928, -0.4265759, -0.3128226, 
    -0.2044405, -0.2650199, -0.2665987, -0.2836234, -0.3516898, -0.6070772, 
    -0.6630179, -0.8218558, -1.090736, -1.261618, -1.461163, -1.627439, 
    -1.725974, -1.633347, -1.443308, -1.262448, -0.9881806, -0.8366019, 
    -0.8734998, -0.9749809, -1.054392, -1.183884, -1.34378, -1.535756, 
    -1.685593, -1.706866, -1.58574, -1.462823, -1.53958, -1.6082, -1.696123, 
    -1.856377, -1.862546, -1.738441, -1.505238, -1.189369, -1.029408, 
    -0.853057, -0.6163383, -0.5048149, -0.1030575, 0.2096872, -0.07496464, 
    -0.05958372, 0.07547486, -0.126283, -0.3188285, -0.4825981, -0.8239392, 
    -1.042494, -0.772686, -0.5694307, -0.681947, -0.5859834, -0.467266, 
    -0.3231091, -0.300225, -0.3156222, -0.3728162, -0.5171683,
  -0.4854786, -0.4319143, -0.362318, -0.1675267, 0.1611031, 0.1361681, 
    -0.0292294, -0.05567777, -0.1291639, -0.600111, -0.7919569, -0.3919404, 
    -0.8243296, -1.075908, -0.5218387, -0.4841599, -0.5776496, -0.6037879, 
    -0.5391078, -0.4899697, -0.5850878, -0.6874638, -0.7157192, -0.7122521, 
    -0.6966438, -0.6824508, -0.6785607, -0.6368456, -0.6119437, -0.6222625, 
    -0.471839, -0.3736954, -0.3432429, -0.3101697, -0.4285126, -0.3732879, 
    -0.1646296, -0.1611792, -0.2271459, -0.3208468, -0.5402156, -0.8020639, 
    -1.015817, -1.346238, -1.599102, -1.668813, -1.638116, -1.533119, 
    -1.549883, -1.512286, -1.43779, -1.281736, -1.009747, -0.7962865, 
    -0.6943984, -0.7835261, -0.7420546, -0.6723608, -0.6785131, -0.7553031, 
    -0.9147595, -1.021726, -1.051771, -1.039939, -1.156198, -1.237806, 
    -1.328952, -1.473354, -1.514044, -1.441697, -1.359128, -1.199379, 
    -1.037253, -0.8581188, -0.4863257, -0.1063448, 0.1725454, 0.2843941, 
    -0.1183238, -0.04706749, 0.1058623, -0.114548, -0.3174129, -0.3316379, 
    -0.6108857, -1.198598, -1.241403, -0.7363739, -0.7586565, -0.6657202, 
    -0.5844214, -0.5284312, -0.4267874, -0.415508, -0.3882294, -0.4221814,
  -0.107842, -0.0755825, -0.008623362, 0.2380559, 0.1792669, 0.08802342, 
    0.02064037, -0.1863251, -0.1094046, -0.2544403, -0.4298638, 0.08888626, 
    0.03032517, -0.2998996, -0.5273082, -0.7039027, -0.6465454, -0.6381955, 
    -0.5217409, -0.4115191, -0.38416, -0.4466763, -0.3868942, -0.2540483, 
    -0.2447872, -0.1549926, -0.2019, -0.2421184, -0.2454882, -0.2655239, 
    -0.2223434, -0.2203741, -0.2480922, -0.1298962, -0.2714815, -0.1416798, 
    0.03341722, -0.03253293, -0.1782196, -0.3846323, -0.6805954, -0.9300094, 
    -0.9761519, -1.199947, -1.318291, -1.406718, -1.478382, -1.417591, 
    -1.466452, -1.348906, -1.079261, -1.003203, -0.883038, -0.6351211, 
    -0.4456842, -0.4406221, -0.3952281, -0.3238251, -0.1075492, 0.06647444, 
    0.01761389, -0.1056285, -0.3636856, -0.5003712, -0.6437635, -0.897702, 
    -1.116712, -1.130662, -1.137709, -1.078414, -0.9157357, -0.879456, 
    -0.6596646, -0.2943006, -0.05539989, 0.268883, 0.421536, 0.1362007, 
    -0.1585258, -0.0394665, 0.09712195, -0.1726367, -0.4419076, -0.3470514, 
    -0.3352673, -0.6052383, -0.9309697, -0.7311649, -0.6009893, -0.475143, 
    -0.4115362, -0.3544722, -0.2973433, -0.2781539, -0.2245088, -0.1644988,
  0.214766, 0.1824088, 0.2174342, 0.1229197, -0.1842259, -0.2107885, 
    0.03239179, -0.03450227, -0.1443493, -0.1445611, -0.3475395, -0.2547497, 
    -0.1268041, -0.4044571, -0.6343393, -0.7584758, -0.6152306, -0.5920701, 
    -0.4104128, -0.2776003, -0.1381979, -0.07224751, -0.06860161, 0.07212162, 
    0.04886341, 0.05584717, 0.03996181, -0.01410723, -0.08700752, 
    -0.03988886, -0.07441044, -0.04169607, 0.1712766, 0.06304002, 
    -0.03625965, -0.08795261, -0.009339333, 0.1491408, -0.2249966, 
    -0.2931108, -0.3868942, -0.6592088, -0.6692023, -0.8078251, -1.007695, 
    -1.108932, -1.178398, -1.127242, -1.02415, -0.8737435, -0.6982226, 
    -0.5947556, -0.4056444, -0.1757622, -0.04221678, 0.003974438, 0.05854797, 
    0.08208275, 0.1886914, 0.2520375, 0.2146842, 0.1582065, -0.06086922, 
    -0.1741018, -0.2975874, -0.3884244, -0.5810184, -0.6814094, -0.7241497, 
    -0.713799, -0.578805, -0.4605432, -0.2634406, -0.007760525, 0.1083045, 
    0.5110054, 0.3697132, -0.04902059, 0.1415232, 0.05228162, -0.02735716, 
    -0.2100067, -0.280694, -0.2125945, -0.2772589, -0.2287893, -0.06197548, 
    -0.06238174, -0.07408428, -0.01622343, -0.01246309, 0.05653095, 
    0.04004335, 0.08940792, 0.07394552, 0.1829467,
  0.2935901, 0.3324573, 0.2746285, 0.00872682, -0.1237764, -0.1113093, 
    0.02171469, 0.03239202, -0.04216814, -0.1354629, -0.4139131, -0.6261044, 
    -0.7267056, -0.9104619, -0.7263799, -0.7542772, -0.5361452, -0.4092407, 
    -0.2088985, -0.0671196, 0.06245422, 0.2363634, 0.2400589, 0.3238325, 
    0.2951851, 0.2544804, 0.1319866, 0.06556416, 0.06317139, 0.1018758, 
    0.04438877, 0.2068396, 0.3790402, 0.4914584, 0.5142612, 0.2086782, 
    0.0177598, 0.2415886, -0.09833622, -0.1546831, -0.1894336, -0.4513144, 
    -0.5137491, -0.6258755, -0.9200811, -0.9304328, -0.8066697, -0.8076296, 
    -0.7117805, -0.6242476, -0.4731898, -0.2312627, 0.03939199, 0.1586461, 
    0.3266959, 0.4380407, 0.5646844, 0.579154, 0.4599481, 0.4812207, 
    0.3562536, 0.1447954, -0.1454229, -0.2557254, -0.3484993, -0.3346648, 
    -0.4822392, -0.4967251, -0.4792113, -0.433085, -0.294528, -0.116549, 
    -0.02419901, -0.05167341, 0.06782532, 0.1840198, 0.1142606, -0.2866019, 
    0.04318324, -0.004603267, 0.01629516, -0.04029667, -0.1903132, 
    -0.2169566, -0.1371226, -0.1037402, 0.03971672, 0.006351471, 0.03597403, 
    0.2072477, 0.2280154, 0.2979045, 0.3511271, 0.4065952, 0.351696, 0.4554725,
  0.3100941, 0.3600771, 0.09412718, 0.01611602, -0.02598977, -0.1993461, 
    0.1077665, 0.05364871, -0.05683279, -0.06414127, -0.2844861, -0.6135391, 
    -0.665817, -0.721839, -0.4985971, -0.5834436, -0.3303347, -0.1495895, 
    -0.03912354, 0.1013389, 0.2075076, 0.3615274, 0.3669147, 0.3783565, 
    0.3333206, 0.4076204, 0.3532104, 0.3157921, 0.2776895, 0.3602901, 
    0.2835159, 0.2575068, 0.2437372, 0.3365431, 0.3822627, 0.5109572, 
    0.3203487, 0.06484699, -0.03709054, 0.01608396, -0.04713249, -0.309453, 
    -0.4500947, -0.6104627, -0.7804494, -0.7628059, -0.5753222, -0.5623174, 
    -0.5107059, -0.2840133, -0.08274364, 0.02205753, 0.1773472, 0.3012404, 
    0.401794, 0.4272332, 0.5034218, 0.4744501, 0.3093624, 0.2575393, 
    0.02140665, -0.1051888, -0.2199016, -0.3154745, -0.3598266, -0.3142862, 
    -0.3328247, -0.2076297, -0.2231898, -0.1685514, -0.0530076, -0.1057744, 
    -0.03157282, -0.02338576, 0.2570341, 0.3086455, 0.08947241, -0.1277966, 
    0.08187133, -0.0464327, -0.05308962, -0.02908254, -0.1405083, -0.2029428, 
    -0.1318326, 0.01846027, 0.09658504, 0.3009639, 0.2676148, 0.372107, 
    0.3683147, 0.410892, 0.4186559, 0.4117222, 0.3070025, 0.4203968,
  0.3911488, 0.4843613, 0.3769885, 0.4585314, 0.2717314, -0.1476535, 
    -0.0175916, 0.03401995, -0.1896293, 0.05695295, 0.1421577, -0.3170544, 
    -0.2958958, -0.2764454, -0.3271618, -0.3469372, -0.1989388, -0.1678843, 
    -0.05707645, 0.02459669, 0.1956415, 0.3563838, 0.4270868, 0.3996129, 
    0.3509793, 0.4121447, 0.492631, 0.4570184, 0.139472, 0.3935909, 
    0.4096222, 0.2790399, 0.08332062, 0.187324, 0.4464388, 0.5560579, 
    0.3864444, 0.07838827, -0.03643918, -0.02426481, 0.0280304, -0.1279917, 
    -0.3220348, -0.5797658, -0.7706513, -1.058542, -0.9964325, -0.7781382, 
    -0.6723599, -0.5372524, -0.3546681, -0.2097788, -0.03510427, 0.1256547, 
    0.210876, 0.3011432, 0.3746295, 0.3831091, 0.3050489, 0.1773963, 
    0.03141642, -0.1050744, -0.2126918, -0.290133, -0.344902, -0.2355762, 
    -0.2648888, -0.2060995, -0.1064253, -0.094625, -0.02426386, 0.06924105, 
    0.2787466, 0.1222032, 0.5033069, 0.5937204, -0.1387341, 0.08569623, 
    0.009394109, 0.008694172, -0.03250039, -0.08526725, -0.1609998, 
    -0.002145469, -0.05299234, -0.1329241, -0.04716539, 0.2181354, 0.2074418, 
    0.2449255, 0.3145709, 0.6446815, 0.5618849, 0.4616895, 0.3283396, 
    0.3939483,
  0.4316597, 0.4245471, 0.3245959, 0.334573, 0.1482125, -0.009404689, 
    -0.04981811, -0.01399451, -0.05046916, 0.148538, 0.4832873, -0.1549451, 
    -0.1778291, 0.04743125, -0.1378227, -0.2266409, -0.05361056, -0.04000354, 
    -0.1398082, -0.0708952, 0.1559112, 0.225003, 0.2299509, 0.1134627, 
    0.02708626, 0.09329724, 0.2457548, 0.1656604, -0.05284542, 0.3240747, 
    0.1224801, 0.05700156, -0.06318074, 0.04145813, 0.3361682, 0.03084597, 
    -0.02831745, 0.06338177, 0.04441977, 0.1065784, -0.07926178, -0.1418107, 
    -0.1494439, -0.4263319, -0.4582005, -0.3860483, -0.1616669, 0.2289739, 
    0.5719271, 0.7859082, 1.034606, 1.154219, 1.057946, 0.9376993, 0.6702185, 
    0.4317093, 0.3011918, 0.1010127, -0.0800581, -0.1846809, -0.1878057, 
    -0.3384891, -0.3134732, -0.2133102, -0.1629848, -0.1169395, -0.0304327, 
    0.06813431, 0.2129748, 0.2354684, 0.2365265, 0.1528351, 0.2397652, 
    0.1276233, 0.5420274, 0.8347685, -0.04143596, -0.04817423, 0.04987264, 
    -0.05128294, -0.1085745, -0.03658557, -0.1147919, -0.1161593, -0.1380997, 
    0.01219416, 0.1024117, 0.2985382, 0.4198761, 0.3911164, 0.253535, 
    0.6415393, 0.5283396, 0.4012563, 0.3077824, 0.4598176,
  0.4876005, 0.3903674, 0.266067, 0.1056669, 0.02441686, 0.0178414, 
    -0.005970433, -0.002698958, -0.1161104, 0.1520211, 0.3754911, 0.0130237, 
    -0.1853651, -0.001706123, -0.03744841, -0.2836075, -0.1875623, 
    -0.1892712, -0.3737113, -0.2902803, -0.1070121, -0.1124483, -0.09804392, 
    0.02693972, -0.07221395, -0.00263384, 0.04344368, -0.1619437, -0.2980276, 
    0.0001493543, -0.07857776, -0.02349974, -0.02340208, -0.07620168, 
    -0.3397758, -0.5290499, -0.3701144, -0.04382825, 0.2628775, 0.2945344, 
    -0.08264697, -0.1373344, -0.1306938, -0.383721, -0.308412, -0.02568102, 
    0.1657746, 0.3250675, 0.5903349, 0.820771, 1.069827, 1.130683, 1.069893, 
    0.9635286, 0.7977409, 0.6083045, 0.4897656, 0.2532749, 0.03608751, 
    -0.2042117, -0.3575325, -0.3535118, -0.4340954, -0.53862, -0.3674936, 
    -0.2734182, -0.1444631, -0.121465, -0.03070974, 0.07859969, 0.1628121, 
    0.2284698, 0.4702503, 0.3746446, 0.1692739, 0.2473661, 0.1197131, 
    -0.04581419, 0.05514609, -0.04833698, -0.01184607, -0.003545344, 
    -0.2898084, -0.4890271, -0.3799126, -0.4040177, -0.09236366, 0.1585478, 
    0.163691, 0.2265491, 0.2218779, 0.3686064, 0.5042997, 0.596471, 
    0.3503121, 0.429023,
  0.1134306, 0.1571314, 0.04726839, -0.003903508, -0.1075819, -0.1092745, 
    0.007978201, -0.04750693, 0.03592409, 0.2496936, 0.1429391, 0.1713732, 
    -0.1369765, -0.3525352, -0.2221642, -0.4367313, -0.7180467, -0.7376277, 
    -0.6140273, -0.555873, -0.3445451, -0.111553, -0.04172802, -0.216794, 
    -0.6736784, -0.4896784, -0.1190401, -0.1592745, -0.2779919, -0.6617, 
    -0.7068655, -0.285544, -0.1602511, -0.3084607, -1.107549, -0.7584118, 
    -0.2995415, -0.1674125, 0.07519794, -0.1231906, -0.3540336, -0.6746553, 
    -0.8215466, -0.6597465, -0.4818008, -0.4526174, -0.3339813, -0.2063608, 
    -0.1954231, -0.25807, -0.216208, -0.171742, -0.1154752, -0.1298308, 
    -0.06314802, -0.1413705, -0.1871881, -0.1606576, -0.1609509, -0.2698054, 
    -0.3533338, -0.3688613, -0.5690889, -0.5684053, -0.276934, -0.09584677, 
    -0.08171915, -0.06764039, 0.1896025, 0.221943, 0.08730745, 0.04228783, 
    -0.04526067, -0.1670706, -0.1177866, 0.03747033, 0.3467968, 0.2135284, 
    6.79493e-005, -0.1604951, -0.1036105, -0.4040012, -0.4902964, -0.4379206, 
    -0.3068982, -0.4197563, -0.1230114, 0.06714141, -0.1291151, 0.08024383, 
    0.1705918, 0.1986029, 0.4421742, 0.3559434, 0.06448859, 0.05778277,
  -0.07151413, 0.07132435, 0.03901637, -0.01487303, -0.1882463, -0.1238579, 
    0.002037525, -0.06798196, 0.1805693, 0.2897327, 0.1675321, 0.1468614, 
    0.09033513, -0.1277804, -0.2231402, -0.4447241, -0.9360471, -1.119755, 
    -1.074117, -0.9303999, -0.430563, -0.153089, -0.18118, -0.6063299, 
    -0.9501266, -1.049769, -1.236081, -0.545505, -0.2852509, -0.809957, 
    -1.378854, -1.576592, -0.676104, -0.2154919, -1.068861, -0.7541638, 
    -0.4821261, -0.3684542, -0.2989554, -0.5644341, -0.5873181, -0.7664686, 
    -0.4510552, -0.16362, -0.3263972, -0.4269176, -0.162106, -0.03191423, 
    -0.1384239, -0.1257453, -0.02984667, -0.1282024, -0.1259727, -0.1818161, 
    -0.196465, -0.393373, -0.5016246, -0.5584283, -0.7604792, -0.9749646, 
    -1.29378, -1.616322, -1.792477, -1.718519, -1.669057, -1.412465, 
    -1.417836, -1.492266, -1.452764, -1.574932, -1.285951, -1.095896, 
    -1.364255, -1.019333, -0.1245739, 0.07526332, 0.0727725, 0.07431889, 
    -0.3305802, -0.4589486, -0.4072723, -0.5644822, -0.3747857, -0.2349417, 
    -0.1450653, -0.1552221, 0.1250681, 0.1159534, 0.02272415, 0.04357409, 
    -0.004457235, 0.1804228, 0.2960804, 0.1823924, 0.07329369, -0.002129555,
  0.09054649, 0.1252954, 0.135875, 0.1204619, 0.02864885, 0.1594269, 
    0.1916206, 0.0213728, 0.06837857, 0.2486842, 0.2522979, 0.2115753, 
    0.09123015, -0.2038054, -0.5222459, -0.6395311, -1.035838, -1.144432, 
    -1.163506, -0.9382124, -0.2617636, -0.1341267, -0.4154291, -1.034406, 
    -1.398027, -1.563977, -1.282548, -0.3502898, -0.4186168, -0.9302378, 
    -1.872962, -2.526934, -1.755238, -0.8967582, -1.055287, -0.741908, 
    -0.7592419, -0.7898247, -0.7045056, -0.5134249, -0.3186659, -0.2645156, 
    0.06437469, -0.2180309, -0.475338, -0.3123822, -0.1053672, -0.2588668, 
    -0.3570442, -0.2829552, -0.1940551, -0.2284465, -0.1846638, -0.1715131, 
    -0.2302365, -0.245276, -0.3116498, -0.5954881, -0.890914, -1.173483, 
    -1.527976, -1.766436, -1.999916, -2.309356, -2.612709, -2.648223, 
    -2.608607, -2.024444, -1.420652, -1.006491, -0.2556615, -0.1381159, 
    -0.7045219, -0.6492476, -0.3512487, -0.4104652, -0.3975897, -0.3382473, 
    -0.3167458, -0.2441854, -0.2417116, -0.1563926, 0.0506382, 0.04087257, 
    0.103796, 0.2069201, 0.3213735, 0.1938343, 0.31789, 0.4221383, 0.3859403, 
    0.4294627, 0.5241895, 0.3856635, -0.02835, -0.07283258,
  0.3635607, 0.3035023, 0.3865587, 0.5067737, 0.7110543, 0.9176623, 
    0.8080758, 0.4471221, 0.3145048, 0.3228707, 0.2884793, 0.4046416, 
    0.2382839, -0.2484347, -0.7452283, -0.4318485, -0.4420719, -0.715868, 
    -0.5782375, -0.3167791, 0.07420588, -0.1652956, -1.140444, -1.811341, 
    -1.767282, -1.018568, 0.01276314, 0.04214144, -0.7046518, -1.420439, 
    -1.645847, -1.441077, -1.545553, -1.517689, -1.194968, -1.196254, 
    -1.313506, -1.051576, -0.6397595, -0.225274, -0.1902637, -0.3610814, 
    -0.2594857, -0.3812141, -0.2072067, -0.1626754, -0.353138, -0.5759239, 
    -0.5712852, -0.5361447, -0.4554319, -0.350338, -0.2500448, -0.196301, 
    -0.2380652, -0.2191205, -0.329423, -0.3955851, -0.450696, -0.608037, 
    -0.7064257, -0.8199182, -1.086715, -1.270814, -1.257793, -1.119724, 
    -0.6999485, -0.1203748, -0.1304985, 0.2152698, 0.5665069, 0.03753537, 
    -0.6104949, 0.0181675, 0.1936731, 0.05997944, 0.004314423, -0.08149147, 
    -0.1093054, -0.1419883, -0.1389441, -0.06986904, 0.02505302, 0.04333019, 
    0.1827183, 0.1683307, 0.2086301, 0.279561, 0.4248891, 0.5066762, 
    0.5159696, 0.6560903, 1.060322, 0.6979356, -0.133656, -0.04127324,
  0.03200155, -0.2255667, -0.2182748, 0.04603171, 0.3484731, 0.511152, 
    0.4417021, 0.3905138, 0.5404, 0.4994983, 0.5178089, 0.4709177, 0.1451521, 
    -0.631882, -1.34876, -1.013864, -0.2595344, -0.1764297, 0.1382666, 
    0.005861282, -0.09836817, -0.4602995, -1.055287, -0.9098606, -0.3733534, 
    0.05394164, 0.1246936, 0.003795147, -0.0665499, -0.648923, -0.6715955, 
    -0.3703262, -0.8115044, -0.9252576, -0.9504206, -1.223093, -1.224705, 
    -0.8418267, -0.4171357, -0.2322073, -0.22612, -0.262773, -0.1706181, 
    -0.1960578, -0.2095342, -0.4710903, -0.7108684, -0.7574344, -0.6309366, 
    -0.4327106, -0.187089, -0.05647373, 0.06574297, 0.08737373, -0.05578995, 
    -0.07636261, -0.1808066, -0.1434855, -0.1593547, -0.1732388, -0.2378712, 
    -0.3088341, -0.250453, -0.2472138, 0.009914637, 0.4476753, 1.152786, 
    1.041605, 0.03784466, 0.115286, 0.4502795, -0.6372204, -0.470716, 
    0.4104528, 0.435811, 0.1434278, -0.05082655, -0.06295204, -0.02178955, 
    -0.1572223, -0.09438086, -0.0451622, 0.06040382, 0.121634, 0.1748252, 
    0.2055702, 0.3028193, 0.4193559, 0.4784055, 0.5828161, 0.6390657, 
    0.8173368, 0.9946155, 0.4014677, -0.1178845, -0.0009899139,
  -0.5752742, -0.7287083, -0.6309052, -0.290801, -0.08746433, 0.2017446, 
    0.4089547, 0.379495, 0.4159534, 0.2633167, 0.1864446, 0.4533396, 
    -0.1178846, -0.6522921, -0.8132133, -0.4952444, -0.3181125, -0.534307, 
    -0.2070441, -0.2275519, -0.4249806, -0.3410128, -0.2372367, 0.05047488, 
    0.3633981, 0.1945341, 0.1318064, 0.8004746, 0.5444202, -0.31961, 
    -0.2708631, -0.1016738, -0.1207654, -0.04168034, -0.3744767, -0.3317513, 
    -0.2234344, -0.1414845, 0.09437132, 0.1152868, 0.04017258, -0.03892851, 
    -0.1255984, -0.2795215, -0.3677702, -0.4443164, -0.5105429, -0.3800578, 
    -0.162138, -0.02909708, 0.05788136, 0.120398, 0.194356, 0.1141315, 
    -0.01036358, 0.04954815, 0.08372784, 0.1064005, 0.1089559, 0.2291374, 
    0.2528028, 0.3293977, 0.3241079, 0.1933942, 0.3715686, 0.6774442, 
    1.004186, 0.910908, -0.1094861, 0.08937454, 0.2146516, -0.5225873, 
    -0.09644794, 0.2465525, -0.06591463, -0.160706, -0.1074667, -0.1500292, 
    -0.2247691, -0.3534632, -0.2297816, -0.1623826, 0.02432013, 0.1480503, 
    0.163496, 0.2708206, 0.2986856, 0.2988482, 0.3745155, 0.5326695, 
    0.5341344, 0.56234, 0.4128447, -0.0727185, -0.4712049, -0.5498182,
  -0.4084611, -0.4451635, -0.2931285, 0.03322244, 0.1336288, 0.4772815, 
    0.5392932, 0.222773, 0.2498401, 0.1395695, 0.2409208, 0.2146676, 
    -0.3112602, -0.1296518, 0.4276884, 0.2667348, -0.06585002, -0.4225228, 
    -0.3369439, -0.2604301, -0.2357393, -0.0230602, 0.02518201, -0.0611949, 
    0.2355984, 0.08621705, -0.05829799, 0.6820341, 0.3573922, 0.03642863, 
    0.6499703, 0.6729846, 0.6388701, 0.9030793, 0.8893584, 0.9991243, 
    0.9105175, 0.8552277, 0.801126, 0.5066276, 0.4108429, 0.2362661, 
    0.003828049, -0.07607126, -0.1212525, -0.189775, -0.1559372, 
    0.0002479553, 0.2061234, 0.358223, 0.5012569, 0.5716338, 0.4614778, 
    0.2602577, 0.2217484, 0.2135453, 0.1836624, 0.1698112, 0.1941442, 
    0.3343787, 0.4311066, 0.5717804, 0.5284045, 0.4707222, 0.6369009, 
    0.5426469, 0.5439811, -0.005368352, -0.4358535, 0.2421093, 0.3605175, 
    0.1778359, 0.3719432, 0.3386259, 0.02259401, -0.3486299, -0.7434542, 
    -0.9447401, -1.032142, -1.048354, -0.8521454, -0.6102509, -0.306963, 
    -0.1204562, 0.02418995, 0.1408076, 0.1445837, 0.2627478, 0.3056026, 
    0.3159537, 0.3792191, 0.3473015, 0.1758652, -0.09644899, -0.3466443, 
    -0.4800916,
  0.2652535, 0.2221708, 0.2370148, 0.1734407, 0.1523793, 0.4333199, 
    0.4094104, 0.2337268, 0.2063017, 0.1555696, 0.2482617, 0.1424179, 
    0.03340149, 0.5105987, 0.3311874, -0.2615042, -0.131947, 0.02347291, 
    -0.07935911, 0.09018856, 0.1567903, 0.3205595, 0.1252797, -0.2597141, 
    -0.07512736, -0.2424939, -0.0829885, 0.5444198, 0.2158395, 0.09469694, 
    0.622122, 0.7508004, 1.046211, 1.192695, 1.58262, 1.511445, 1.185094, 
    1.073212, 0.81623, 0.4973172, 0.4710474, 0.4087918, 0.3133495, 0.268688, 
    0.1653838, 0.1631868, 0.2969756, 0.402477, 0.3799183, 0.3289254, 
    0.3032422, 0.3805046, 0.3797717, 0.3310251, 0.3004265, 0.2375193, 
    0.2233596, 0.188333, 0.2046905, 0.2673206, 0.2901561, 0.4393746, 
    0.5675322, 0.576045, 0.3946977, 0.169909, 0.1852076, -0.2766898, 
    -0.2149708, 0.4207056, 0.3409374, 0.1564483, 0.1772652, 0.04292274, 
    -0.1233207, -0.2648735, -0.4003878, -0.6154594, -0.9019828, -0.9519342, 
    -0.9333956, -0.9505017, -0.8615857, -0.7718071, -0.606019, -0.4142873, 
    -0.2873178, -0.1178679, -0.05601931, -0.00535202, 0.06945276, 0.1095901, 
    0.1401234, 0.1322293, 0.1943551, 0.2541533,
  -0.0894016, -0.1624155, -0.3320119, -0.3099582, 0.0362497, 0.4055691, 
    0.1542838, -0.05553079, -0.1236136, -0.310674, 0.1592803, 0.2349966, 
    0.1723824, 0.1145048, -0.128773, -0.3386365, -0.1406221, -0.1048312, 
    -0.005807683, 0.3104683, 0.1866238, 0.006431878, 0.04259682, 0.1067086, 
    0.198066, 0.09171849, 0.4709664, 0.7088244, -0.02664095, -0.2468071, 
    0.12012, 0.5211942, 0.7700549, 0.5366241, 1.064082, 0.7660835, 0.5198921, 
    0.1611031, 0.06582308, 0.1402209, 0.0748564, 0.1142444, 0.2230495, 
    0.2458525, 0.2552763, 0.2904651, 0.303014, 0.3986031, 0.4305529, 
    0.3175484, 0.1854684, 0.1789742, 0.1987495, 0.2275745, 0.1726426, 
    0.08154607, -0.002080917, -0.1291479, -0.1653458, -0.179473, -0.1633598, 
    0.1244495, 0.39639, 0.1636267, 0.1122262, 0.07165027, 0.09477806, 
    -0.179994, -0.2152478, -0.03303751, -0.06503621, -0.1494601, -0.2834281, 
    -0.3890921, -0.2707002, -0.08004284, 0.367923, 0.455195, 0.1774445, 
    -0.04884148, -0.3304167, -0.5702932, -0.6700978, -0.7985322, -0.832826, 
    -0.7404919, -0.5827121, -0.4453588, -0.2881484, -0.1577933, -0.2297821, 
    -0.1198866, 0.347122, 0.664635, 0.4774931, 0.2609729,
  -0.9675913, -0.750176, -0.6099255, -0.6534802, -0.210495, -0.1519501, 
    -0.4462047, -0.8671358, -0.8016736, -0.5495251, -0.4709607, -0.5403943, 
    -0.5189102, -0.4356089, -0.00455451, 0.1552273, -0.2188447, -0.507761, 
    0.07978815, 0.5734729, 0.2207711, -0.07740641, -0.02667358, 0.06653932, 
    0.002020836, -0.07988, 0.1905465, 0.245999, -0.1470837, -0.1085421, 
    0.169811, 0.1873726, 0.2588896, 0.2806507, 0.5750188, 0.6575711, 
    0.3866563, 0.07508409, -0.06493843, -0.02234459, -0.1519012, -0.2770965, 
    -0.368633, -0.3792126, -0.196465, -0.1321096, -0.135967, 0.0157094, 
    0.1240258, 0.1138859, 0.08161044, -0.02016354, -0.1804172, -0.20348, 
    -0.1752574, -0.2170054, -0.3034151, -0.4251599, -0.44238, -0.4431124, 
    -0.4147107, -0.2344699, 0.04914045, 0.3633659, 0.1220078, -0.2028453, 
    -0.2849743, -0.3578423, -0.49168, -0.1550427, 0.1140979, 0.1268584, 
    -0.1315726, -0.2862114, -0.2331679, -0.1173311, 0.07739544, 0.2048202, 
    0.3574901, 0.2410021, 0.06064749, 0.0506053, -0.06611013, -0.2955375, 
    -0.4536102, -0.6344209, -0.6084118, -0.4424615, -0.4304497, -0.4672822, 
    -0.5091118, -0.4736788, -0.1158012, 0.4140328, 0.5682642, -0.2974906,
  -1.179636, -0.7463188, -0.9547331, -0.7551568, -0.4849905, -0.454115, 
    -0.7589652, -0.8789523, -0.5664523, -0.2802706, -0.3470187, -0.632061, 
    -0.4823703, 0.07811156, 0.3357125, 0.352639, 0.02802992, 0.1692899, 
    0.7111519, 0.6744983, 0.3558785, 0.165221, 0.09923786, 0.03904903, 
    -0.05805385, 0.08649361, 0.3628771, 0.264456, -0.1492484, -0.01811242, 
    0.3433131, 0.4115263, 0.3608589, 0.1524279, -0.07935917, -0.1201957, 
    -0.08852291, -0.1344376, -0.08979213, -0.0597465, -0.1546849, -0.3716929, 
    -0.5833628, -0.5974414, -0.5489883, -0.5629854, -0.6210253, -0.6346161, 
    -0.6930306, -0.677959, -0.5243456, -0.4207001, -0.3674617, -0.370961, 
    -0.4441862, -0.41712, -0.4096162, -0.4337699, -0.4498022, -0.4591279, 
    -0.4935517, -0.4064424, -0.1665821, 0.1811714, 0.004804432, -0.3975395, 
    -0.4054985, -0.2247368, -0.2221977, -0.1848443, -0.07843131, 0.01364219, 
    0.09905885, 0.1645049, 0.118769, 0.1887889, 0.04035091, -0.08404636, 
    -0.1657522, -0.09960651, 0.0839715, 0.2595081, 0.2647657, 0.1964221, 
    0.2159052, 0.1108594, 0.004918575, -0.05525398, -0.2648082, -0.4652638, 
    -0.4459605, -0.5750628, -0.6747693, -0.4735647, -0.5800753, -1.016159,
  -1.15291, -0.7686334, -0.6939424, -0.6438936, -0.4097302, -0.4241345, 
    -0.4360814, -0.2357396, -0.01866603, -0.06656623, -0.245391, -0.252227, 
    0.03079713, 0.397122, 0.4878772, 0.4581734, 0.4506051, 0.5934762, 
    0.6163278, 0.423652, 0.3372913, 0.2846708, 0.1120308, -0.06394571, 
    -0.2112602, -0.2693006, -0.2972953, -0.4288057, -0.4581516, 0.005504131, 
    0.3028674, 0.156985, -0.0991838, -0.2803032, -0.4640921, -0.4829399, 
    -0.4197237, -0.5175265, -0.623451, -0.5254855, -0.4663547, -0.4405246, 
    -0.433428, -0.4989552, -0.7523575, -0.9495575, -1.038766, -1.123532, 
    -1.19225, -1.157468, -1.021286, -0.8331513, -0.5803032, -0.3881316, 
    -0.3252087, -0.2448535, -0.2671194, -0.3103647, -0.3158984, -0.3533497, 
    -0.3370087, -0.1836722, -0.1122692, -0.01542711, -0.1791151, -0.3211073, 
    -0.263718, -0.1355278, -0.07904987, -0.0914197, -0.1126436, 0.04101849, 
    0.2919788, 0.2019561, 0.2463732, 0.1155952, -0.06532955, -0.1437638, 
    -0.03113329, 0.1724966, 0.1819043, 0.3495636, 0.3490267, 0.3177114, 
    0.2631221, 0.1955113, 0.05182648, -0.06957674, -0.2360969, -0.4139123, 
    -0.4544077, -0.6407032, -0.999541, -1.368698, -1.651934, -1.681589,
  -0.4050264, -0.4844859, -0.5011687, -0.1896942, 0.05706668, -0.01313186, 
    -0.06685948, 0.1049342, 0.1922063, 0.05358356, -0.06850305, 0.06398404, 
    0.4006702, 0.7281767, 0.7150255, 0.5782089, 0.4784856, 0.3378446, 
    0.09557545, -0.05681705, -0.08518589, -0.1464001, -0.2389458, -0.2752739, 
    -0.3087212, -0.3488742, -0.3382783, -0.2255828, 0.007196665, 0.04437149, 
    -0.322035, -0.7590792, -0.861846, -0.7745902, -0.7874157, -0.7951956, 
    -0.6248668, -0.4746716, -0.3365531, -0.3915009, -0.5663057, -0.6723441, 
    -0.6999809, -0.7122694, -0.8244923, -0.9337536, -0.9809871, -1.060755, 
    -0.9981904, -0.8566537, -0.7528944, -0.6137342, -0.4114716, -0.2508755, 
    -0.2318816, -0.3046517, -0.4544725, -0.5467906, -0.5244107, -0.4752407, 
    -0.3247852, -0.1130178, 0.1226588, 0.01647425, -0.2157849, -0.2301241, 
    -0.244333, -0.3700494, -0.347751, -0.1589328, 0.07596314, 0.2059436, 
    0.2635121, 0.1837757, 0.03288043, -0.08040082, -0.06262779, 0.08571219, 
    0.1655464, 0.1327013, 0.07189405, 0.2614772, 0.2502794, 0.4018748, 
    0.4904165, 0.4593778, 0.2694693, 0.03611994, -0.1325812, -0.1885548, 
    -0.1450481, -0.1152148, -0.2401824, -0.5159147, -0.6857553, -0.6200814,
  0.08372664, -0.1552379, -0.1077604, 0.1075389, 0.2204621, 0.225214, 
    0.2682643, 0.4246118, 0.5485542, 0.5788437, 0.5343289, 0.4871935, 
    0.4541045, 0.4134794, 0.3435088, 0.2962104, 0.2463732, 0.1467639, 
    -0.08500683, -0.2781223, -0.3566867, -0.3717583, -0.3904594, -0.4255506, 
    -0.4895318, -0.5410616, -0.503057, -0.332387, -0.1421196, -0.2353814, 
    -0.561016, -0.7900851, -0.7383598, -0.6953422, -0.7734346, -0.7184379, 
    -0.4285941, -0.1994601, -0.07512724, -0.234307, -0.356768, -0.3394991, 
    -0.467559, -0.2788545, -0.1884249, -0.1682588, -0.2667452, -0.3248345, 
    -0.2683893, -0.2037082, -0.1188445, -0.1165659, -0.1278942, -0.1923311, 
    -0.3780406, -0.5389454, -0.5785451, -0.5161266, -0.4394338, -0.3247693, 
    -0.1912735, 0.06828082, 0.01476526, -0.04361725, -0.05855823, 0.05823803, 
    0.132278, 0.1668156, 0.2545927, 0.3432971, 0.3900908, 0.3970406, 
    0.3767769, 0.3079131, 0.2870471, 0.3989611, 0.4811223, 0.5016139, 
    0.3660508, 0.2612659, 0.3420601, 0.3143749, 0.4596545, 0.5870306, 
    0.6565781, 0.5731797, 0.3664093, 0.223326, 0.2351594, 0.2838736, 
    0.3200226, 0.3399935, 0.3400745, 0.2177927, 0.2230825, 0.2179394,
  0.1898137, 0.1638372, 0.1716335, 0.466995, 0.6412135, 0.7570176, 0.7109565, 
    0.8129421, 0.6941761, 0.6480822, 0.6098011, 0.5275419, 0.4524444, 
    0.5197295, 0.5891141, 0.6379424, 0.6023303, 0.4291532, 0.1620145, 
    -0.09801149, -0.2391086, -0.326576, -0.436309, -0.5950491, -0.6855441, 
    -0.6668428, -0.4575818, -0.2138318, -0.1540499, -0.3695934, -0.788783, 
    -1.010967, -0.9161756, -0.6125947, -0.3879691, -0.2663057, -0.2095025, 
    -0.1849744, -0.07459021, -0.09462631, -0.07476926, -0.08396518, 
    -0.0423474, 0.07467735, 0.3374866, 0.4705757, 0.4874541, 0.4507352, 
    0.3949248, 0.3347848, 0.2751656, 0.197773, 0.1857288, 0.1805042, 
    0.0638212, -0.07019579, -0.166436, -0.188197, -0.1032361, -0.0100069, 
    0.09785438, 0.09428966, 0.1949248, 0.175231, 0.1830105, 0.1736356, 
    0.2377795, 0.3749378, 0.5095243, 0.5204781, 0.482734, 0.5495797, 
    0.4680693, 0.6521189, 0.8426787, 1.01636, 1.048733, 0.9649277, 0.7536322, 
    0.7747099, 0.6554552, 0.7682972, 0.6921253, 0.6267608, 0.6824573, 
    0.6561878, 0.4606636, 0.3399277, 0.3972518, 0.5285351, 0.5957875, 
    0.6262238, 0.6480663, 0.5943389, 0.4646997, 0.4536159,
  0.5188667, 0.3342476, 0.3785021, 0.4951851, 0.6105824, 0.5739612, 
    0.7339221, 0.7388537, 0.7488148, 0.7949411, 0.7920765, 0.6896514, 
    0.5618356, 0.4742542, 0.433499, 0.4095569, 0.2667349, 0.0661, -0.1894503, 
    -0.4184216, -0.6137668, -0.7590466, -0.806296, -0.7857067, -0.6867159, 
    -0.5486462, -0.4742973, -0.4413708, -0.5684542, -0.7715954, -0.9576144, 
    -0.9190401, -0.6146456, -0.2952934, -0.1664358, -0.1719372, -0.1704561, 
    -0.1502088, -0.1302379, -0.1027965, -0.09848344, -0.04713255, 0.06691368, 
    0.2197782, 0.3437693, 0.3623728, 0.3375356, 0.3044789, 0.4272165, 
    0.5889027, 0.6437528, 0.6081897, 0.7271677, 0.6425322, 0.5362823, 
    0.3543648, 0.2520211, 0.2920113, 0.2999378, 0.2597196, 0.2677435, 
    0.2717799, 0.2370956, 0.227493, 0.2064807, 0.1938342, 0.2388212, 
    0.3778023, 0.5662789, 0.6452177, 0.6420927, 0.3876819, 0.5957385, 
    0.7325062, 0.7253771, 0.6167347, 0.9238635, 0.9884144, 0.6295114, 
    0.7157907, 0.9462756, 0.8490751, 0.6936393, 0.597594, 0.5494655, 
    0.8443062, 0.8717802, 0.8792672, 0.9244332, 1.017923, 1.066149, 1.061331, 
    1.056855, 1.110029, 1.037714, 0.7659208,
  0.8552926, 0.8641304, 0.8138537, 1.016344, 1.069127, 1.090693, 0.8225615, 
    0.9372262, 0.8796741, 0.8395536, 0.7560738, 0.6661161, 0.5518746, 
    0.4642769, 0.3529, 0.2538115, 0.09723598, -0.09750676, -0.3711885, 
    -0.628594, -0.8221163, -0.8295545, -0.7124809, -0.5481743, -0.4475883, 
    -0.3918916, -0.4434053, -0.4940075, -0.5146944, -0.5447237, -0.467738, 
    -0.3381482, -0.209893, -0.1512667, -0.139255, -0.1877576, -0.1324027, 
    -0.07009806, -0.04335651, -0.09106159, -0.1587862, -0.1281547, 
    -0.0479138, 0.04676394, 0.08546835, 0.08677042, 0.1318877, 0.3199899, 
    0.5099313, 0.6938667, 0.7556019, 0.4218617, 0.6282417, 0.4868355, 
    0.3767118, 0.2945667, 0.2306995, 0.1820666, 0.1699248, 0.1464221, 
    0.07527956, 0.09098593, 0.1862333, 0.313219, 0.4362659, 0.5183948, 
    0.597301, 0.6685413, 0.6538277, 0.5997099, 0.5650745, 0.6234241, 
    0.6970569, 0.6868681, 0.3558785, 0.1962268, 0.2087105, 0.4985055, 
    0.4336455, 0.3223174, 0.03880507, 0.03764927, 0.09329677, 0.1665227, 
    0.292923, 0.3550153, 0.5683132, 0.8349636, 0.9086615, 0.9074736, 
    0.8482289, 0.9633005, 0.7740426, 0.7971058, 0.8377144, 0.861917,
  0.7224801, 0.8341174, 0.9205595, 0.9570992, 0.9294626, 1.22847, 1.229251, 
    1.078942, 0.8995471, 0.7266955, 0.5995796, 0.5571317, 0.5215198, 
    0.4410673, 0.1784371, -0.02074909, -0.2267549, -0.4057751, -0.5235811, 
    -0.5993136, -0.581768, -0.4709119, -0.3265759, -0.191973, -0.1154758, 
    -0.07094443, -0.04884154, -0.01866573, -0.0001760721, -0.001917541, 
    -0.01895863, -0.0415172, -0.04275441, -0.002145648, 0.05298138, 
    -0.01947963, -0.1297334, -0.1436821, -0.177699, -0.1647758, -0.1079885, 
    0.007554948, 0.1451038, 0.2993681, 0.4394885, 0.65679, 0.8775094, 
    0.9631051, 0.9539416, 0.5659859, 0.3726265, 0.2864286, 0.2766632, 
    0.523717, 0.4981636, 0.4214711, 0.3854846, 0.3181669, 0.312454, 
    0.4940621, 0.6484892, 0.8164904, 0.9798043, 1.121145, 1.16081, 1.083597, 
    0.9265165, 0.7484566, 0.5840035, 0.3104195, 0.4155465, 0.4101754, 
    0.3791533, 0.1605497, 0.06149375, -0.06785196, -0.0943656, -0.07579473, 
    -0.07647827, -0.06269243, -0.1071911, -0.08959663, 0.001598001, 
    0.03258753, 0.07610971, 0.08522421, 0.07526326, 0.07552367, 0.1563993, 
    0.2019722, 0.1584013, 0.191344, 0.2414091, 0.2782906, 0.4039254, 0.5683297,
  0.1863474, 0.3645863, 0.5384631, 0.6818388, 0.7893258, 0.772415, 0.6150256, 
    0.3967803, 0.1976428, 0.0537138, -0.05240601, -0.1273572, -0.2073865, 
    -0.2885225, -0.3896618, -0.7762341, -0.5002738, -0.489141, -0.4440727, 
    -0.665199, -0.5297823, -0.3677707, -0.2523734, -0.1851373, -0.1465955, 
    -0.1405083, -0.1199679, -0.1078422, -0.1125785, -0.08285856, -0.06648481, 
    0.01564407, 0.1337428, 0.266865, 0.3631866, 0.1971056, 0.2474475, 
    0.2984403, 0.7059927, 0.9318063, 0.7175971, 0.8698107, 0.9336127, 
    0.969355, 0.9946479, 1.024596, 1.024368, 0.9506213, 0.8278512, 0.711331, 
    0.6020861, 0.521536, 0.5103543, 0.5660347, 0.6227241, 0.6889351, 
    0.7615914, 0.8000354, 0.8145862, 0.8307158, 0.8394886, 0.8397652, 
    0.7782906, 1.039293, 0.8428739, 0.5955921, 0.3816109, 0.2104196, 
    0.08992797, 0.004820555, 0.08581012, 0.1493193, 0.08200155, 0.1893421, 
    0.1659859, 0.1872262, 0.1797392, 0.1969755, 0.1996285, 0.07806265, 
    0.015172, 0.07550728, -0.02021199, -0.01710325, -0.02362996, -0.03803426, 
    -0.07192093, -0.08282596, -0.0281547, 0.03551716, -0.04713255, 
    -0.007549223, -0.06230181, -0.04929727, -0.0301241, 0.04240194,
  -0.353171, -0.3871716, -0.4064425, -0.3851535, -0.3582816, -0.3476695, 
    -0.4312309, -0.4963838, -0.5454561, -0.5712537, -0.5969861, -0.6284477, 
    -0.6260876, -0.6035942, -0.5621554, -0.5172498, -0.4906384, -0.4193819, 
    -0.3530896, -0.2844535, -0.2373017, -0.2254202, -0.1949842, -0.1559868, 
    -0.1314914, -0.1157854, -0.07125401, -0.001120329, 0.05164647, 0.1112819, 
    0.178714, 0.2892443, 0.3037137, 0.374498, 0.4245957, 0.60373, 0.7738795, 
    0.8892115, 0.9869658, 1.055732, 1.138056, 1.174042, 1.154316, 1.078665, 
    0.9643258, 0.8271188, 0.6911488, 0.5704292, 0.4912951, 0.4564155, 
    0.4535673, 0.4715034, 0.5211455, 0.5720731, 0.608027, 0.6218291, 
    0.6028512, 0.5653837, 0.5232126, 0.4505889, 0.3434274, 0.2137073, 
    0.08955365, 0.07544231, 0.05641568, 0.2378283, 0.2066434, 0.2144884, 
    0.2338408, 0.2941272, 0.3804716, 0.4812854, 0.5481638, 0.5422717, 
    0.5718127, 0.3455269, 0.4128609, 0.2857774, 0.1409208, 0.02908814, 
    -0.04029667, -0.06733114, -0.04672566, -0.02743854, -0.003366292, 
    0.005373955, -0.004114985, -0.000762105, -0.01104859, -0.01565468, 
    -0.04187539, -0.1990369, -0.1366182, -0.1711072, -0.2800753, -0.3298799,
  -0.3836885, -0.4146781, -0.4513806, -0.4156547, -0.412432, -0.3747693, 
    -0.383005, -0.3613253, -0.3681937, -0.338197, -0.3111788, -0.2926241, 
    -0.2733696, -0.2513806, -0.2306612, -0.2144503, -0.1859021, -0.1559704, 
    -0.1269991, -0.1004853, -0.07190454, -0.08679724, -0.1127414, 
    -0.07590866, 0.0283556, 0.2082548, 0.2742703, 0.3609565, 0.4784045, 
    0.5625353, 0.6071154, 0.6499702, 0.7029487, 0.7627958, 0.8241403, 
    0.8630074, 0.8677275, 0.8398141, 0.7906604, 0.7257841, 0.6528186, 
    0.5747424, 0.4928902, 0.4293161, 0.3699086, 0.3341338, 0.3190296, 
    0.3191598, 0.334801, 0.3551787, 0.3741565, 0.3862496, 0.3924019, 
    0.3773141, 0.3443876, 0.2961943, 0.2626168, 0.2241077, 0.2047229, 
    0.1916045, 0.1911975, 0.2112171, 0.2282255, 0.2548043, 0.286445, 
    0.3185901, 0.3469267, 0.3469104, 0.3398954, 0.3344918, 0.3279488, 
    0.5948107, 0.4767118, 0.3067575, 0.2767606, 0.2212756, 0.1565295, 
    0.09313437, 0.02876261, -0.02833372, -0.0735974, -0.112432, -0.1314913, 
    -0.1452771, -0.1708956, -0.1919405, -0.2382296, -0.2720512, -0.2883109, 
    -0.2918429, -0.2766899, -0.274932, -0.2655896, -0.2843722, -0.3112764, 
    -0.3391899,
  -0.3257133, -0.3006807, -0.2908826, -0.2717908, -0.235251, -0.1961398, 
    -0.1659965, -0.1423637, -0.127227, -0.1128715, -0.104766, -0.1004529, 
    -0.1001274, -0.09905313, -0.1039197, -0.1033012, -0.09882526, 
    -0.07618529, -0.03860392, 0.01139608, 0.07098269, 0.1303739, 0.1924508, 
    0.2518259, 0.3170602, 0.3959501, 0.463219, 0.5055529, 0.5584338, 
    0.6257353, 0.6795764, 0.7351917, 0.7861519, 0.8223987, 0.8466825, 
    0.8610542, 0.8675483, 0.8465362, 0.8074248, 0.7589059, 0.706139, 
    0.6518584, 0.5974801, 0.5421416, 0.4898954, 0.4453642, 0.3998238, 
    0.353193, 0.3111194, 0.2728056, 0.2359892, 0.1930693, 0.1615751, 
    0.1221708, 0.07711875, 0.04192993, 0.009768486, -0.01155311, -0.02808958, 
    -0.02545288, -0.009827852, 0.008498967, 0.02702111, 0.04228802, 
    0.04858685, 0.06107056, 0.07910442, 0.09808229, 0.1099638, 0.121829, 
    0.1270048, 0.1217639, 0.1129586, 0.09054643, 0.08498001, 0.04769167, 
    -0.001185298, -0.0671358, -0.1157361, -0.1766573, -0.2355603, -0.2850883, 
    -0.2913546, -0.3172822, -0.3103486, -0.3586071, -0.3941378, -0.4157036, 
    -0.4305473, -0.4423148, -0.442982, -0.4160453, -0.3967094, -0.3807589, 
    -0.3550915, -0.341029,
  -0.2868786, -0.2511202, -0.2106742, -0.1735649, -0.1320772, -0.09447956, 
    -0.0577608, -0.03035196, -0.01051146, 0.01395143, 0.0400582, 0.06533489, 
    0.08841433, 0.1111357, 0.1279325, 0.149775, 0.1729521, 0.1937854, 
    0.2153349, 0.2414579, 0.2726917, 0.2931344, 0.3182158, 0.3509631, 
    0.3734729, 0.4019885, 0.4263212, 0.4463407, 0.4729358, 0.4958199, 
    0.5161812, 0.5357125, 0.5509468, 0.5599638, 0.5626168, 0.5558297, 
    0.5446969, 0.5339872, 0.5141793, 0.4934762, 0.4588896, 0.4246448, 
    0.3899931, 0.3587594, 0.3220081, 0.2845732, 0.2489937, 0.2143095, 
    0.1812203, 0.1532581, 0.1179228, 0.08458945, 0.06268188, 0.03637981, 
    0.00916627, -0.01853555, -0.04150106, -0.06521523, -0.08334675, 
    -0.100225, -0.1163708, -0.1281547, -0.1469047, -0.1609184, -0.1811983, 
    -0.1972302, -0.2155408, -0.2367973, -0.2527315, -0.2714815, -0.2937797, 
    -0.3157849, -0.3448865, -0.3762015, -0.4010713, -0.4311494, -0.4550427, 
    -0.4841769, -0.5055147, -0.5254203, -0.5441215, -0.5555473, -0.5612439, 
    -0.5652966, -0.5643852, -0.5562797, -0.5445935, -0.531003, -0.5089327, 
    -0.4862602, -0.4606905, -0.435544, -0.4032524, -0.3818005, -0.3534314, 
    -0.3228976,
  -0.4758687, -0.4520569, -0.4270732, -0.4021548, -0.3787662, -0.357705, 
    -0.3398012, -0.3253807, -0.3144756, -0.3074933, -0.3040918, -0.303473, 
    -0.3053613, -0.309788, -0.3154683, -0.3217835, -0.3286028, -0.3349671, 
    -0.3399639, -0.3442612, -0.3474507, -0.3490944, -0.348834, -0.3462138, 
    -0.3406634, -0.3313375, -0.318284, -0.3008847, -0.2786031, -0.2514057, 
    -0.2195535, -0.183063, -0.1434469, -0.1019111, -0.05700469, -0.01255488, 
    0.03207397, 0.07611632, 0.1181089, 0.1574968, 0.1941019, 0.2275978, 
    0.2575295, 0.284043, 0.3070085, 0.3262959, 0.3333108, 0.3420348, 
    0.3490663, 0.3254011, 0.3303652, 0.2929463, 0.2701759, 0.3465919, 
    0.3272562, 0.339447, 0.3406677, 0.3303161, 0.296999, 0.2505474, 
    0.2535748, 0.257318, 0.23419, 0.2041116, 0.1765404, 0.1485782, 0.1197853, 
    0.08371782, 0.05118179, 0.03181362, 0.006650925, -0.02404594, 
    -0.05882788, -0.183063, -0.07090425, -0.106679, -0.08439732, -0.2982159, 
    -0.2184467, -0.2425356, -0.2754788, -0.3120832, -0.3483138, -0.3856673, 
    -0.4190817, -0.4517641, -0.4808006, -0.5052638, -0.5246487, -0.5385804, 
    -0.5461812, -0.5488505, -0.5449605, -0.5337629, -0.5177803, -0.4978738,
  -0.05088544, -0.03561825, -0.02468085, -0.02127915, -0.02433904, 
    -0.0323143, -0.0438703, -0.05588201, -0.06717747, -0.07756156, 
    -0.08898729, -0.1008525, -0.1123435, -0.1250879, -0.1389877, -0.1542546, 
    -0.1707585, -0.1896875, -0.2117739, -0.2404199, -0.2742736, -0.3159242, 
    -0.3643289, -0.4159894, -0.4610415, -0.4970279, -0.5221901, -0.5382876, 
    -0.5492086, -0.5545144, -0.5523014, -0.5431218, -0.5265856, -0.5008693, 
    -0.4636135, -0.4150457, -0.3564358, -0.2907939, -0.222939, -0.1570697, 
    -0.104531, -0.06318998, -0.03312808, 0.01156598, 0.0274837, 0.006552696, 
    0.06161499, 0.07295942, 0.08199263, 0.06091499, 0.09781289, 0.1459899, 
    0.09325552, 0.1740823, 0.04449272, 0.2959414, 0.3241153, 0.3283954, 
    0.3736758, 0.3764749, 0.3756933, 0.3659444, 0.3191018, 0.2473574, 
    0.1722269, 0.1163352, 0.04968441, -0.0232811, -0.0375551, -0.03887355, 
    -0.02243477, -0.017389, -0.01590788, -0.02497363, -0.05243134, 
    -0.0759341, -0.09860641, -0.1504948, -0.1651433, -0.2072978, -0.2529359, 
    -0.2524965, -0.2943907, -0.3061261, -0.3569565, -0.349534, -0.3136454, 
    -0.2976131, -0.2788472, -0.2574606, -0.2297754, -0.1980534, -0.1597717, 
    -0.1275616, -0.09735322, -0.0715723,
  0.1551042, 0.1261169, 0.09528986, 0.08467789, 0.08799821, 0.09719416, 
    0.1087176, 0.1192319, 0.1250588, 0.1263283, 0.1189064, 0.1067808, 
    0.09309256, 0.07321954, 0.04179072, -0.004693508, -0.06691742, 
    -0.1496482, -0.2497129, -0.3493061, -0.4301009, -0.4620831, -0.4089258, 
    -0.2862529, -0.1935285, -0.1681377, -0.2121648, -0.2809309, -0.3542218, 
    -0.4339256, -0.5227437, -0.6280172, -0.744277, -0.835, -0.8897691, 
    -0.9029198, -0.8753643, -0.8092995, -0.7142477, -0.6011944, -0.4870501, 
    -0.3627996, -0.2100973, -0.1207581, -0.04997396, -0.04553044, 
    -0.05197579, -0.06214827, -0.06921208, -0.08286768, -0.09688136, 
    -0.1049055, -0.1050356, -0.09408188, -0.06940737, -0.03259075, 
    -0.0150128, 0.004127622, 0.01846683, 0.04177415, 0.05372071, 0.04885423, 
    0.02844405, -0.01016259, -0.06768209, -0.1433006, -0.2283267, -0.297858, 
    -0.3393779, -0.3451884, -0.3277897, -0.2915103, -0.2413801, -0.2049218, 
    -0.2013897, -0.1928448, -0.2149315, -0.2998436, -0.2926494, -0.3155338, 
    -0.3492249, -0.3915589, -0.3959858, -0.4132059, -0.4007711, -0.4337952, 
    -0.3988831, -0.291038, -0.2032614, -0.08552074, 0.03580141, 0.1110778, 
    0.1999612, 0.2470641, 0.2424092, 0.2123961,
  0.2513609, 0.2026949, 0.1947689, 0.1732197, 0.1558208, 0.1455178, 
    0.1376405, 0.1367774, 0.1585872, 0.1914649, 0.2109147, 0.2089618, 
    0.2000588, 0.2016375, 0.2005145, 0.1716733, 0.1161721, 0.03570342, 
    -0.03677368, -0.0656147, -0.1198635, -0.2007713, -0.249681, -0.2646222, 
    -0.2532129, -0.2305402, -0.220986, -0.204401, -0.1977441, -0.2197328, 
    -0.2809146, -0.3748925, -0.5021546, -0.6534733, -0.7987694, -0.936269, 
    -1.069521, -1.1753, -1.240062, -1.266755, -1.224094, -1.07958, 
    -0.8306704, -0.4964252, -0.2563701, -0.1419983, -0.3256409, -0.2480208, 
    -0.2610415, -0.3322492, -0.4005922, -0.4260969, -0.4178447, -0.3941633, 
    -0.348216, -0.3191307, -0.3147036, -0.1660547, -0.1349183, -0.08029604, 
    -0.01392221, 0.1046977, 0.2191508, 0.3580182, 0.4309671, 0.4537375, 
    0.3969662, 0.2614522, 0.1460876, 0.06080151, -0.009641647, -0.05007124, 
    -0.08234668, -0.1165915, -0.08807564, -0.170742, -0.1985251, -0.1673079, 
    -0.1225649, -0.224404, -0.1023826, -0.07051396, -0.05065751, -0.04889965, 
    -0.08753908, -0.1540103, -0.2450256, -0.3040099, -0.2982483, -0.2412658, 
    -0.09247065, 0.03441763, 0.2184505, 0.3119397, 0.3245053, 0.2822366,
  0.07430983, 0.00276041, -0.04413128, -0.06748676, -0.04087591, -0.05557251, 
    -0.01530552, 0.04509497, 0.1018982, 0.1651626, 0.2825127, 0.3947859, 
    0.4833431, 0.4933858, 0.433701, 0.5044534, 0.5448344, 0.4180439, 
    0.2802508, 0.1606219, 0.2735939, 0.280673, 0.2134218, 0.1459255, 
    0.05274439, -0.04035473, -0.08353472, -0.1309314, -0.1772685, -0.2173724, 
    -0.2564678, -0.2825258, -0.3112528, -0.383193, -0.5169985, -0.6776267, 
    -0.8346748, -0.9403384, -0.98124, -0.9853906, -0.947093, -0.8490624, 
    -0.680491, -0.4448469, -0.2136617, -0.08353508, -0.1796615, -0.1663638, 
    -0.2424543, -0.2946842, -0.3319563, -0.3505598, -0.3421614, -0.3296126, 
    -0.3108789, -0.291608, -0.3085351, -0.291429, -0.2268294, -0.1497946, 
    -0.04416326, 0.05324885, 0.1245867, 0.1942645, 0.2403909, 0.2754005, 
    0.2949969, 0.2977474, 0.3121029, 0.3133398, 0.2644957, 0.1801692, 
    0.1433692, 0.1102962, 0.08822596, -0.02178383, -0.1097883, -0.1916893, 
    -0.2054914, -0.2672426, -0.08835259, 0.03903987, 0.1842872, 0.2986428, 
    0.3613705, 0.3737565, 0.3386328, 0.2930274, 0.2569435, 0.2508075, 
    0.3513608, 0.2280531, 0.3428812, 0.3353133, 0.2158303, 0.1978774,
  0.1012633, 0.05461597, -0.205605, -0.2374897, -0.2198958, -0.1657777, 
    -0.1709208, -0.04616499, -0.1199441, -0.2107158, -0.2409892, -0.2213926, 
    -0.170351, -0.02930307, 0.06897163, 0.1979592, 0.3685156, 0.374424, 
    0.2795023, 0.175791, 0.07973027, 0.1231217, 0.2881279, 0.3749619, 
    0.4547462, 0.516921, 0.5332937, 0.4978781, 0.3902931, 0.2498951, 
    0.1096125, -0.03273773, -0.1079655, -0.1924381, -0.2620015, -0.335309, 
    -0.3741107, -0.4071679, -0.4147849, -0.3621807, -0.3292542, -0.2930725, 
    -0.3028545, -0.2639713, -0.215843, -0.1711164, -0.07736639, 0.03679389, 
    0.1809344, 0.2722266, 0.2806088, 0.2872006, 0.3085386, 0.3559668, 
    0.3800552, 0.3690858, 0.2823832, 0.1545024, 0.01493549, -0.07360649, 
    -0.08775043, -0.0423727, -0.01732373, -0.05692339, -0.1130757, 
    -0.1451559, -0.1593812, -0.1516666, -0.1418521, -0.1166241, -0.1473372, 
    -0.1244043, -0.05399418, 0.06382811, 0.172585, 0.2055275, 0.1790138, 
    0.1455177, -0.0100975, -0.06478494, -0.04041982, 0.02128255, 0.117816, 
    0.2171325, 0.3312599, 0.419232, 0.5029885, 0.6004819, 0.6876564, 
    0.7541115, 0.8122982, 0.8312111, 0.8476663, 0.7924089, 0.6199646, 
    0.3852642,
  0.6851336, 0.4701108, 0.2582131, 0.1331642, 0.05497396, 0.02128255, 
    0.02471685, 0.05066085, 0.04924506, 0.04070002, 0.02069677, -0.0415591, 
    -0.1106185, -0.2171286, -0.3318913, -0.3827699, -0.3862855, -0.3564841, 
    -0.2786685, -0.2114159, -0.1272525, -0.01638001, 0.1079202, 0.2609963, 
    0.388731, 0.4893653, 0.5637466, 0.6672136, 0.7409439, 0.7689065, 
    0.7446389, 0.6892357, 0.7057233, 0.5769792, 0.5463157, 0.3948998, 
    0.2825134, 0.2030699, 0.1120381, 0.0357523, 0.02387071, 0.08558941, 
    0.197129, 0.2824317, 0.3346779, 0.376605, 0.3990009, 0.4776303, 
    0.6182715, 0.8066828, 0.9032981, 1.013715, 1.025596, 1.105837, 1.15115, 
    1.215668, 1.134141, 1.017393, 0.8820412, 0.7455015, 0.6651304, 0.6947856, 
    0.7553487, 0.7697692, 0.7587996, 0.7963805, 0.8481221, 0.9752216, 
    1.073903, 1.026736, 0.9374776, 0.7049906, 0.6281514, 0.5513284, 0.431488, 
    0.3903906, 0.430397, 0.4765885, 0.4690202, 0.4676204, 0.4890399, 
    0.4514425, 0.4157655, 0.373626, 0.3486915, 0.3776791, 0.4425063, 
    0.4974707, 0.5510352, 0.5417579, 0.5672135, 0.6738052, 0.8045998, 
    0.8721454, 0.9031512, 0.8349221,
  0.9392025, 0.807904, 0.6408303, 0.4555275, 0.3022401, 0.1812277, 0.1078553, 
    0.06044316, 0.06023097, 0.1126723, 0.2227473, 0.3429782, 0.3907814, 
    0.3223732, 0.1969336, 0.08664703, -0.002805948, -0.02116537, 0.01018214, 
    0.06700182, 0.1469173, 0.222259, 0.35167, 0.468776, 0.5316014, 0.4949479, 
    0.4358008, 0.4407487, 0.5637141, 0.7461686, 0.9030048, 1.053493, 
    1.068255, 1.247748, 1.497568, 1.538926, 1.274684, 1.379209, 1.347959, 
    1.427337, 1.512233, 1.767019, 1.915635, 2.166953, 2.498415, 2.492718, 
    2.286322, 2.054209, 1.731813, 1.683148, 1.78432, 1.733881, 1.65486, 
    1.570665, 1.38004, 1.298171, 1.402126, 1.498057, 1.717963, 1.886827, 
    2.06666, 2.165456, 2.277435, 2.288747, 2.245486, 2.186078, 2.076638, 
    2.039236, 2.146055, 2.200466, 2.108018, 2.035004, 2.038845, 2.002744, 
    1.882953, 1.851427, 1.869427, 1.948513, 2.035606, 2.004535, 1.765391, 
    1.404486, 1.172683, 1.041384, 0.942621, 0.8596454, 0.8023703, 0.7508075, 
    0.684597, 0.6240337, 0.5888286, 0.6206808, 0.6848409, 0.7838807, 
    0.9161398, 0.9668233,
  1.161469, 1.142588, 1.210378, 1.24057, 1.147292, 1.144362, 1.104259, 
    1.143598, 1.17374, 1.176036, 1.106049, 1.077842, 1.358246, 1.629079, 
    1.978656, 2.256407, 2.295111, 2.394965, 2.407383, 1.829047, 0.9101501, 
    0.5375099, 0.4731226, 0.6180768, 0.9422464, 1.307237, 1.509727, 1.709109, 
    1.913096, 2.003412, 1.843076, 1.693777, 1.57571, 1.606341, 1.721251, 
    1.853102, 1.918532, 1.871088, 1.832237, 1.929698, 2.099961, 2.176931, 
    2.129128, 1.958441, 1.860166, 1.88253, 1.868174, 1.705593, 1.592654, 
    1.660882, 1.808995, 1.885101, 1.908913, 1.950987, 1.946706, 1.826622, 
    1.707807, 1.709987, 1.769655, 1.840504, 1.956244, 2.093011, 2.171657, 
    2.165977, 2.165423, 2.232383, 2.278217, 2.287445, 2.242735, 2.183197, 
    2.143907, 2.088486, 1.966726, 1.813991, 1.774668, 1.87055, 1.875987, 
    1.723805, 1.590179, 1.635654, 1.755365, 1.786077, 1.80154, 1.908539, 
    1.784369, 1.662087, 1.603737, 1.491693, 1.180544, 1.002826, 0.9831648, 
    1.06601, 1.145844, 1.083555, 0.9684672, 1.07737,
  1.54612, 1.386468, 1.157855, 1.014773, 0.9788189, 0.9341903, 0.8759212, 
    0.8077569, 0.6426854, 0.5940857, 0.5696392, 0.5602961, 0.6181898, 
    0.7431412, 0.8730412, 1.007854, 1.128803, 1.243305, 1.447423, 1.687169, 
    1.883865, 1.752289, 1.383036, 1.335589, 1.422488, 1.594803, 1.756423, 
    1.861665, 1.964269, 2.07195, 2.157562, 2.136778, 2.026946, 1.876197, 
    1.772341, 1.765863, 1.762624, 1.690473, 1.585199, 1.575336, 1.685606, 
    1.728916, 1.591091, 1.375401, 1.302354, 1.362721, 1.383832, 1.233132, 
    1.058197, 1.139642, 1.3685, 1.540603, 1.636566, 1.743142, 1.828005, 
    1.825596, 1.755902, 1.713112, 1.613535, 1.541221, 1.665782, 1.92055, 
    2.053852, 2.008473, 1.991319, 2.055219, 2.100238, 2.093467, 2.047113, 
    1.962641, 1.928753, 1.914838, 1.80014, 1.631455, 1.603314, 1.597617, 
    1.308652, 0.8864198, 0.6553326, 0.7027926, 0.89013, 1.004859, 1.060687, 
    0.9821386, 1.001295, 1.085248, 1.195404, 1.478135, 1.648366, 1.675319, 
    1.636501, 1.555609, 1.620502, 1.538177, 1.482677, 1.521804,
  1.124978, 1.083539, 0.9812756, 0.8540626, 0.7618423, 0.7420831, 0.7480888, 
    0.7437921, 0.7125425, 0.700839, 0.7204361, 0.7343683, 0.6802015, 
    0.6005478, 0.5656033, 0.5996695, 0.7087517, 0.859745, 0.9650993, 
    0.9845638, 0.9925566, 1.064009, 1.185768, 1.297601, 1.342996, 1.375596, 
    1.42991, 1.466644, 1.512282, 1.621429, 1.718989, 1.774864, 1.811159, 
    1.762136, 1.617475, 1.497261, 1.430609, 1.346738, 1.263584, 1.267816, 
    1.365652, 1.380349, 1.199538, 1.0289, 0.9876566, 0.9958439, 0.9539003, 
    0.8610125, 0.6828713, 0.5492454, 0.6006937, 0.8138287, 1.040179, 
    1.307334, 1.552582, 1.665798, 1.639284, 1.489545, 1.23948, 1.039756, 
    1.033002, 1.274213, 1.54433, 1.681862, 1.71946, 1.709955, 1.683978, 
    1.626068, 1.571788, 1.512136, 1.505641, 1.586387, 1.626524, 1.631146, 
    1.619704, 1.347552, 0.7477479, 0.6509542, 0.880332, 0.9209738, 0.6809673, 
    0.5978451, 0.6302996, 0.4845467, 0.3747816, 0.4441338, 0.6103621, 
    0.774766, 0.8878508, 1.003525, 1.149668, 1.243694, 1.247845, 1.220289, 
    1.191676, 1.159792,
  1.141156, 1.087005, 1.111549, 1.110475, 1.041221, 0.9571223, 0.934238, 
    0.9478617, 0.9334898, 0.9047298, 0.8745542, 0.8047628, 0.6687593, 
    0.5378838, 0.4992776, 0.5126228, 0.5609646, 0.6391211, 0.6654081, 
    0.7062607, 0.7889261, 0.7511501, 0.6206484, 0.6172304, 0.7705994, 
    0.9834738, 1.204762, 1.310069, 1.309793, 1.311453, 1.283164, 1.220615, 
    1.233881, 1.237624, 1.17314, 1.111779, 1.008849, 0.8603621, 0.708457, 
    0.6162205, 0.7140718, 0.7352152, 0.4164653, 0.1478128, 0.181016, 
    0.1652446, -0.001633644, -0.1157777, -0.2011781, -0.2454653, -0.2201073, 
    -0.07982397, 0.1083108, 0.3458596, 0.6471617, 0.9470966, 1.104698, 
    1.078884, 0.8812276, 0.6334572, 0.4890401, 0.4405537, 0.5135679, 
    0.7024026, 0.8896911, 1.131439, 1.302533, 1.28917, 1.199018, 1.098594, 
    0.9753518, 0.8955016, 0.8678322, 0.9059997, 0.9807558, 0.7565699, 
    0.2632751, 0.2532005, 0.4847107, 0.3372011, -0.02337837, -0.0137105, 
    0.05111647, -0.1188216, -0.2067447, -0.1544991, -0.04294205, 0.1482363, 
    0.3345156, 0.5181408, 0.7771091, 1.024391, 1.195078, 1.303867, 1.337802, 
    1.258539,
  1.437526, 1.330527, 1.245811, 1.18292, 1.177744, 1.208099, 1.195062, 
    1.141335, 1.048448, 0.9855084, 0.9539652, 0.931602, 0.9146585, 0.8818951, 
    0.8434672, 0.7478619, 0.6679463, 0.6549087, 0.5666275, 0.4828711, 
    0.5495529, 0.5567007, 0.4368763, 0.3507252, 0.344264, 0.4013929, 
    0.5170832, 0.5834246, 0.5885353, 0.5762148, 0.5492935, 0.5238543, 
    0.5047302, 0.4337187, 0.3739853, 0.3899679, 0.3272715, 0.2630148, 
    0.2625751, 0.1498957, 0.1406507, 0.1719174, -0.2107649, -0.61096, 
    -0.6646872, -0.5911198, -0.5904522, -0.7682679, -0.9955463, -0.9834538, 
    -0.7560282, -0.580719, -0.5069075, -0.454043, -0.2451236, 0.1193295, 
    0.3990332, 0.5156187, 0.3710872, 0.1520278, 0.004990339, -0.0734272, 
    -0.0031147, 0.1704202, 0.2080181, 0.3462017, 0.6111429, 0.7052348, 
    0.7567325, 0.6591082, 0.3988543, 0.2025657, 0.09817076, 0.07208061, 
    0.140554, 0.1021748, -0.08093023, -0.1539285, -0.07349253, -0.2317443, 
    -0.3761454, -0.2834697, -0.3040915, -0.3945374, -0.3794818, -0.4367085, 
    -0.4418359, -0.2152896, 0.01972008, 0.1729426, 0.3510509, 0.5905204, 
    0.8810649, 1.147943, 1.340212, 1.460084,
  0.9098573, 0.9059834, 0.9177999, 0.9518166, 1.058457, 1.153477, 1.058702, 
    1.017246, 0.9896908, 0.9034605, 0.8492613, 0.8549743, 0.9042091, 
    0.8654075, 0.7539654, 0.5980897, 0.424408, 0.3369079, 0.2723899, 
    0.2100687, 0.178184, 0.07416344, -0.02809906, -0.1510477, -0.3170319, 
    -0.4196835, -0.4679918, -0.4219952, -0.2564354, -0.1909876, -0.2297897, 
    -0.2236223, -0.1832409, -0.1483459, -0.143219, -0.149437, -0.2567778, 
    -0.3174219, -0.2511783, -0.3471904, -0.3935776, -0.4129786, -0.7759175, 
    -1.222109, -1.390826, -1.317145, -1.054043, -0.8879783, -1.090322, 
    -1.353262, -1.318545, -1.087685, -0.8691471, -0.7713768, -0.6744528, 
    -0.5510643, -0.5495346, -0.6418846, -0.7613506, -0.9374251, -0.9227765, 
    -0.8895247, -0.7616758, -0.5101624, -0.4815001, -0.3299215, -0.04984331, 
    0.08995152, 0.2801862, 0.2788672, -0.01353168, -0.251781, -0.4341207, 
    -0.555768, -0.6147685, -0.6900454, -0.6913474, -0.6033916, -0.341152, 
    -0.2526755, -0.4051657, -0.4549377, -0.4615133, -0.4343321, -0.3549705, 
    -0.3424702, -0.2843161, -0.1602926, -0.1270895, -0.08044243, -0.05031538, 
    -0.04396772, 0.09719419, 0.35429, 0.5701108, 0.7751727,
  0.4389586, 0.4444275, 0.5094342, 0.6424417, 0.794281, 0.803998, 0.5547628, 
    0.4153097, 0.2670186, 0.1207294, 0.1174581, 0.1623476, 0.237087, 
    0.2107358, 0.1098897, 0.02958369, -0.09452128, -0.2539124, -0.4713278, 
    -0.6357157, -0.6617739, -0.7136457, -0.8668685, -1.082102, -1.279644, 
    -1.354547, -1.355638, -1.296409, -1.131972, -1.153343, -1.126748, 
    -0.8779359, -0.7268786, -0.6291895, -0.5702209, -0.5447822, -0.56039, 
    -0.5225971, -0.5104878, -0.591738, -0.6422586, -0.6810932, -0.9547095, 
    -1.316624, -1.516868, -1.534658, -1.490745, -1.342991, -1.258112, 
    -1.491543, -1.646247, -1.578392, -1.509902, -1.469619, -1.438727, 
    -1.351585, -1.291039, -1.290355, -1.320498, -1.483844, -1.475218, 
    -1.404955, -1.337848, -1.12359, -0.9921453, -0.8072982, -0.6263411, 
    -0.5696678, -0.3048401, -0.162034, -0.2695699, -0.4320209, -0.6742256, 
    -0.77932, -0.890094, -0.8947003, -0.6274966, -0.3843813, -0.379401, 
    -0.1676821, -0.04632801, -0.05371714, -0.1122786, -0.2101139, -0.2638086, 
    -0.2462144, -0.210325, -0.3302634, -0.4930887, -0.5835834, -0.6347394, 
    -0.5861712, -0.5109434, -0.2716045, 0.01137114, 0.2377377,
  0.08614278, 0.1402278, 0.2376889, 0.3307717, 0.3492775, 0.3383237, 
    0.2597106, 0.07517254, -0.2696189, -0.6170962, -0.5312238, -0.5879459, 
    -0.6792544, -0.5688214, -0.4889549, -0.5721906, -0.671149, -0.785602, 
    -0.9578677, -1.136253, -1.278424, -1.426178, -1.639817, -1.726699, 
    -1.788206, -1.835521, -1.689525, -1.578066, -1.557998, -1.682607, 
    -1.567943, -1.060765, -0.8223532, -0.6533916, -0.5796285, -0.5204, 
    -0.4708068, -0.5237532, -0.5318099, -0.5354395, -0.6529684, -0.9152079, 
    -0.9346251, -0.9390037, -1.179629, -1.314948, -1.449599, -1.591152, 
    -1.647874, -1.873721, -2.054889, -2.100771, -2.177122, -2.101146, 
    -2.002074, -1.839866, -1.51542, -1.342682, -1.233779, -1.244782, 
    -1.293952, -1.309902, -1.293382, -1.161448, -1.094668, -1.098314, 
    -1.194375, -1.14322, -0.8221257, -0.6450262, -0.6042707, -0.7009666, 
    -0.8045799, -0.8056543, -0.9411848, -0.7774315, -0.2519594, -0.04502571, 
    -0.2584862, -0.1631085, -0.01605454, -0.04277974, -0.1638409, -0.3586489, 
    -0.473574, -0.5421125, -0.6135969, -0.8259506, -0.968268, -1.032672, 
    -1.102399, -0.9132552, -0.7957587, -0.6204331, -0.3462954, -0.1699929,
  -0.1685771, -0.08154953, 0.01444674, 0.01029658, 0.04857755, 0.3686134, 
    0.37029, 0.1747658, -0.2500226, -0.8197817, -0.794066, -0.7767801, 
    -0.9895406, -0.7732644, -0.4668517, -0.5845764, -0.7446837, -0.8837299, 
    -0.9953022, -1.044635, -1.106793, -1.146572, -1.19527, -1.122939, 
    -1.13954, -1.355882, -1.430101, -1.4697, -1.473704, -1.592617, -1.473021, 
    -1.020514, -0.9517153, -0.7561749, -0.7515038, -0.6234276, -0.4023826, 
    -0.4657615, -0.6362205, -0.60624, -0.5930402, -1.009642, -1.22442, 
    -1.193024, -1.309251, -1.375527, -1.354857, -1.531956, -1.748851, 
    -1.866722, -1.949404, -1.776602, -1.670921, -1.775137, -1.776162, 
    -1.699746, -1.428164, -1.255182, -1.185179, -1.160342, -1.312279, 
    -1.410244, -1.397907, -1.430198, -1.498053, -1.367064, -1.263157, 
    -1.175153, -0.8785057, -0.5601463, -0.3104393, -0.2552635, -0.3134177, 
    -0.420742, -0.50222, -0.3287823, -0.04457033, 0.1223406, -0.03172815, 
    -0.03810853, 0.0004168749, -0.1393456, -0.2610254, -0.379238, -0.7600486, 
    -0.9555727, -0.7803776, -0.7901103, -0.9861878, -0.8452049, -0.855768, 
    -0.8047426, -0.6785383, -0.5432193, -0.3793195, -0.3415753,
  -0.1914449, -0.04572535, 0.04489946, 0.07821655, 0.311159, 0.5125261, 
    0.3876889, 0.06958961, -0.2901269, -0.8461163, -0.7943094, -0.40082, 
    -0.6539776, -0.5627995, -0.2937236, -0.4462953, -0.4365296, -0.4891829, 
    -0.7258363, -0.874095, -0.8747783, -0.7939839, -0.7934794, -0.8030658, 
    -0.8254132, -0.97193, -1.12346, -1.1982, -1.114508, -1.117682, 
    -0.8456113, -0.5747132, -0.6897523, -0.645823, -0.6906636, -0.6878803, 
    -0.341787, -0.2300847, -0.4116597, -0.5752994, -0.5908266, -0.8174379, 
    -1.034397, -1.156744, -1.127838, -1.091331, -0.9889874, -0.9601786, 
    -1.114785, -1.129449, -1.279905, -1.224843, -1.09802, -1.241917, 
    -1.178945, -1.179303, -1.016136, -0.8023176, -0.8544172, -0.9813215, 
    -1.123639, -1.108112, -1.076308, -1.14099, -1.156533, -0.916966, 
    -0.6975974, -0.661025, -0.4807193, -0.3564026, -0.2610738, -0.1326883, 
    -0.1505597, -0.1463764, -0.1318092, -0.1093489, 0.06830454, 0.05471379, 
    -0.174648, -0.02891266, 0.1790137, -0.08211923, -0.3780661, -0.2477767, 
    -0.6972724, -0.9120504, -0.857265, -0.5661845, -0.7438703, -0.6943419, 
    -0.6495993, -0.6841695, -0.5621154, -0.5381572, -0.4544168, -0.373883,
  -0.001307964, 0.08474302, 0.2211528, 0.4539648, 0.6020607, 0.4431739, 
    0.264235, 0.05569053, -0.09264922, -0.4142805, -0.4407451, 0.08005536, 
    -0.06657541, -0.280573, -0.135911, -0.2453022, -0.3408751, -0.3978906, 
    -0.4683819, -0.5630274, -0.5505104, -0.5386124, -0.5032616, -0.5101309, 
    -0.5482807, -0.6284895, -0.6630759, -0.6186752, -0.4392476, -0.3184633, 
    -0.1951885, -0.3248925, -0.4966369, -0.3277245, -0.4766173, -0.4787173, 
    -0.2302632, -0.0128479, -0.1516988, -0.2521546, -0.3840556, -0.5747786, 
    -0.4666243, -0.5846739, -0.6444886, -0.6157122, -0.5720599, -0.391396, 
    -0.3794169, -0.4194071, -0.5120015, -0.6318419, -0.5933654, -0.4760966, 
    -0.3481994, -0.3815653, -0.2691791, -0.2448142, -0.2436585, -0.3079977, 
    -0.4849508, -0.6248922, -0.7486393, -0.6971903, -0.6769431, -0.6302307, 
    -0.4990296, -0.3983619, -0.2789288, -0.1570044, -0.02056313, 0.1226015, 
    0.1287374, 0.3375268, 0.3170838, 0.3442155, 0.5317806, -0.01115537, 
    -0.3967675, -0.06333637, 0.2211851, -0.2447653, -0.4766824, -0.1993387, 
    -0.4590394, -0.6022363, -0.4782286, -0.3794818, -0.5068421, -0.6090393, 
    -0.5754614, -0.6113667, -0.5648985, -0.5053935, -0.3901429, -0.2076397,
  0.04973364, 0.09100962, 0.1852639, 0.3466572, 0.4576759, 0.1739359, 
    0.147145, 0.1472597, -0.02119756, -0.2618067, -0.4767642, -0.06844711, 
    -0.1133853, -0.2921448, -0.04941988, 0.03239918, -0.1297431, -0.2907782, 
    -0.3543682, -0.4254961, -0.3804102, -0.4177799, -0.4202385, -0.46171, 
    -0.3638906, -0.2632227, -0.1500883, -0.08392572, 0.03695631, 0.1475525, 
    0.09237671, -0.1174703, 0.003851414, 0.002321482, -0.04038668, 
    -0.03678989, -0.03936195, 0.2914, -0.08605766, 0.01949215, 0.1491475, 
    -0.03791285, -0.02415943, -0.09699488, -0.2615781, -0.1849346, 
    -0.1546283, -0.1742249, -0.110146, -0.1091533, -0.08016539, -0.0833559, 
    -0.05360365, 0.08751011, 0.168613, 0.1936951, 0.2218366, 0.03635454, 
    0.09157848, 0.1029396, -0.06885386, -0.1558332, -0.2308493, -0.1355042, 
    -0.2292223, -0.2137103, -0.1110735, 0.03441763, 0.07024145, 0.1872172, 
    0.2461367, 0.3201928, 0.381309, 0.4830995, 0.4711361, 0.6208105, 
    0.3531675, -0.3541079, -0.08498359, 0.09084666, 0.108034, -0.1921284, 
    -0.3034403, 0.07701206, -0.3015695, -0.2623923, 0.08402681, -0.1322494, 
    -0.2154202, -0.259398, -0.3070707, -0.3604722, -0.3788476, -0.2502503, 
    -0.1664777, -0.07251549,
  0.07727242, 0.1684184, 0.2182877, 0.2474709, 0.2859637, -0.00440073, 
    -0.00264287, 0.1512146, -0.00423789, -0.1122296, -0.4578841, -0.3168194, 
    -0.3112855, -0.4223204, -0.1050844, -0.03470659, -0.1040268, -0.1122627, 
    -0.1602602, -0.2755594, -0.2063389, -0.2224684, -0.1785555, -0.183177, 
    0.006991386, 0.09784508, 0.09869099, 0.1840429, 0.2930436, 0.3270931, 
    0.3257751, 0.2594342, 0.2279553, 0.2631941, 0.4732842, 0.2764425, 
    0.1087012, 0.482204, 0.1054301, 0.04865837, 0.2310648, 0.1888285, 
    -0.02020454, -0.04326773, -0.159153, -0.1150937, 0.02849293, 0.02116919, 
    0.03015327, 0.05228901, 0.09852886, 0.2046161, 0.4051208, 0.5317812, 
    0.6322041, 0.4814882, 0.367393, 0.3017516, 0.2727318, 0.2293234, 
    0.1144958, 0.02842808, -0.08342075, -0.05827427, -0.05291939, 0.07022476, 
    -0.008453369, 0.1505632, 0.2370377, 0.356976, 0.378005, 0.4489522, 
    0.4841733, 0.3649187, 0.520062, 0.23834, 0.008571148, -0.3061749, 
    -0.01680321, 0.06052423, 0.006520331, 0.01636708, -0.1443257, 
    -0.01913118, -0.05964184, -0.1031313, 0.2066836, 0.2027926, 0.1041765, 
    0.0233984, -0.03093052, -0.0241766, -0.01354837, 0.02022505, 0.09104204, 
    0.1274028,
  0.1121359, 0.1693294, 0.09831721, 0.270746, 0.4399514, 0.1156673, 
    0.06641603, 0.197943, 0.03072309, -0.01820278, -0.4416404, -0.5184305, 
    -0.3540916, -0.3504128, -0.0762105, -0.02974224, -0.02197838, 0.02453804, 
    0.1122818, 0.02749968, -0.009072304, -0.05337572, -0.033144, -0.0387435, 
    0.03773737, 0.1279235, 0.2177992, 0.3306575, 0.3347273, 0.4626727, 
    0.4759703, 0.2708273, 0.2091246, 0.1415629, 0.327354, 0.4147239, 
    0.238503, 0.0949316, 0.0003845692, -0.02671528, 0.08495474, 0.2312436, 
    0.1739035, 0.1136498, 0.1181092, 0.1442323, 0.1665955, 0.2401142, 
    0.1479921, 0.1250591, 0.1934509, 0.2923603, 0.4151797, 0.4309349, 
    0.5486269, 0.5308852, 0.486794, 0.3716083, 0.1735129, 0.06682301, 
    -0.1292868, -0.1127992, -0.09619808, -0.08097982, -0.1552153, -0.0519433, 
    0.05782223, 0.2316022, 0.2602315, 0.367816, 0.4020934, 0.3426371, 
    0.2721291, 0.1525166, 0.3128517, 0.2263446, 0.04022825, -0.1706116, 
    0.07862321, -0.0355044, -0.1360905, 0.1360123, -0.07723629, -0.1169658, 
    -0.1271877, 0.05725241, 0.1513448, 0.4224219, 0.2947688, 0.2302504, 
    0.2759376, 0.1766863, 0.1254005, 0.07059956, 0.1111593, 0.1804628,
  0.2035096, 0.2062111, 0.05349299, 0.2646911, 0.516156, 0.1657327, 
    0.09994489, 0.222194, 0.02917695, 0.1221132, 0.03972363, -0.2853254, 
    -0.1827371, -0.162441, -0.1326559, -0.1483469, -0.07720327, -0.03885746, 
    0.1523051, 0.1372495, 0.1316671, 0.1434999, 0.1620708, 0.1938252, 
    0.360085, 0.3589292, 0.3159122, 0.4206967, 0.1999614, 0.514854, 
    0.5656676, 0.2438254, 0.04286528, 0.04727554, 0.3260517, 0.428102, 
    0.3246844, -0.05635401, -0.06675422, -0.05542636, -0.06543565, 0.1109476, 
    0.1529393, -0.03172827, -0.3242087, -0.4362206, -0.5626531, -0.4254293, 
    -0.2617574, -0.1399803, 0.04141569, 0.2898703, 0.4790468, 0.6006122, 
    0.6201272, 0.6293235, 0.4627705, 0.2657328, 0.1792579, 0.02271509, 
    -0.1352763, -0.111774, -0.2450585, -0.2093811, -0.15095, -0.04981089, 
    0.06545639, 0.05349302, 0.1972432, 0.2520123, 0.2862077, 0.3576436, 
    0.3969338, 0.3284765, 0.1795346, 0.3608661, -0.08840156, 0.01469091, 
    0.08034846, 0.06760454, 0.04926127, -0.1120342, -0.1459049, -0.02292299, 
    -0.06914687, -0.02422476, 0.04916382, 0.4153256, 0.5623312, 0.44835, 
    0.445518, 0.4401631, 0.2843685, 0.2011008, 0.1629171, 0.2054789,
  0.2195085, 0.1150978, -0.00959301, 0.1450455, 0.0539161, -0.08237922, 
    0.03557307, 0.1442645, 0.1269631, 0.2253516, 0.3974873, -0.1449445, 
    -0.1040265, 0.052256, -0.04100561, -0.1622134, -0.1551981, -0.193691, 
    -0.09857368, 0.02284551, 0.04286504, 0.01625347, 0.08322954, 0.1485777, 
    0.3068297, 0.3109639, 0.155804, 0.1395607, 0.07528681, 0.3136332, 
    0.09929374, 0.04286471, -0.09636053, 0.05806684, 0.2976174, -0.005768061, 
    -0.01154606, -0.04141261, -0.3123922, -0.1317449, -0.3026428, -0.3612692, 
    -0.2930236, -0.08553672, -0.1625388, -0.1085346, 0.03599668, 0.2711203, 
    0.5185163, 0.6846128, 0.7886982, 0.747406, 0.5495219, 0.3814392, 
    0.1722598, 0.06845093, -0.1358461, -0.1236062, -0.204205, -0.2379947, 
    -0.05143833, -0.07918882, -0.1056051, -0.02707291, 0.05619478, 
    0.02261782, 0.05622768, 0.1214294, 0.2425883, 0.2304626, 0.3724871, 
    0.3601335, 0.2564065, 0.2048602, -0.03682256, 0.5357684, 0.04934239, 
    -0.07393214, 0.1202085, 0.2616311, 0.0679462, -0.08226562, -0.1489648, 
    -0.2327538, -0.1560934, 0.02385426, 0.2905536, 0.5626569, 0.8388283, 
    0.7432556, 0.7137635, 0.6901467, 0.3827574, 0.3063579, 0.2520447, 
    0.2844498,
  0.3408303, 0.1341244, 0.04260445, 0.01337242, -0.05363584, -0.1055564, 
    -0.02040024, 0.06171238, 0.07232438, 0.2608336, 0.4759213, -0.142438, 
    -0.1907778, 0.01511431, -0.1372945, -0.2958885, -0.3814679, -0.5009503, 
    -0.5404522, -0.3651268, -0.2520083, -0.1575747, -0.07508761, 0.02707697, 
    0.1496193, 0.3245541, 0.2320902, -0.04704413, 0.001067758, -0.05651677, 
    -0.1265363, 0.009791819, -0.07171859, -0.277741, -0.522158, -0.8825747, 
    -0.8797262, -0.7324281, -0.4060769, -0.04631138, -0.1362534, -0.1615462, 
    0.1360286, 0.4403418, 0.703916, 0.9173601, 0.976068, 1.035589, 1.071869, 
    1.066237, 1.087934, 0.8772726, 0.6873312, 0.4289165, 0.2123961, 
    0.1082134, -0.04198217, -0.1342835, -0.09769535, -0.06156206, -0.2408261, 
    -0.1837139, -0.02529907, -0.1764388, -0.07858658, 0.0658958, 0.07382202, 
    0.07142949, 0.1352313, 0.1937598, 0.2410093, 0.3329852, 0.4896582, 
    0.3123801, -0.1576233, 0.07684928, 0.1012467, -0.007379234, 0.06620458, 
    0.1209246, 0.1647071, 0.03373402, -0.4630924, -0.7594461, -0.6378317, 
    -0.4256897, 0.1186624, 0.5047786, 0.7487237, 0.7829525, 0.7966407, 
    0.7404883, 0.7342384, 0.802663, 0.5015398, 0.4432229,
  0.09761727, 0.1065855, 0.04898453, -0.04878581, -0.1829979, -0.09139645, 
    0.06320989, 0.1260027, 0.2651303, 0.3047463, 0.4184344, 0.1170996, 
    -0.5260153, -0.3963447, -0.2201071, -0.4440651, -0.7496805, -0.8839257, 
    -0.9275291, -0.7362857, -0.4978902, -0.3252182, -0.4313049, -0.4031477, 
    -0.2995017, -0.122972, 0.02971375, 0.01978531, 0.1041768, -0.5514872, 
    -0.764622, -0.30694, -0.4678288, -0.8157616, -1.355687, -1.124469, 
    -1.002252, -0.6661844, -0.2527568, -0.1229231, -0.06019515, 0.3376239, 
    0.583685, 0.2334083, 0.1245378, 0.07837892, -0.2031963, -0.3386128, 
    -0.4592021, -0.5267313, -0.3650777, -0.2391338, -0.07876587, -0.1566956, 
    -0.2228413, -0.3406961, -0.3452697, -0.4457581, -0.3088603, -0.2374897, 
    -0.2535058, 0.1445248, -0.03197265, -0.08421862, 0.1503842, 0.1600198, 
    0.08469416, 0.1181414, 0.1676857, 0.1235449, -0.04728842, 0.1164165, 
    0.1130147, -0.3230855, -0.1561098, 0.04854506, 0.09478521, 0.1975847, 
    -0.07129541, -0.03068662, -0.02974284, -0.2913959, -0.5404358, 
    -0.6604228, -0.2302474, -0.05938137, 0.1613707, 0.5501401, 0.5771257, 
    0.4769789, 0.4477313, 0.4260026, 0.6441669, 0.580251, 0.1325947, 
    0.07077837,
  0.03487313, 0.07745123, -0.01229489, -0.3215392, -0.5707095, -0.2815332, 
    -0.02118158, 0.01465845, 0.1866147, 0.04304376, 0.3395605, 0.1195736, 
    -0.4114807, -0.3931212, -0.2706928, -0.5376205, -1.033714, -1.196393, 
    -1.26887, -0.9991107, -0.4832745, -0.23526, -0.4783583, -0.6056709, 
    -0.4333067, -0.3654523, -0.2008686, 0.1506937, 0.2456319, -0.5668354, 
    -1.24859, -1.474273, -0.7686262, -0.3331932, -1.195791, -0.979173, 
    -0.7510806, -0.4759828, -0.3177635, -0.1101789, 0.1921974, 0.3707131, 
    -0.01613587, -0.5425192, -0.5772687, -0.7733786, -0.922044, -0.9820373, 
    -0.9662821, -0.8803933, -0.6871481, -0.7467673, -0.8475323, -0.9945376, 
    -0.9319396, -0.9640036, -0.9077373, -0.9982975, -0.8756574, -0.7672426, 
    -0.7268456, -0.7237531, -1.080492, -0.8062401, -0.8002018, -0.88985, 
    -0.7835839, -0.7677469, -1.13609, -1.554482, -1.463906, -1.198867, 
    -1.653489, -1.598525, -0.2618716, -0.05077136, -0.1199936, 0.1444271, 
    -0.2765036, -0.3821673, -0.2611222, -0.4020081, -0.3924704, -0.1443261, 
    0.09476888, 0.0719012, 0.1962176, 0.351198, 0.2966084, 0.1907492, 
    0.1728127, 0.2041283, 0.1763773, 0.2236104, 0.1639748, -0.02458334,
  0.07157576, 0.09426451, 0.1326435, 0.1158304, 0.2858827, 0.6451271, 
    0.6136817, 0.300905, 0.2439064, 0.410085, 0.4421325, 0.01115894, 
    -0.2492249, -0.6044824, -0.7015364, -0.5832257, -1.00178, -1.1788, 
    -1.315761, -0.9869208, -0.2732, -0.3643298, -0.919343, -1.034023, 
    -0.5599017, -0.2503486, -0.01385689, -0.006435156, -0.156842, -0.5608459, 
    -1.259576, -1.807558, -1.382265, -0.699209, -0.862718, -0.6022688, 
    -0.4606997, -0.3307031, -0.2237694, -0.06639647, -0.4430238, -0.9099347, 
    -1.210553, -1.054905, -0.8777728, -1.161041, -1.045107, -0.959446, 
    -0.6913476, -0.6460834, -0.6339417, -0.6998758, -0.6566792, -0.523818, 
    -0.4261131, -0.4854064, -0.6101465, -0.7172747, -0.6321187, -0.8202372, 
    -1.294635, -1.749388, -1.833665, -1.700413, -1.820482, -1.798672, 
    -1.80624, -1.624258, -1.663532, -1.360602, -0.5678612, -0.2358787, 
    -0.914606, -1.130296, -0.6931872, -0.7336006, -0.4081268, -0.2802782, 
    -0.196703, -0.1750717, -0.2610087, -0.2114968, -0.1187568, -0.06021118, 
    -0.05969048, 0.04743862, 0.1919372, 0.1763769, 0.1497985, 0.2738708, 
    0.288584, 0.3160257, 0.3380473, 0.2932227, 0.08501959, -0.1256739,
  0.5030375, 0.68917, 0.77667, 0.9493915, 1.400889, 1.567604, 1.185296, 
    0.646836, 0.3630797, 0.4933207, 0.3723409, 0.09924507, -0.1973209, 
    -0.6491112, -0.7921777, -0.2740626, -0.2770567, -0.4621305, -0.6207094, 
    -0.4164438, -0.02095366, -0.4392805, -1.242666, -1.089459, -0.475234, 
    -0.1228089, 0.1185485, -0.2604716, -0.7546451, -1.351325, -1.386367, 
    -0.8787824, -0.9874902, -1.132445, -0.7648013, -0.2547427, 0.0607357, 
    0.1969173, -0.1199447, -0.6330957, -1.269847, -1.480573, -1.280866, 
    -1.105686, -1.142649, -1.200494, -1.006419, -1.104189, -0.9182024, 
    -0.9237852, -0.8318911, -0.667275, -0.4377012, -0.2531309, -0.3365946, 
    -0.4134173, -0.5809145, -0.5345278, -0.5940161, -0.8898335, -0.9914131, 
    -0.9613502, -0.9634502, -1.242047, -1.331761, -1.56931, -1.338597, 
    -0.8073142, -0.9063866, -0.04920883, 0.4577085, 0.1243101, -0.7655985, 
    -0.2604876, 0.01986647, -0.09880257, 0.09288216, -0.08721352, -0.1204329, 
    -0.1771879, -0.1880755, -0.1003804, -0.001291752, 0.03332758, 0.1983013, 
    0.2209578, 0.1713314, 0.2497816, 0.2410583, 0.367393, 0.4322853, 
    0.8648701, 1.105219, 0.4715105, 0.06895506, 0.08218765,
  0.6163186, 0.5320249, 0.4047301, 0.3542418, 0.6256936, 0.6563575, 
    0.4865496, 0.5296484, 0.4385679, 0.2997007, 0.2315367, 0.1748636, 
    -0.003212571, -0.4340884, -0.6648501, -0.3665427, 0.05686235, 
    -0.02391529, -0.2286682, -0.2745352, -0.2521381, -0.56568, -0.6100487, 
    0.05142617, 0.5076921, 0.2902443, -0.03864568, -0.4348208, -0.4078514, 
    -0.5313703, -0.2666731, 0.4258239, 0.2814552, 0.2106382, 0.3096942, 
    0.4289651, 0.4743915, 0.1814227, -0.3753481, -0.9034731, -1.159056, 
    -1.110683, -1.054336, -1.12569, -0.9403706, -0.7874575, -0.8254452, 
    -0.913662, -0.6546936, -0.4916077, -0.2749243, 0.0350523, 0.3129654, 
    0.3010187, 0.1045995, 0.01705074, -0.1051664, -0.08994818, -0.2294655, 
    -0.3210511, -0.2909565, -0.3454485, -0.4171124, -0.553896, -0.5228256, 
    -0.5755922, 0.2521258, 0.3551531, -0.3314191, 0.1865496, 0.309629, 
    -0.7038798, -0.7152567, 0.0274353, 0.2815533, -0.006858349, -0.1519265, 
    -0.2324286, -0.1631408, -0.3206282, -0.1313214, 0.00365591, 0.1186132, 
    0.1620378, 0.1588311, 0.1079369, 0.1156187, 0.2040143, 0.1504173, 
    0.2854595, 0.3406188, 0.6617938, 0.6915138, 0.2093037, 0.2893328, 
    0.5301044,
  0.01115918, -0.1640687, -0.05938101, 0.04641318, 0.03628874, 0.282774, 
    0.6283789, 0.7154395, 0.445469, 0.2458107, 0.3217057, 0.6048279, 
    -0.03205377, -0.3787336, -0.1455792, -0.07422531, -0.08151698, 
    -0.4037657, -0.4650135, -0.420661, -0.4518452, -0.3623762, -0.1323956, 
    0.1779397, 0.2679461, 0.1686623, -0.1500064, -0.3218325, 0.3309996, 
    0.2739354, 0.1907003, 0.2813579, 0.1917416, 0.8262143, 0.9877213, 
    0.9824314, 0.6368263, 0.1260192, -0.02861953, -0.1165266, -0.2883849, 
    -0.3371153, -0.2605042, -0.1825747, 0.02907896, -0.04745102, -0.1312723, 
    -0.03159809, 0.02732134, 0.1096296, 0.1870708, 0.3359632, 0.4381604, 
    0.3440037, 0.243011, 0.1684017, 0.09685183, 0.05966139, 0.04445934, 
    0.08342505, 0.06744146, 0.140049, 0.06947613, -0.0500716, 0.0606707, 
    0.5085225, 1.178005, 0.8413838, 0.08479181, 0.4141213, -0.198818, 
    -0.8710833, -0.3309803, 0.2920189, 0.01854897, -0.2286854, -0.1503325, 
    -0.2440009, -0.2371159, -0.3954816, -0.1666565, -0.08159781, -0.00645113, 
    0.09953785, 0.04719448, 0.1110616, 0.04717779, 0.006634235, 0.05189848, 
    0.1723084, 0.1550722, 0.1667421, 0.05101895, 0.008033991, 0.1055762, 
    0.1209896,
  -0.03202105, -0.0167706, 0.0793395, 0.1446228, 0.07771182, 0.2682065, 
    0.5773374, 0.4692482, 0.1559995, 0.1111264, 0.3336523, 0.09296238, 
    -0.4092023, -0.07116508, 0.7772723, 0.420827, -0.1187889, -0.2837303, 
    -0.3425194, -0.2997948, -0.01209939, 0.1241147, 0.07276416, -0.2006407, 
    -0.01094389, 0.1268328, -0.322679, 0.05704105, 0.716465, 0.4200783, 
    0.3603616, 0.6321551, 0.7891376, 1.094476, 1.140733, 1.008864, 0.7042255, 
    0.6005144, 0.7209573, 0.6582131, 0.5342059, 0.3706484, 0.442409, 
    0.6421328, 0.8107848, 0.714561, 0.5704041, 0.5041442, 0.4925718, 
    0.6962342, 0.8044534, 0.9092546, 0.9272394, 0.8363543, 0.7683201, 
    0.5830989, 0.5215597, 0.4211693, 0.3706317, 0.3695574, 0.4436464, 
    0.5678325, 0.3297298, 0.2365986, 0.4856873, 0.6661558, 1.081976, 
    0.5220965, 0.3848248, 0.37973, -0.203229, -0.2128639, 0.273757, 
    0.5987241, 0.2682067, -0.06222963, -0.2343651, -0.5408105, -0.6403872, 
    -0.6927309, -0.5275614, -0.4113667, -0.2993715, -0.166966, -0.105052, 
    0.02720737, -0.05453062, -0.07754517, -0.1207418, -0.1321025, 0.01863003, 
    0.0699811, 0.1118915, 0.1737078, -0.04512354, -0.1554589,
  0.3056577, 0.2534766, 0.06836963, -0.2603741, -0.1279519, 0.2446061, 
    0.4140397, 0.2746356, 0.04424822, 0.07732081, -0.113662, -0.5854393, 
    -0.4485412, 0.362689, 0.4399838, -0.2392964, -0.3791242, -0.1051332, 
    -0.09660465, 0.08718461, 0.1543882, 0.07860708, -0.1519916, -0.4316795, 
    -0.2535871, -0.4159732, -0.7027082, 0.2394304, 0.9104103, 0.5981054, 
    0.6194599, 0.7790951, 0.8076596, 0.9647563, 1.162299, 1.023025, 
    0.7430766, 0.8858337, 0.8912535, 0.6432068, 0.5573664, 0.5168228, 
    0.6369567, 0.7504654, 0.7649021, 0.7610943, 0.6997986, 0.6734314, 
    0.8307068, 0.964138, 0.9219666, 0.9442809, 0.867018, 0.8294048, 
    0.8232031, 0.7300715, 0.6877217, 0.5038676, 0.3942809, 0.4209247, 
    0.5235779, 0.6460057, 0.5548929, 0.6006124, 0.3929791, 0.4450459, 
    0.6153908, 0.4475521, 0.2594502, -0.01052046, -0.2544663, 0.1035257, 
    0.3883726, 0.5090107, 0.1828224, 0.01101255, 0.1540787, -0.09572589, 
    -0.3065331, -0.3640852, -0.4525942, -0.5749413, -0.5380597, -0.3944073, 
    -0.269521, -0.1588764, -0.1580303, -0.1081929, -0.1079979, -0.1011457, 
    0.0005955696, 0.03724909, 0.1845641, 0.3403255, 0.3931089, 0.3868102,
  0.05393231, -0.2174218, -0.5290917, -0.4667379, -0.1424217, 0.1125422, 
    -0.05016875, -0.3045962, -0.442894, -0.4382391, -0.3649311, -0.2833068, 
    0.06348664, 0.2584574, 0.01810908, -0.1720442, -0.08395827, -0.02088869, 
    0.09512711, 0.3173438, -0.1106021, -0.2626528, -0.1393781, -0.2206444, 
    -0.03358383, 0.008278191, 0.107513, 0.9498633, 1.094541, 0.5496843, 
    0.4957292, 0.5308204, 0.542653, 0.5617775, 0.7353614, 0.5314226, 
    0.2833107, 0.2648375, 0.3607033, 0.2528908, 0.248708, 0.3552184, 
    0.4399675, 0.3248309, 0.1887956, 0.2516537, 0.3558693, 0.4173439, 
    0.576605, 0.7528744, 0.8494889, 0.8764096, 0.8135189, 0.8383723, 
    0.8325621, 0.6462501, 0.485687, 0.3035091, 0.2287369, 0.2100521, 
    0.2455014, 0.4447039, 0.5492125, 0.2950788, 0.243223, 0.3567154, 
    0.5572366, 0.3911721, 0.09574559, -0.236481, -0.1645571, 0.2475848, 
    0.2993426, 0.05521825, -0.1691958, -0.03941059, 0.3673278, 0.3841574, 
    0.276768, 0.1873312, 0.02444053, -0.000803709, 0.05899382, -0.008030534, 
    -0.1395244, -0.1991926, -0.1477929, -0.08293283, -0.05803013, 
    -0.02575493, -0.004775047, 0.1002216, 0.467116, 0.859987, 0.8869077, 
    0.7110127,
  -0.5623107, -0.721344, -1.024941, -0.958584, -0.3562238, -0.3121808, 
    -0.5173078, -0.8506737, -0.8392479, -0.6154847, -0.4472395, -0.1846092, 
    -0.09203076, -0.215631, 0.3248309, 0.4228451, 0.0500102, -0.2352927, 
    0.06924826, 0.2705505, -0.1142318, -0.1718812, -0.01179022, -0.07909164, 
    0.1240982, 0.2289649, 0.1108335, 0.2374448, 0.3074969, 0.2167417, 
    0.2200783, 0.1057391, 0.148366, 0.1396421, 0.04675472, -0.01026026, 
    -0.03443021, -0.05096665, -0.0300031, -0.08423483, 0.01311219, 0.0776304, 
    0.06106114, 0.09325516, 0.1346778, 0.09136724, 0.06016612, 0.1707778, 
    0.3979261, 0.6120538, 0.6021253, 0.4590752, 0.3805763, 0.4024186, 
    0.3465594, 0.194769, 0.1340594, 0.0937764, 0.04664081, -0.01445931, 
    -0.0414452, 0.1018004, 0.2513285, 0.4411559, 0.2256446, 0.09756851, 
    0.01088238, -0.1358626, -0.3725976, -0.5332257, -0.2511457, 0.04237646, 
    -0.06657538, -0.1790102, -0.1663151, -0.1726627, -0.202692, -0.09305668, 
    -0.006369829, -0.06600547, -0.1312561, 0.06070352, 0.1618431, 0.1079853, 
    0.02173877, -0.1733465, -0.2593651, -0.1277734, -0.1191305, -0.1356672, 
    -0.1470441, -0.1785057, 0.09880549, 0.5527119, 0.71889, 0.03278986,
  -0.828213, -0.7263898, -0.9398501, -0.6542544, -0.4229229, -0.3854232, 
    -0.8202049, -1.065696, -0.8862692, -0.482949, -0.2233462, -0.2903383, 
    -0.2206445, 0.1622659, 0.5215429, 0.4521093, 0.09450865, 0.2112404, 
    0.5598569, 0.374424, 0.08000672, 0.07310563, -0.03439763, -0.1659082, 
    -0.01921225, -0.008421183, -0.2110579, -0.1371971, 0.01281917, 
    0.04779637, 0.0667578, 0.07688153, 0.1527116, 0.1112728, -0.07378578, 
    -0.09230775, -0.1733463, -0.2432194, -0.2811749, -0.2602114, -0.3160709, 
    -0.2686751, -0.2605696, -0.1970601, -0.1288147, -0.1807027, -0.1568258, 
    0.00494194, 0.1898379, 0.3204527, 0.3373637, 0.3320904, 0.3417256, 
    0.2606382, 0.09799194, 0.01075244, -0.01929331, -0.09489536, -0.1290751, 
    -0.144114, -0.1661682, -0.07010698, 0.1485941, 0.3035091, -0.01914698, 
    -0.4153058, -0.3897199, -0.2150942, -0.285895, -0.3459697, -0.217324, 
    -0.1160708, -0.051813, 0.1475199, 0.1731706, 0.008424759, -0.1438378, 
    -0.1091211, -0.162034, -0.08395791, 0.105593, 0.2313089, 0.1532328, 
    0.1093853, 0.07671928, -0.06952095, -0.1622784, -0.1344624, -0.2199931, 
    -0.2927797, -0.2719467, -0.3528222, -0.3707584, -0.2404198, -0.4064028, 
    -0.6511295,
  -0.991966, -0.7365299, -0.5354394, -0.4678124, -0.4140526, -0.4612694, 
    -0.3796449, -0.2080303, 0.02305686, 0.07623076, -0.004270673, 0.03425471, 
    0.3190854, 0.5844826, 0.5845802, 0.3747333, 0.2641212, 0.2692319, 
    0.1487077, -0.01592445, -0.03167954, -0.05259424, -0.2204815, -0.2985578, 
    -0.2252017, -0.2549869, -0.3554751, -0.3624085, -0.4459537, -0.4631412, 
    -0.2764876, 0.009319782, 0.1974874, 0.2608011, 0.126263, -0.06950521, 
    -0.222793, -0.3744528, -0.5451397, -0.7290591, -0.9998761, -0.9798241, 
    -0.8558981, -0.704905, -0.5706928, -0.3916731, -0.1695371, -0.03552055, 
    0.08995104, 0.1690855, 0.1186295, 0.109189, 0.1096616, 0.02680016, 
    -0.1527081, -0.3154354, -0.4359603, -0.4301333, -0.3435941, -0.3135638, 
    -0.2805238, -0.0764873, 0.03261113, 0.03985345, -0.2874899, -0.5155988, 
    -0.3751529, -0.243675, -0.2845441, -0.150934, 0.1035256, 0.2684019, 
    0.390342, 0.3360613, 0.2026139, 0.01382816, -0.01372719, -0.02609706, 
    0.05931962, 0.4282002, 0.6893656, 0.8404074, 0.6474223, 0.5368917, 
    0.3501725, 0.142849, -0.02909231, -0.1713438, -0.3501039, -0.4559956, 
    -0.3833394, -0.4058328, -0.5791891, -0.7952378, -1.041168, -1.159739,
  -0.5432026, -0.5294983, -0.4175355, -0.2330139, -0.04998994, 0.107497, 
    0.2442973, 0.4050233, 0.4905537, 0.4853292, 0.4844013, 0.5941182, 
    0.7147889, 0.6595315, 0.4456317, 0.3263936, 0.2732524, 0.08067405, 
    -0.1569726, -0.1992904, -0.1608461, -0.2486066, -0.4101789, -0.5297916, 
    -0.5146223, -0.4108136, -0.3270572, -0.3052146, -0.3409895, -0.2223861, 
    -0.02984047, 0.02684927, 0.02942061, -0.01118803, -0.1292546, -0.3109441, 
    -0.3526269, -0.3554101, -0.4421289, -0.684528, -0.7205627, -0.527643, 
    -0.252887, -0.06569624, -0.01320601, -0.01052046, -0.01421499, 
    -0.03454447, -0.07827806, -0.1734924, -0.242373, -0.216331, -0.1306548, 
    -0.0965066, -0.2228413, -0.364264, -0.4696841, -0.516396, -0.5439677, 
    -0.5086327, -0.2755432, -0.104157, 0.04372728, -0.1937564, -0.4697819, 
    -0.4770736, -0.4213933, -0.3716048, -0.2425195, 0.03222013, 0.1828713, 
    0.1670184, 0.1645933, 0.1939389, 0.1083107, 0.0543555, 0.1284603, 
    0.2663672, 0.4611264, 0.6377703, 0.6395606, 0.7609149, 0.5728455, 
    0.7032979, 0.6608667, 0.4127378, 0.09594107, -0.1790428, -0.2492738, 
    -0.1477113, -0.06750298, -0.007362843, -0.01917982, -0.2288799, 
    -0.4678445, -0.5400288,
  0.07356143, -0.0157125, 0.0004823208, 0.1283305, 0.3509054, 0.5133891, 
    0.5519145, 0.6044698, 0.7185812, 0.8369566, 0.9058043, 0.885801, 
    0.7339621, 0.4846943, 0.2631772, 0.1996193, 0.2181576, 0.1992122, 
    0.1667745, 0.1019633, 0.005543709, -0.05303383, -0.1217675, -0.2109278, 
    -0.3100326, -0.2625227, -0.2073302, -0.2075911, -0.1930077, -0.1194563, 
    -0.0370667, 0.02660477, 0.1356707, 0.1729429, 0.02922547, -0.1998924, 
    -0.3138735, -0.2709862, -0.06934229, 0.0008074343, 0.2041767, 0.3146746, 
    0.3387957, 0.2395769, 0.2842386, 0.2887633, 0.2208436, 0.1538839, 
    0.06145239, -0.02204394, -0.07816362, -0.097646, -0.1839581, -0.3756571, 
    -0.6052794, -0.7276592, -0.7611389, -0.7017479, -0.6585345, -0.5500548, 
    -0.3582096, -0.1234113, -0.1809633, -0.2761133, -0.233242, -0.1218162, 
    0.01542306, 0.1583433, 0.3349056, 0.4242938, 0.3656024, 0.3240987, 
    0.4172951, 0.5171161, 0.5322363, 0.4617773, 0.6986265, 0.9217222, 
    1.023057, 0.9846454, 0.946462, 0.7264423, 0.8983988, 0.9809511, 
    0.9194112, 0.7355571, 0.4272726, 0.1420999, 0.06526041, 0.2060323, 
    0.3862734, 0.5392847, 0.6148205, 0.4531512, 0.2274027, 0.08894253,
  0.3257101, 0.4391704, 0.4930277, 0.6661394, 0.7724385, 0.874717, 0.7553648, 
    0.6830504, 0.6276792, 0.5907651, 0.5916277, 0.5523863, 0.4753844, 
    0.450954, 0.4262794, 0.4137632, 0.3968523, 0.3834571, 0.3179789, 
    0.2123311, 0.1555599, 0.157741, 0.1819922, 0.07673502, -0.05954421, 
    -0.08753908, -0.08817375, -0.1234112, -0.1287824, -0.07241857, 
    0.06141925, 0.1941667, 0.2853776, 0.3175718, 0.1756449, -0.04492823, 
    -0.1771222, -0.1166242, 0.151019, 0.3237891, 0.4266211, 0.3505309, 
    0.3651466, 0.3864683, 0.3799416, 0.504372, 0.6003355, 0.6082782, 
    0.5302347, 0.345355, 0.1531023, -0.09297514, -0.337718, -0.5486394, 
    -0.7369531, -0.8604231, -0.8503482, -0.7254947, -0.5415266, -0.3685935, 
    -0.2504945, -0.2611393, -0.2073467, -0.1040263, 0.06539059, 0.1578549, 
    0.284515, 0.4666438, 0.6356544, 0.6479104, 0.5877216, 0.6812274, 
    0.4877217, 0.6304461, 0.774945, 1.020925, 1.270664, 1.430983, 1.349701, 
    1.181423, 0.868939, 1.048903, 1.093532, 1.041205, 1.024424, 1.03279, 
    0.9589132, 0.7906513, 0.7050233, 0.6987569, 0.6873963, 0.6698017, 
    0.6392841, 0.5194275, 0.3509378, 0.3882098,
  0.3706969, 0.3273699, 0.2918069, 0.3494238, 0.3391376, 0.2803811, 
    0.2396096, 0.2965106, 0.3721617, 0.3879331, 0.3688414, 0.3709735, 
    0.3338642, 0.2615822, 0.2233335, 0.1963804, 0.2166928, 0.2900001, 
    0.2481219, 0.152842, 0.03386414, -0.08386046, -0.1301821, -0.1527733, 
    -0.1177961, 0.01084977, 0.1087827, 0.1326271, 0.1554626, 0.2839129, 
    0.4263444, 0.5181739, 0.4834898, 0.3449482, 0.1458921, 0.00316748, 
    0.006959796, 0.1309671, 0.2295834, 0.2526139, 0.2746354, 0.2859637, 
    0.3693622, 0.5068296, 0.5637631, 0.5021256, 0.3899187, 0.2957944, 
    0.2177019, 0.05341148, -0.1067446, -0.2455304, -0.2324771, -0.2129133, 
    -0.2306216, -0.2571839, -0.2748924, -0.2518293, -0.1800193, -0.03921527, 
    0.08643556, 0.1845963, 0.3010843, 0.3595313, 0.4300393, 0.5084572, 
    0.6263121, 0.8280861, 0.9606219, 0.9202735, 0.7754982, 0.4846454, 
    0.5790627, 0.6552508, 0.7746356, 0.8048764, 1.170388, 1.214512, 
    0.8098896, 0.6678647, 0.6078387, 0.6110125, 0.5401303, 0.4155535, 
    0.3794369, 0.5844174, 0.6591896, 0.7400815, 0.8043557, 0.8459898, 
    0.8423766, 0.8078551, 0.7722757, 0.7497822, 0.6798766, 0.510492,
  0.2919534, 0.3200458, 0.3492286, 0.5032651, 0.4258237, 0.3334735, 
    0.2946063, 0.3161232, 0.3745542, 0.35945, 0.3115822, 0.2875425, 
    0.2914813, 0.310687, 0.2984637, 0.2971942, 0.3085223, 0.3648537, 
    0.3473245, 0.268467, 0.151898, 0.1198993, 0.1617938, 0.2537208, 
    0.3587013, 0.3685158, 0.332855, 0.2759376, 0.2481707, 0.2894305, 
    0.3790789, 0.3899839, 0.3012632, 0.1753517, 0.0685972, 0.008652687, 
    -0.003098786, -0.0003806949, -0.03182602, -0.06978174, -0.07713851, 
    -0.04922511, 0.01001966, 0.07816762, 0.1178485, 0.06626976, 0.03799808, 
    0.0505631, 0.04932618, 0.01661134, -0.01997721, -0.08983397, 0.0212338, 
    0.001849055, -0.03034484, -0.05332667, -0.01774724, 0.06089859, 
    0.2305275, 0.3516538, 0.3756284, 0.4084572, 0.4648048, 0.5255308, 
    0.5986103, 0.6821877, 0.7510028, 0.7589292, 0.6332456, 0.4615985, 
    0.381911, 0.4574806, 0.5703062, 0.6890074, 0.5025327, 0.5587664, 
    0.4947202, 0.5795997, 0.3589292, 0.12973, -0.09168923, -0.09574211, 
    -0.1756899, -0.1824441, -0.2448628, -0.2634664, -0.273314, -0.1521058, 
    0.1222916, 0.3751074, 0.508669, 0.6103126, 0.527728, 0.4881122, 0.439691, 
    0.3545998,
  -0.04526994, 0.05435565, 0.1853777, 0.3238869, 0.4202736, 0.4769468, 
    0.5688576, 0.6247984, 0.6240985, 0.6202248, 0.6413999, 0.619118, 
    0.6074318, 0.5695739, 0.5865172, 0.5290789, 0.5146909, 0.5188739, 
    0.5430437, 0.5517189, 0.5083921, 0.4822853, 0.4863544, 0.492116, 
    0.4797951, 0.3239357, 0.1739194, 0.03352225, -0.06558245, -0.1052472, 
    -0.08659494, -0.06815413, -0.05122703, -0.04149395, -0.1180564, 
    -0.1720442, -0.2926333, -0.3982973, -0.4982322, -0.5370017, -0.5491762, 
    -0.4699607, -0.3252179, -0.1624249, -0.004840314, 0.1216083, 0.2072366, 
    0.2378843, 0.2199643, -0.01120418, -0.02656901, -0.01577795, -0.04769528, 
    0.2331641, 0.2879981, 0.2978126, 0.3052345, 0.3128681, 0.2422951, 
    0.3559344, 0.3779559, 0.3956317, 0.4244403, 0.5227964, 0.6080177, 
    0.6502215, 0.6124936, 0.5448016, 0.4501238, 0.3159767, 0.4929462, 
    0.6224872, 0.6828225, 0.5482521, 0.6255959, 0.3102964, 0.3301369, 
    0.1760353, 0.03764012, -0.08211899, -0.09712553, -0.1093976, -0.2309307, 
    -0.3125876, -0.4198141, -0.3955795, -0.3215233, -0.2009339, -0.07865196, 
    0.03874707, 0.02953482, -0.005881846, -0.04476523, -0.120449, -0.1369204, 
    -0.1176007,
  0.1083272, 0.2801369, 0.4842061, 0.6796811, 0.8504656, 0.9532163, 
    0.9840268, 0.936631, 0.8589779, 0.7733986, 0.6850685, 0.6041279, 
    0.5271258, 0.4294208, 0.3332131, 0.2666115, 0.1670834, 0.1644305, 
    0.1515399, 0.2115985, 0.1219827, 0.02323592, -0.07096994, -0.142731, 
    -0.1951395, -0.2876037, -0.3801333, -0.4527245, -0.4843325, -0.4763085, 
    -0.4359601, -0.3576887, -0.2418846, -0.1393129, -0.1109275, -0.05943036, 
    -0.03879225, -0.09686518, -0.180817, -0.09372425, 0.004811168, 
    0.07045245, 0.13139, 0.1699967, 0.2723243, 0.3426042, 0.3822365, 
    0.4035906, 0.3149678, 0.2444437, 0.09397137, 0.03804684, 0.03036451, 
    0.09568036, 0.1459897, 0.1788999, 0.2194598, 0.2765725, 0.3324157, 
    0.4096616, 0.4780047, 0.5579526, 0.608506, 0.799782, 0.7880308, 
    0.7477476, 0.6558856, 0.5397072, 0.460622, 0.3410582, 0.4792092, 
    0.513926, 0.3800229, 0.4288673, 0.3313413, 0.2203062, 0.1632912, 
    0.0239194, -0.03233051, -0.02738285, -0.01758456, -0.1088767, -0.131826, 
    -0.1138736, -0.06364566, -0.003994003, -0.01177388, -0.03141916, 
    -0.05560541, -0.05628884, -0.1176332, -0.1571027, -0.1361392, 
    -0.09178686, -0.06481749, -0.002138376,
  0.4802507, 0.6031674, 0.6529558, 0.6591733, 0.6429298, 0.5717384, 
    0.5065528, 0.448724, 0.3726662, 0.270355, 0.1687437, 0.07361025, 
    -0.01999313, -0.1005109, -0.2202048, -0.2806052, -0.2959048, -0.318268, 
    -0.4200583, -0.5341372, -0.6063865, -0.6341858, -0.642096, -0.599355, 
    -0.5331607, -0.6120342, -0.4777894, -0.3596256, -0.2307191, -0.07394862, 
    0.02946937, 0.2086849, 0.2680273, 0.2326921, 0.1939714, 0.1976497, 
    0.2163022, 0.3031021, 0.4004167, 0.474961, 0.5735776, 0.6795021, 
    0.7197853, 0.7391049, 0.7278094, 0.6855081, 0.6364031, 0.5712339, 
    0.5298927, 0.5051206, 0.5181903, 0.5539976, 0.5695574, 0.6002541, 
    0.6005145, 0.5968198, 0.5859474, 0.5578387, 0.5359148, 0.5143166, 
    0.4875262, 0.4618263, 0.4740334, 0.5273862, 0.6029721, 0.8062437, 
    0.8271584, 0.8291766, 0.8063413, 0.7707945, 0.7234312, 0.7343524, 
    0.6825783, 0.5755634, 0.5307229, 0.3243589, 0.2253354, 0.1742611, 
    0.1347106, 0.1031678, 0.06791377, 0.05704117, 0.09987962, 0.1238218, 
    0.1201434, 0.06643224, -0.001503825, -0.07196283, -0.1359113, -0.1988672, 
    -0.2109438, -0.1982974, -0.06136703, 0.004827619, 0.140098, 0.328607,
  0.1891212, 0.2365986, 0.2739195, 0.2706644, 0.3102964, 0.2621681, 
    0.2048113, 0.09592463, 0.003265128, -0.03262354, -0.0759341, -0.1351138, 
    -0.1820376, -0.2256899, -0.245384, -0.296035, -0.3014874, -0.341087, 
    -0.38277, -0.4305077, -0.4489648, -0.4284894, -0.3864158, -0.3125063, 
    -0.1910219, -0.1408429, -0.05116189, 0.04472029, 0.1135354, 0.09131855, 
    0.09701514, 0.1706318, 0.2253355, 0.2596617, 0.3023375, 0.3647236, 
    0.4249938, 0.4747496, 0.512624, 0.5455992, 0.5807718, 0.6025979, 
    0.6183694, 0.6115172, 0.5921161, 0.5628517, 0.5309669, 0.4978127, 
    0.4719989, 0.4553647, 0.4519142, 0.4540301, 0.4482033, 0.4401629, 
    0.4378354, 0.4380307, 0.4474221, 0.453965, 0.4512795, 0.4360289, 
    0.4205829, 0.3966083, 0.3813088, 0.3648537, 0.3432555, 0.3400654, 
    0.3239845, 0.314577, 0.2839943, 0.2602475, 0.202549, 0.1830828, 
    0.09795928, 0.1156351, 0.06343782, 0.03671247, 0.01457703, -0.00918591, 
    -0.01540345, -0.04614878, -0.07385075, -0.09666978, -0.1418357, 
    -0.2018619, -0.2787663, -0.3274314, -0.3752017, -0.3801661, -0.3360579, 
    -0.2944564, -0.2291241, -0.1645409, -0.1141991, -0.01721013, 0.07364272, 
    0.1271095,
  -0.1015363, -0.07884751, -0.06774724, -0.0620018, -0.05661444, -0.06921209, 
    -0.06942368, -0.08016586, -0.09308904, -0.1095278, -0.1150942, -0.121686, 
    -0.1458071, -0.174339, -0.203408, -0.2381411, -0.2571841, -0.2590233, 
    -0.2537987, -0.2382062, -0.2116437, -0.1832746, -0.1639875, -0.1225324, 
    -0.08971986, -0.02907535, 0.0009701848, 0.0305438, 0.02927423, 
    0.04112315, 0.06823906, 0.1056252, 0.1386004, 0.1579038, 0.1597267, 
    0.1690529, 0.1876238, 0.2086525, 0.222422, 0.2303647, 0.2285093, 
    0.2171974, 0.1959409, 0.1712013, 0.1423927, 0.112868, 0.08345717, 
    0.05652033, 0.02823257, 0.007741034, -0.02258122, -0.05830714, 
    -0.08127263, -0.09979478, -0.1037336, -0.1014875, -0.1019432, 
    -0.09670231, -0.09730452, -0.1011782, -0.0951561, -0.08849919, 
    -0.07791977, -0.06834947, -0.06688461, -0.07860336, -0.107591, 
    -0.1337303, -0.1502668, -0.1584211, -0.1772687, -0.1829328, -0.1818423, 
    -0.1830467, -0.1722882, -0.2164777, -0.26166, -0.3048404, -0.3211164, 
    -0.3509667, -0.3926657, -0.4332095, -0.4835025, -0.5129296, -0.4703677, 
    -0.4670962, -0.4829816, -0.5302961, -0.5163312, -0.519147, -0.4929263, 
    -0.4261619, -0.3529523, -0.2668032, -0.1856997, -0.1360252,
  -0.2952538, -0.2794497, -0.2605207, -0.2415916, -0.2273664, -0.2193586, 
    -0.2147687, -0.2093163, -0.2031965, -0.1949933, -0.1892153, -0.1823631, 
    -0.1742577, -0.1702049, -0.1609276, -0.160423, -0.1628807, -0.1544172, 
    -0.1470116, -0.1343814, -0.1249738, -0.1190168, -0.1118879, -0.101634, 
    -0.09531886, -0.09351222, -0.09056626, -0.07676417, -0.06704737, 
    -0.05407538, -0.03802718, -0.02692693, -0.01341783, 0.002304837, 
    0.01112644, 0.01674166, 0.02857438, 0.03169939, 0.03479183, 0.03449884, 
    0.03427097, 0.027549, 0.01555353, 0.008408368, -0.0002016723, 
    -0.01395491, -0.02433905, -0.04328436, -0.0598371, -0.07328108, 
    -0.09317043, -0.1074283, -0.1230533, -0.129173, -0.1400617, -0.1574771, 
    -0.1644269, -0.1650942, -0.1626529, -0.1564191, -0.1462954, -0.1406802, 
    -0.139964, -0.1406965, -0.1373436, -0.133535, -0.1301821, -0.124339, 
    -0.122565, -0.1262922, -0.1336001, -0.1391828, -0.1464094, -0.1573143, 
    -0.1755109, -0.1941633, -0.2164451, -0.2433332, -0.2640526, -0.2815331, 
    -0.3006737, -0.311188, -0.3220767, -0.3322818, -0.3368879, -0.3466535, 
    -0.3483136, -0.3518781, -0.3485903, -0.3436913, -0.3543683, -0.351048, 
    -0.3395897, -0.3221092, -0.3105533, -0.3065493,
  -0.4232118, -0.4088886, -0.3925154, -0.3744006, -0.3545761, -0.3325059, 
    -0.3092312, -0.2846869, -0.2597845, -0.2341335, -0.2072453, -0.1801783, 
    -0.1527698, -0.1253123, -0.09800029, -0.07147002, -0.04567242, 
    -0.02103138, 0.001820087, 0.02354956, 0.04348755, 0.06117964, 0.07727623, 
    0.09176254, 0.1058083, 0.1189747, 0.1315074, 0.1427541, 0.1529269, 
    0.1620584, 0.1702127, 0.177146, 0.1829734, 0.187139, 0.1871397, 
    0.1866353, 0.1844699, 0.1803522, 0.1741185, 0.1652642, 0.1540175, 
    0.1402806, 0.1235325, 0.1043595, 0.08241916, 0.05862331, 0.02405405, 
    0.001104593, -0.0261097, -0.0477891, -0.06292486, -0.06626177, 
    -0.1160178, -0.1837916, -0.1749873, -0.2194681, -0.2416687, -0.2623568, 
    -0.2480979, -0.2254252, -0.2536163, -0.3022981, -0.2794137, -0.2938185, 
    -0.2941103, -0.2932634, -0.2983923, -0.3059764, -0.3138208, -0.3041205, 
    -0.3030138, -0.3095241, -0.3165388, -0.2881861, -0.2703309, -0.314342, 
    -0.2696962, -0.328372, -0.3555036, -0.363512, -0.3754902, -0.3888202, 
    -0.4025412, -0.4161968, -0.4287944, -0.4397645, -0.4487815, -0.4563336, 
    -0.4611673, -0.4638042, -0.4641948, -0.4635611, -0.458499, -0.4528022, 
    -0.4462585, -0.4353867,
  -0.6781113, -0.6454943, -0.5956733, -0.5378444, -0.4759467, -0.4133978, 
    -0.3537461, -0.3010443, -0.2563503, -0.2185573, -0.1843776, -0.1511745, 
    -0.1188666, -0.0903998, -0.06779242, -0.05237913, -0.04477823, 
    -0.04292238, -0.04428983, -0.0467968, -0.05136943, -0.05851436, 
    -0.07042837, -0.09276009, -0.1285014, -0.1820655, -0.2433772, -0.3062196, 
    -0.3684926, -0.4272647, -0.4822297, -0.5288591, -0.5604835, -0.576076, 
    -0.573081, -0.5491719, -0.504365, -0.4428091, -0.3692241, -0.2881043, 
    -0.2011261, -0.1158391, -0.02252865, -0.02269149, 0.009144664, 
    0.03805089, 0.03704214, 0.03437304, 0.03028774, 0.01476026, -0.02028179, 
    -0.06356049, -0.02905464, -0.04192972, 0.03464866, -0.0964222, 
    -0.08624983, -0.07604504, -0.07060862, -0.06419611, -0.07461119, 
    -0.07885933, -0.09471369, -0.1081729, -0.1420436, -0.1956563, -0.2319031, 
    -0.265123, -0.2697781, -0.2520371, -0.229446, -0.2044948, -0.1727403, 
    -0.1592311, -0.1207871, -0.1320664, -0.09707296, -0.08125281, 
    -0.03126907, -0.04349232, -0.02540898, 0.0282526, -0.01766157, 
    0.001479149, 0.03839254, 0.007338524, -0.0879097, -0.1698594, -0.258759, 
    -0.3551126, -0.4496441, -0.534996, -0.6000834, -0.655015, -0.6863956, 
    -0.6930529,
  -0.6476752, -0.6728218, -0.6409857, -0.5923366, -0.537584, -0.4902207, 
    -0.455211, -0.4270371, -0.398375, -0.366295, -0.3291531, -0.296894, 
    -0.2718775, -0.2587428, -0.2573752, -0.2677753, -0.2897973, -0.3292665, 
    -0.3795762, -0.4291363, -0.4656277, -0.4662292, -0.4009956, -0.3025743, 
    -0.2425157, -0.2449571, -0.2718937, -0.2989935, -0.3309922, -0.3817086, 
    -0.4495957, -0.5366883, -0.6490583, -0.7833519, -0.9061232, -0.9871922, 
    -1.016668, -0.9966316, -0.9268723, -0.8105974, -0.6714048, -0.477313, 
    -0.2333026, -0.0902853, 0.0165664, 0.06025124, 0.07768297, 0.06961, 
    0.03876689, -0.0162624, -0.08138285, -0.1369655, -0.1601914, -0.1465196, 
    -0.1030788, -0.06281197, -0.03349864, 0.003447771, 0.04514718, 0.1029269, 
    0.1535616, 0.1684868, 0.1401827, 0.08927131, 0.03694391, -0.009198606, 
    -0.05512968, -0.1027207, -0.1383002, -0.1629584, -0.1824734, -0.1931829, 
    -0.1949081, -0.1614447, -0.139114, -0.1166693, -0.09642193, -0.10692, 
    -0.0739122, -0.03816998, -0.005048156, 0.02931058, 0.08752966, 0.1216605, 
    0.2067683, 0.2470515, 0.2704732, 0.2640605, 0.2182264, 0.1906714, 
    0.0180316, -0.1239114, -0.2772641, -0.4172225, -0.5238302, -0.606106,
  -0.0207057, -0.1167498, -0.2110863, -0.3004251, -0.3814149, -0.4258809, 
    -0.4364445, -0.4322456, -0.4172392, -0.3912625, -0.3652858, -0.3501817, 
    -0.3419135, -0.3316758, -0.3281927, -0.3373724, -0.3687853, -0.4794133, 
    -0.6574571, -0.801599, -0.7865419, -0.7897801, -0.7661967, -0.6487002, 
    -0.4649605, -0.3421088, -0.2952662, -0.2536323, -0.2138046, -0.1949895, 
    -0.2028673, -0.2196966, -0.2450709, -0.2781115, -0.3249538, -0.4254582, 
    -0.5829773, -0.7403507, -0.8276877, -0.8488951, -0.8067083, -0.7124043, 
    -0.5149107, -0.2633815, -0.1005554, 0.0116837, 0.002373457, 0.09198952, 
    0.08975971, 0.06946349, 0.02569735, -0.0342637, -0.1156114, -0.145071, 
    -0.1452338, -0.1168159, -0.01842725, -0.1071479, -0.08706379, 
    -0.03133345, 0.004734278, 0.07945752, 0.1163716, 0.1755672, 0.1925592, 
    0.2152152, 0.2212868, 0.207387, 0.1661925, 0.1120911, 0.06269264, 
    0.01217175, -0.04749632, -0.09298706, -0.08877206, -0.1370144, 
    -0.1670926, -0.1683457, -0.1987494, -0.2672064, -0.2069688, -0.1438178, 
    -0.09993756, -0.02225208, 0.08419335, 0.1836725, 0.25169, 0.2987769, 
    0.3739071, 0.5173643, 0.5813131, 0.6123028, 0.5353007, 0.4012351, 
    0.2455549, 0.09672546,
  -0.08489799, -0.004917622, 0.02249146, 0.06323051, 0.04078579, -0.08125305, 
    -0.2077012, -0.2806511, -0.3298526, -0.2759786, -0.2370625, -0.1895523, 
    -0.1538434, -0.1561542, -0.1715198, -0.1109076, -0.08411741, -0.05055594, 
    -0.01123311, -0.01712513, -0.1158714, -0.1371441, -0.1767273, -0.2395048, 
    -0.333384, -0.4197288, -0.4160018, -0.3801289, -0.3600931, -0.3707867, 
    -0.3731306, -0.3544292, -0.3369167, -0.3294785, -0.3020537, -0.2786648, 
    -0.2580429, -0.2349637, -0.2184272, -0.2480983, -0.3089054, -0.3276551, 
    -0.2889993, -0.1975932, -0.1136098, 0.02742267, 0.051934, 0.2098931, 
    0.3164198, 0.3732229, 0.3875133, 0.3735485, 0.3019342, 0.2176406, 
    0.1509252, 0.1128879, 0.1075006, 0.1147271, 0.187302, 0.2747858, 
    0.3613743, 0.4367813, 0.5369927, 0.6926244, 0.8226862, 0.9065237, 
    0.9662081, 0.9793428, 0.9829562, 0.9391572, 0.7367814, 0.5371389, 
    0.4322882, 0.3287077, 0.2767551, 0.3535941, 0.290248, 0.2573217, 
    0.1966933, 0.1664362, 0.08546285, 0.1339004, 0.1540338, 0.1916641, 
    0.1899876, 0.1536269, 0.1186335, 0.09867895, 0.09348702, 0.1011531, 
    0.1253562, 0.09807754, 0.08429146, 0.09597778, -0.005032063, -0.04656744,
  -0.037503, 0.06158638, -0.1611185, -0.02752471, 0.0281229, 0.1478169, 
    0.1210592, -0.02363539, -0.09697533, -0.1777527, -0.2810404, -0.3526063, 
    -0.3727069, -0.2695656, -0.2217793, -0.1665871, 0.01264393, -0.01129824, 
    -0.04450142, 0.00592196, -0.06183505, 0.02615309, 0.2058887, 0.4336243, 
    0.413703, 0.3500309, 0.2730618, 0.2088842, 0.1194963, 0.03204632, 
    -0.05335426, -0.06466675, -0.05481958, -0.04240131, -0.0396843, 
    -0.05644751, -0.09936762, -0.1122417, -0.1197128, -0.01562738, 
    0.07288218, 0.1268046, 0.1578093, 0.1655898, 0.1289688, 0.142608, 
    0.1996393, 0.250746, 0.3457167, 0.4468888, 0.5518855, 0.6352352, 
    0.7217419, 0.8003393, 0.8321915, 0.8102188, 0.7382631, 0.6715956, 
    0.6626928, 0.6882141, 0.7148581, 0.7357564, 0.763849, 0.8010721, 
    0.8473611, 0.8876934, 0.9444315, 0.9978496, 1.042462, 1.06559, 0.9907686, 
    0.835251, 0.5919406, 0.3964166, 0.282175, 0.2754043, 0.3840957, 
    0.5071751, 0.5229628, 0.4898086, 0.3347955, 0.3708632, 0.4375787, 
    0.5300592, 0.5502577, 0.4913222, 0.3874323, 0.2431777, 0.1122207, 
    0.09128968, 0.07421613, 0.07000059, 0.09926486, 0.08228886, 0.05312252, 
    0.01021862,
  0.5719862, 0.5689752, 0.5077448, 0.460821, 0.420782, 0.4196099, 0.4651016, 
    0.5052546, 0.4907038, 0.4195449, 0.341013, 0.2746881, 0.1748996, 
    0.0487442, -0.03696561, -0.04363847, 0.06611073, 0.1019994, 0.0873509, 
    0.05273172, 0.09555399, 0.2381646, 0.4098933, 0.5238581, 0.5708632, 
    0.593715, 0.6755508, 0.7038387, 0.6561333, 0.592006, 0.6405895, 
    0.7392552, 0.8076968, 0.6585097, 0.6426082, 0.5850887, 0.5400696, 
    0.5112281, 0.5312955, 0.5380177, 0.5468724, 0.5439258, 0.5550756, 
    0.5742325, 0.6181452, 0.6375462, 0.6588189, 0.7220515, 0.8354305, 
    1.039972, 1.165672, 1.321954, 1.417462, 1.538409, 1.583868, 1.566794, 
    1.466306, 1.35252, 1.276886, 1.20182, 1.13421, 1.062497, 1.028074, 
    1.024786, 1.012855, 0.9842091, 1.030889, 1.100991, 1.124038, 1.154018, 
    1.253725, 1.24212, 1.003725, 0.7205873, 0.4005837, 0.2562635, 0.247865, 
    0.2602348, 0.2832329, 0.3370903, 0.323077, 0.3179011, 0.3617811, 
    0.4755185, 0.6403458, 0.7776016, 0.8557761, 0.847345, 0.7364233, 
    0.6102512, 0.4762669, 0.4158012, 0.4185356, 0.4547009, 0.4937472, 
    0.5559055,
  0.9557271, 0.9923971, 1.001072, 0.956362, 0.8678691, 0.7709126, 0.7259581, 
    0.7054341, 0.7148907, 0.7619283, 0.8192201, 0.9099908, 0.9879365, 
    0.9609998, 0.892087, 0.8296845, 0.8149387, 0.8537084, 0.9332498, 
    0.9347146, 0.9019186, 0.8181295, 0.7681127, 0.8481913, 1.040558, 1.27687, 
    1.496759, 1.665264, 1.747296, 1.849868, 2.066892, 2.310788, 2.540622, 
    2.734372, 2.936553, 2.868487, 2.434307, 2.424476, 2.473256, 2.471124, 
    2.348484, 2.220799, 2.245099, 2.55672, 2.844138, 3.021514, 2.998826, 
    2.760235, 2.500274, 2.379864, 2.279766, 2.250615, 1.954895, 1.897817, 
    1.704571, 1.641078, 1.704049, 1.670276, 1.863669, 1.912791, 1.907696, 
    1.994627, 2.058282, 2.123044, 2.196465, 2.302553, 2.375664, 2.281279, 
    2.061325, 1.85003, 1.765915, 1.833591, 2.014467, 2.094105, 1.945309, 
    1.778008, 1.608818, 1.673304, 1.707955, 1.692998, 1.604376, 1.304278, 
    0.9765766, 0.920229, 0.9810691, 1.086521, 1.25488, 1.404685, 1.471596, 
    1.448646, 1.323338, 1.152439, 1.021189, 0.9492977, 0.9028947, 0.9155085,
  1.395766, 1.389337, 1.361781, 1.431655, 1.514793, 1.45117, 1.428155, 
    1.430498, 1.621222, 1.719316, 1.766176, 1.928545, 2.265395, 2.550795, 
    2.793813, 2.903025, 2.950925, 2.969106, 2.966176, 2.690216, 1.95208, 
    1.50776, 1.346807, 1.375436, 1.692282, 2.086586, 2.484991, 2.705059, 
    2.910967, 3.03644, 3.225828, 3.313751, 3.458884, 3.51074, 3.492559, 
    3.439043, 3.464759, 3.457501, 3.36821, 3.307907, 3.331116, 3.392787, 
    3.532077, 3.619122, 3.617201, 3.602325, 3.458054, 3.181443, 2.856508, 
    2.734616, 2.762139, 2.731117, 2.612546, 2.531394, 2.544838, 2.55667, 
    2.543764, 2.589272, 2.63032, 2.55283, 2.360415, 2.140834, 2.059861, 
    2.134486, 2.201593, 2.201055, 2.20628, 2.23364, 2.213344, 2.139597, 
    2.033884, 1.944724, 1.899965, 1.89741, 1.970473, 2.058266, 2.02337, 
    1.854929, 1.704392, 1.691421, 1.763654, 1.769936, 1.749281, 1.860707, 
    1.740231, 1.587757, 1.512904, 1.613441, 1.761227, 1.7735, 1.696351, 
    1.652048, 1.637269, 1.541908, 1.479327, 1.392722,
  2.672377, 2.799363, 2.644838, 2.469968, 2.338361, 2.248533, 2.09754, 
    1.940053, 1.875275, 1.725421, 1.605532, 1.544561, 1.577211, 1.635839, 
    1.754784, 1.923354, 2.008884, 2.041746, 2.232259, 2.545637, 2.980027, 
    2.91201, 2.695848, 2.29803, 2.097298, 2.161816, 2.350097, 2.453417, 
    2.4687, 2.500421, 2.550161, 2.569773, 2.620554, 2.724152, 2.749233, 
    2.745376, 2.807664, 2.941355, 3.107859, 3.235805, 3.328741, 3.336993, 
    3.304815, 3.280173, 3.236228, 3.150778, 2.985479, 2.718617, 2.428464, 
    2.304473, 2.360463, 2.422816, 2.380727, 2.273874, 2.17031, 2.091811, 
    2.054392, 1.977878, 1.924607, 1.916111, 1.905808, 1.847524, 1.743227, 
    1.70309, 1.772296, 1.85418, 1.896417, 1.943471, 2.004603, 2.075518, 
    2.160349, 2.169301, 2.039874, 1.913718, 1.954148, 1.959894, 1.746727, 
    1.478155, 1.34915, 1.412547, 1.631623, 1.777277, 1.80545, 1.686489, 
    1.752276, 1.902586, 2.124152, 2.35397, 2.63351, 2.864289, 3.077977, 
    3.173777, 3.091225, 2.874021, 2.654767, 2.542104,
  2.396775, 2.400893, 2.305401, 2.19339, 2.155483, 2.125356, 2.04147, 
    1.897101, 1.734861, 1.527114, 1.354327, 1.270066, 1.187042, 1.059779, 
    0.9735661, 0.9546366, 0.9732733, 1.033545, 1.061995, 1.07259, 1.165119, 
    1.244579, 1.228662, 1.170475, 1.096418, 1.076252, 1.223615, 1.413997, 
    1.458413, 1.429556, 1.439777, 1.411766, 1.444823, 1.63758, 1.809455, 
    1.85073, 1.827147, 1.775796, 1.758657, 1.905304, 2.130531, 2.188637, 
    2.137384, 2.13045, 2.158933, 2.119138, 1.977797, 1.832175, 1.657483, 
    1.486585, 1.414612, 1.520391, 1.638701, 1.579749, 1.391615, 1.224998, 
    1.121905, 1.112611, 1.06507, 0.9968076, 1.031589, 1.149151, 1.16904, 
    1.044495, 0.9126916, 0.8924608, 0.9567676, 1.03958, 1.128138, 1.267233, 
    1.560463, 1.821498, 1.873744, 1.838393, 1.793276, 1.599492, 1.238491, 
    1.307907, 1.477211, 1.567365, 1.500876, 1.560072, 1.675421, 1.642104, 
    1.606687, 1.644269, 1.697964, 1.693634, 1.687498, 1.760577, 1.867332, 
    2.000128, 2.132012, 2.207257, 2.244839, 2.316713,
  1.929018, 1.865786, 1.770994, 1.665233, 1.618081, 1.591779, 1.522459, 
    1.369773, 1.143943, 0.9349427, 0.7559872, 0.6383276, 0.5906391, 
    0.5779114, 0.6039696, 0.5924301, 0.5500793, 0.5821438, 0.5937157, 
    0.5640936, 0.6471024, 0.6437817, 0.4498682, 0.373127, 0.435709, 
    0.4161777, 0.4351711, 0.5876455, 0.703742, 0.7596827, 0.8342438, 
    0.8605947, 0.8479319, 0.8206377, 0.7220364, 0.5946922, 0.5194969, 
    0.4484358, 0.3596497, 0.3701315, 0.5610652, 0.7071433, 0.6049299, 
    0.4754047, 0.5343394, 0.5299287, 0.4449525, 0.4196911, 0.4248028, 
    0.3559711, 0.3012671, 0.4029758, 0.5594051, 0.5901992, 0.5447726, 
    0.4229953, 0.315834, 0.3162897, 0.3153458, 0.1226048, -0.04643822, 
    -0.0825057, -0.01172161, 0.1201963, 0.2135725, 0.3190575, 0.3840957, 
    0.3316221, 0.2777162, 0.3187804, 0.4543924, 0.6730447, 0.8003554, 
    0.8682423, 0.9446583, 0.7927876, 0.4515605, 0.5840955, 0.704505, 
    0.636147, 0.5408502, 0.7665019, 1.033364, 1.082062, 1.065021, 1.012628, 
    0.9954896, 1.007289, 1.016973, 1.070604, 1.163084, 1.310577, 1.499705, 
    1.687563, 1.822377, 1.925486,
  1.094057, 1.169383, 1.209031, 1.188442, 1.179262, 1.214321, 1.172296, 
    0.9867654, 0.7583952, 0.6986461, 0.7161269, 0.6042295, 0.4253073, 
    0.3211718, 0.2873015, 0.2919087, 0.335073, 0.4580388, 0.5068498, 
    0.4194813, 0.3943176, 0.3329887, 0.07805729, -0.2056332, -0.35464, 
    -0.3528662, -0.309165, -0.2369156, -0.1097832, -0.0746603, -0.1593285, 
    -0.2707214, -0.3477564, -0.4682474, -0.5891457, -0.6238632, -0.7618341, 
    -0.9704447, -0.9813175, -0.9252949, -0.8736677, -0.7757511, -0.8280792, 
    -0.8831077, -0.8021669, -0.7272482, -0.7102892, -0.7678576, -0.8898628, 
    -0.8397162, -0.6896021, -0.5924013, -0.4544621, -0.3335962, -0.2417994, 
    -0.1965847, -0.2280624, -0.2324076, -0.2706237, -0.4203961, -0.5005717, 
    -0.5573263, -0.6477237, -0.6954942, -0.6949077, -0.5970564, -0.5089698, 
    -0.5181174, -0.443882, -0.3295426, -0.261167, -0.1209493, 0.02228022, 
    0.02634907, -0.01635981, -0.09305191, -0.1998072, -0.2382181, -0.202395, 
    -0.2023301, -0.1603541, 0.06430435, 0.1614561, 0.1466126, 0.1597471, 
    0.1612449, 0.2774234, 0.5039029, 0.7191715, 0.8606586, 0.8887677, 
    0.8858376, 0.9288068, 0.9139466, 0.9312639, 1.014533,
  0.5424786, 0.5629702, 0.5624003, 0.5164356, 0.6154108, 0.7842412, 
    0.9145799, 0.9826465, 0.8573871, 0.7071919, 0.670017, 0.5407853, 
    0.3501763, 0.1841774, 0.1001611, 0.09848404, 0.1080213, 0.1696424, 
    0.2313457, 0.1765757, 0.00733757, -0.2655458, -0.4790554, -0.6690292, 
    -0.9957867, -1.21719, -1.401922, -1.590399, -1.533823, -1.490399, 
    -1.612746, -1.746275, -1.844078, -1.861184, -1.86999, -1.758564, 
    -1.720494, -1.796291, -1.677737, -1.5459, -1.575523, -1.575442, 
    -1.733889, -1.878501, -1.878306, -1.868134, -1.751516, -1.630521, 
    -1.799189, -1.902444, -1.713073, -1.487926, -1.156514, -0.8718295, 
    -0.8589549, -0.9037628, -0.9237981, -0.8676291, -0.8286967, -0.925946, 
    -0.8953471, -0.8528504, -0.9518735, -1.072382, -1.226418, -1.201939, 
    -1.043719, -0.9478536, -0.8614764, -0.8391132, -0.8410993, -0.7807641, 
    -0.7554383, -0.7781925, -0.783906, -0.7452493, -0.6331568, -0.5852571, 
    -0.4996934, -0.4877636, -0.6385611, -0.7423693, -0.7101433, -0.5646193, 
    -0.416491, -0.2335641, 0.0395813, 0.2764785, 0.4127259, 0.4821582, 
    0.5019169, 0.4837546, 0.4379201, 0.3578916, 0.343504, 0.4628234,
  -0.07410717, -0.04368782, 0.01715231, 0.004229784, 0.02252412, 0.01765704, 
    -0.04098582, 0.117836, 0.1690893, 0.007126331, -0.02028251, 0.01453185, 
    -0.05441332, -0.1936064, -0.3278511, -0.4238951, -0.4703796, -0.4747903, 
    -0.5182965, -0.6392763, -0.7520528, -1.013316, -1.369256, -1.552264, 
    -1.7584, -1.960288, -2.214194, -2.38309, -2.376776, -2.611818, -2.67951, 
    -2.558465, -2.548471, -2.338771, -2.196356, -2.082684, -1.7862, 
    -1.356351, -1.196064, -1.40015, -1.54455, -1.739357, -2.278062, 
    -2.641588, -2.618004, -2.547073, -2.572903, -2.455162, -2.41138, 
    -2.500149, -2.395674, -2.280488, -2.104902, -1.758482, -1.532571, 
    -1.365416, -1.32497, -1.269029, -1.136233, -1.228339, -1.392727, 
    -1.364211, -1.212193, -1.033759, -0.9988625, -0.9553244, -0.9045267, 
    -0.9304557, -0.9976587, -1.132718, -1.16631, -1.194598, -1.255373, 
    -1.162242, -1.074449, -0.8963566, -0.5424343, -0.2878444, -0.5062689, 
    -0.443655, -0.4105658, -0.6071316, -0.7479356, -0.761233, -0.6632351, 
    -0.3591825, -0.1984401, -0.2325714, -0.2007833, -0.1515484, -0.04454994, 
    0.04379702, 0.008168697, -0.07207298, -0.1875191, -0.1803246,
  -0.9590195, -0.9678903, -0.836884, -0.7528183, -0.5209498, -0.1511582, 
    -0.04432231, -0.09907496, -0.1816921, -0.3320339, -0.3453151, -0.3499375, 
    -0.4407908, -0.4626818, -0.5589707, -0.8192735, -0.9994329, -1.101988, 
    -1.165676, -1.323701, -1.407539, -1.396764, -1.644143, -1.918085, 
    -2.171894, -2.277753, -2.321699, -2.402705, -2.43669, -2.742548, 
    -2.467011, -1.766783, -1.64385, -1.302298, -1.101353, -0.9698106, 
    -0.8953639, -0.9316757, -0.9315782, -1.110435, -1.211445, -1.592158, 
    -2.021487, -2.249514, -2.498343, -2.569518, -2.674742, -2.743378, 
    -2.615448, -2.683596, -2.674482, -2.582441, -2.57497, -2.386542, 
    -2.12082, -1.825849, -1.499498, -1.254771, -1.119892, -1.16221, 
    -1.159817, -1.107489, -1.062242, -0.9558296, -0.9201851, -0.9127307, 
    -0.9277046, -0.9943225, -1.102265, -1.221324, -1.220592, -1.218655, 
    -1.179283, -1.154934, -1.20373, -0.9404972, -0.3938666, -0.04013936, 
    -0.4334987, -0.3866724, -0.2637885, -0.366702, -0.5185902, -0.7532091, 
    -0.9300973, -0.5296901, -0.2287787, -0.3636094, -0.4299179, -0.6354842, 
    -0.8660675, -0.9488959, -1.049433, -0.938463, -0.9751489, -1.039732,
  -1.131318, -1.098978, -0.9842314, -0.882782, -0.5535184, -0.06919211, 
    0.2495091, 0.1817031, -0.1414252, -0.2829781, -0.2002954, -0.2109728, 
    -0.4979999, -0.5436387, -0.4013529, -0.6851587, -0.9322124, -1.203811, 
    -1.305699, -1.196096, -1.186883, -1.143166, -1.174693, -1.254592, 
    -1.442206, -1.560174, -1.553762, -1.662584, -1.62069, -1.713121, 
    -1.420283, -1.040774, -1.128551, -0.9371449, -0.9272975, -0.7499538, 
    -0.5285996, -0.6920925, -0.8529326, -0.8913115, -0.8734728, -1.263772, 
    -1.614423, -1.607457, -1.864147, -1.958743, -1.90303, -1.976191, 
    -1.989375, -1.973034, -2.001988, -1.898343, -1.901272, -1.97873, 
    -1.815335, -1.589212, -1.284182, -1.043329, -1.030943, -0.9535182, 
    -0.8049181, -0.7527045, -0.8228053, -0.7775905, -0.7070339, -0.6261094, 
    -0.6049994, -0.7321152, -0.8503932, -0.9551621, -1.047301, -1.063317, 
    -1.047285, -0.977005, -0.7518259, -0.4406928, -0.1883978, 0.2040665, 
    0.05973041, -0.1833684, -0.1119818, -0.2584662, -0.3717314, -0.4057806, 
    -0.9146184, -1.096585, -0.7431016, -0.8639838, -1.169664, -1.321324, 
    -1.381871, -1.335159, -1.394746, -1.313772, -1.266995, -1.241051,
  -0.7950382, -0.6707058, -0.4742858, -0.257961, -0.06619734, -0.09409446, 
    0.01650119, 0.07128644, -0.1464057, -0.5163434, -0.2368348, 0.1125298, 
    -0.3319681, -0.5529494, -0.3813992, -0.6677604, -0.8429222, -0.9577184, 
    -1.074352, -0.9545112, -0.7673855, -0.635664, -0.6360869, -0.6537781, 
    -0.6998234, -0.8105173, -0.826158, -0.911037, -0.7625515, -0.7056661, 
    -0.4640975, -0.3544621, -0.5998065, -0.5156109, -0.6910343, -0.7153993, 
    -0.3516468, -0.3204781, -0.4975286, -0.7551459, -0.7533711, -0.8449895, 
    -1.044029, -1.0119, -0.8992701, -0.8367045, -0.7843771, -0.7351744, 
    -0.8240743, -0.9022319, -1.141555, -1.285321, -1.297171, -1.38415, 
    -1.1876, -1.08747, -1.037893, -0.8691106, -0.7936218, -0.7215031, 
    -0.7659531, -0.6967149, -0.6296576, -0.5465198, -0.4765328, -0.425426, 
    -0.4005886, -0.4696803, -0.4357121, -0.4980814, -0.5614278, -0.5279319, 
    -0.5991564, -0.5260763, -0.3210635, -0.02640247, 0.09280324, 0.2284479, 
    0.1419895, -0.04883075, 0.1356419, 0.05180407, -0.2787786, -0.3834822, 
    -1.249579, -1.679104, -1.510288, -1.270494, -1.531285, -1.495413, 
    -1.45718, -1.368785, -1.277802, -1.21068, -1.050556, -0.8969264,
  -0.1808128, -0.004412651, 0.2363098, 0.4425104, 0.3139296, -0.0349474, 
    -0.1265326, -0.1334984, -0.05517769, -0.3632026, -0.2137554, 0.4228327, 
    0.1156549, -0.2551947, -0.2034369, -0.3208528, -0.4958515, -0.6193709, 
    -0.6461287, -0.6488142, -0.5096865, -0.3168478, -0.1908226, -0.1655455, 
    -0.1448421, -0.2205749, -0.1993999, -0.1901073, 0.005384922, 0.1055803, 
    0.2472637, 0.1758926, -0.1919942, -0.3135767, -0.5110378, -0.5389023, 
    -0.3298523, -0.2024441, -0.2468939, -0.3713403, -0.4796252, -0.5108433, 
    -0.2744498, -0.3119335, -0.2630239, -0.1453314, -0.1413927, 0.03115034, 
    -0.05040932, -0.2409201, -0.4218774, -0.5467629, -0.4588079, -0.4285669, 
    -0.434638, -0.5277524, -0.4584985, -0.3008487, -0.2961934, -0.2422714, 
    -0.2108748, -0.1714869, -0.1904812, -0.08045483, -0.02876186, 
    -0.05553627, -0.02428675, -0.07710218, -0.141295, -0.1933293, -0.1728215, 
    -0.1180201, -0.1330113, 0.1408019, 0.1935363, 0.5006485, 0.5811821, 
    0.1662409, -0.03206635, -0.05773383, 0.009632796, 0.05509162, 0.08541393, 
    -0.128778, -0.7060566, -1.30552, -1.199905, -1.071959, -1.23651, 
    -1.156969, -1.095462, -0.9935246, -0.7762232, -0.6240749, -0.4043818, 
    -0.2815623,
  0.2667947, 0.287693, 0.3678685, 0.508526, 0.2543105, -0.1743191, 
    -0.2491565, -0.1463726, -0.003403664, -0.230422, -0.2827988, 0.2686823, 
    0.1728002, -0.1523137, -0.2105331, -0.3235044, -0.3804216, -0.4712105, 
    -0.3872576, -0.2476578, -0.05153179, 0.06054401, 0.1250305, 0.09278774, 
    0.1077452, 0.03915882, 0.1119452, 0.1885061, 0.3219857, 0.371726, 
    0.3545556, 0.2756815, 0.1684871, -0.02301693, -0.1062846, -0.0654974, 
    -0.1211934, 0.2181616, -0.06030464, -0.02444839, 0.03795338, 0.002699852, 
    0.1688285, 0.125421, 0.04745913, 0.1541476, 0.1371069, 0.08603191, 
    0.1396627, 0.04451275, 0.01783657, -0.0760603, -0.08271694, -0.105227, 
    -0.1142926, -0.04962826, 0.06589937, 0.0897603, 0.05344868, 0.1765604, 
    0.3279271, 0.2880683, 0.1701474, 0.2458315, 0.1958642, 0.1674623, 
    0.1784163, 0.2136536, 0.1779428, 0.2256327, 0.1854801, 0.1975565, 
    0.2066059, 0.3397765, 0.3253074, 0.4260717, 0.3294082, -0.06522077, 
    0.02206767, -0.05690372, -0.1445013, -0.1306341, -0.006073475, 
    0.02307749, -0.4555688, -0.7167501, -0.6915874, -0.6834655, -0.6980648, 
    -0.6370788, -0.5526714, -0.4576845, -0.2782736, -0.09738255, 0.03790474, 
    0.1089001,
  0.349997, 0.2599902, 0.2372369, 0.5049289, 0.5324518, 0.1322238, 
    -0.08066678, 0.07828569, -0.03105664, -0.1333029, -0.2603705, 0.1296363, 
    0.1327772, -0.1111679, 0.01562309, -0.1492863, -0.171031, -0.1677437, 
    -0.1110697, -0.0004739761, 0.1563625, 0.2096004, 0.257452, 0.2642069, 
    0.3422661, 0.2827454, 0.2940569, 0.3599262, 0.3729138, 0.3790021, 
    0.4041967, 0.3883278, 0.5003066, 0.4947557, 0.5073702, 0.3174777, 
    0.1833315, 0.566339, 0.190671, -0.1287613, -0.02176428, 0.06375027, 
    0.07312489, 0.1769834, 0.1182909, 0.01952934, -0.01432467, 0.02955532, 
    0.251121, 0.2460418, 0.1996236, 0.1323538, 0.2088513, 0.2316375, 
    0.2423797, 0.2700329, 0.2993627, 0.3463511, 0.3274059, 0.2957664, 
    0.2728982, 0.2516732, 0.1568332, 0.1931124, 0.1998839, 0.3770962, 
    0.2889628, 0.3882127, 0.346694, 0.3752084, 0.3407683, 0.4475226, 
    0.5163879, 0.4017391, 0.4512181, 0.1388646, 0.02994528, -0.01378846, 
    0.01353905, 0.05011129, -0.0264512, -0.03011322, -0.04105067, 0.08858824, 
    -0.2675972, -0.3795104, -0.2143736, -0.1728535, -0.2206402, -0.247642, 
    -0.1565776, -0.07858276, 0.07112408, 0.1827445, 0.2729626, 0.2809873,
  0.2218239, 0.2099584, 0.04584697, 0.1049132, 0.3924127, 0.3654271, 
    0.2384902, 0.4399869, 0.3003724, 0.002504349, -0.2962584, -0.06050014, 
    0.0907526, -0.151792, 0.0125947, -0.08929253, -0.08751822, -0.1513042, 
    -0.02539253, 0.1359029, 0.2554502, 0.2409811, 0.2606754, 0.3218889, 
    0.372117, 0.3553529, 0.4171205, 0.5188618, 0.4206519, 0.3847303, 
    0.3507299, 0.154995, 0.1666155, 0.1702616, 0.3952451, 0.6260066, 
    0.4211402, 0.2233052, 0.06038094, -0.03411651, -0.08247328, -0.1692238, 
    -0.03058529, 0.08124685, 0.1439257, 0.1149387, 0.1219044, 0.1924944, 
    0.1737108, 0.0231576, -0.004039764, -0.07220268, 0.09905386, 0.2787089, 
    0.3792949, 0.3890595, 0.417933, 0.3938608, 0.2529273, 0.1910462, 
    0.1269188, 0.1097636, 0.009388924, 0.1478658, 0.1702776, 0.3127418, 
    0.3088031, 0.4507141, 0.4242973, 0.5526338, 0.5489402, 0.4536929, 
    0.4199357, 0.2726212, 0.24697, 0.1570286, 0.05820051, -0.04536402, 
    0.108054, 0.1750787, -0.01133084, -0.02373314, 0.06614304, -0.0895853, 
    -0.2195821, -0.1704125, -0.0483582, 0.03453445, 0.0001120567, 
    -0.03224516, 0.06060934, 0.06793308, 0.1812315, 0.1683736, 0.2242656, 
    0.1817689,
  0.2020317, 0.2371718, 0.05278051, 0.05689907, 0.2391739, 0.2201959, 
    -0.04347594, 0.3829076, 0.4425919, 0.1680317, -0.06155825, -0.2161484, 
    0.1572406, 0.01446676, -0.130259, -0.2542663, -0.1549821, -0.1527858, 
    0.06677818, 0.08528376, 0.2699032, 0.3819966, 0.4431295, 0.5401673, 
    0.6404443, 0.6111636, 0.628921, 0.6047506, 0.1741669, 0.2203259, 
    0.2899714, 0.2147107, 0.05322075, -0.0662291, 0.2248514, 0.3985171, 
    0.2387832, -0.05060485, -0.03091085, 0.04791415, 0.03726959, -0.1759462, 
    -0.2396345, -0.4427433, -0.4907901, -0.4564481, -0.5674019, -0.4246278, 
    -0.1585641, -0.05688715, 0.1466608, 0.305532, 0.5216126, 0.6155906, 
    0.6098285, 0.6215625, 0.4783673, 0.3514466, 0.3165007, 0.308558, 
    0.2527637, 0.2100716, 0.1253223, 0.2137666, 0.2158995, 0.3056936, 
    0.4222307, 0.4450827, 0.4507957, 0.4711885, 0.4248023, 0.5125957, 
    0.5160615, 0.3692844, 0.1171361, 0.1761042, -0.08512634, -0.04948181, 
    -0.04557556, 0.2293268, 0.432582, -0.1440945, -0.05869389, -0.03987885, 
    -0.04762554, -0.09049654, -0.08878779, 0.1383443, 0.2175422, 0.00868845, 
    0.01420593, -0.006512642, 0.08808374, 0.102797, 0.18172, 0.1679168,
  0.2151666, 0.1787896, -0.03183889, 0.09325886, 0.09989953, -0.004820347, 
    -0.07506774, 0.07117249, 0.1916803, 0.3532848, 0.2082174, -0.2287951, 
    0.1382951, 0.03419316, -0.1578965, -0.2691915, -0.3325384, -0.3791685, 
    -0.03300977, 0.1043274, 0.2135072, 0.2912414, 0.4356101, 0.5337543, 
    0.6853333, 0.5972636, 0.3309056, 0.209405, 0.02097714, 0.2295706, 
    0.04609111, 0.04594463, -0.1227403, -0.2538439, 0.0247044, -0.01886657, 
    -0.03123637, -0.08076436, -0.1603384, 0.08414507, -0.07047725, 
    -0.2500834, -0.2785833, -0.4083035, -0.2926946, 0.01845503, 0.2883279, 
    0.6736305, 0.9552226, 0.9087377, 0.7570138, 0.6556945, 0.6326466, 
    0.5711722, 0.4645486, 0.4649396, 0.4021788, 0.3628874, 0.2659473, 
    0.3330216, 0.4613266, 0.3759418, 0.2918758, 0.221108, 0.347312, 
    0.2633438, 0.2214003, 0.2461729, 0.3516908, 0.4056942, 0.4367323, 
    0.4256647, 0.1716608, 0.1113905, 0.001722693, 0.4553361, -0.04983991, 
    -0.08799092, -0.100084, 0.2615533, 0.4720514, -0.08056903, -0.1943713, 
    -0.1938179, -0.01954985, -0.0324564, 0.2075491, 0.4100409, 0.3752093, 
    0.1557274, 0.2162409, 0.1209614, 0.08832788, 0.06775403, 0.1798151, 
    0.3034804,
  0.3685031, 0.2659323, 0.04449677, 0.06983769, 0.05733782, -0.0256536, 
    -0.004901722, -0.02482361, 0.0996393, 0.3783991, 0.352227, -0.2310736, 
    -0.07962504, 0.02924526, -0.1083196, -0.3758816, -0.4747097, -0.6146185, 
    -0.5029975, -0.2692249, -0.1703313, -0.0441758, 0.1806614, 0.2432591, 
    0.3131321, 0.3335911, 0.1331352, -0.02972269, -0.1603054, -0.2125189, 
    -0.3144394, -0.002964878, -0.04739847, -0.4145371, -0.7958684, 
    -0.9621283, -0.8135606, -0.6891134, -0.3077011, 0.027879, -0.1141142, 
    -0.1078476, 0.1696589, 0.1659155, 0.4328586, 0.8498509, 1.212709, 
    1.486391, 1.565867, 1.440785, 1.26437, 1.12228, 0.9966607, 0.728806, 
    0.5979462, 0.5576472, 0.4991188, 0.3921852, 0.3642397, 0.4629374, 
    0.4537082, 0.3336234, 0.3596988, 0.2800763, 0.3104308, 0.2150698, 
    0.2211723, 0.177976, 0.1003064, 0.1686009, 0.1999811, 0.1808079, 
    0.2686986, 0.2825332, -0.1575384, -0.01979446, -0.1308946, 0.00383848, 
    -0.0594753, 0.1646133, 0.336114, 0.06487358, -0.5150416, -0.471633, 
    -0.2459493, -0.07179642, 0.2153134, 0.3463359, 0.495343, 0.3440237, 
    0.2779107, 0.2075818, 0.3051242, 0.4259902, 0.4146783, 0.5026013,
  0.1379366, 0.09557033, -0.01702738, 0.004212976, -0.006708503, -0.09241784, 
    -0.02687436, 0.04083383, 0.2645482, 0.3557755, 0.4079401, 0.08464909, 
    -0.5521021, -0.2598822, -0.1395044, -0.4284205, -0.5585638, -0.774791, 
    -0.7959498, -0.5498235, -0.328306, -0.1388204, -0.1333518, -0.1644559, 
    -0.1748564, -0.1386093, 0.01809645, -0.1051296, -0.2369817, -0.7813823, 
    -0.9638529, -0.4663438, -0.6765978, -0.8769557, -1.648879, -1.541669, 
    -1.081399, -0.7084336, -0.3311062, -0.3052437, -0.3075221, -0.2529974, 
    0.01046282, -0.07636988, -0.3422391, -0.2944686, -0.08874011, 0.04117584, 
    0.05868936, 0.1840475, 0.3407044, 0.5185201, 0.6423972, 0.5003562, 
    0.4766419, 0.5151348, 0.5666158, 0.497442, 0.5024219, 0.3266573, 
    0.3406222, 0.4736627, 0.3987766, 0.247442, 0.03591859, 0.03707418, 
    -0.1121446, -0.273603, -0.2349476, -0.100996, -0.04389858, -0.05729389, 
    -0.03633022, -0.2507186, 0.0917623, 0.03739968, -0.1330923, 0.4094374, 
    -0.01691345, -0.1290229, -0.0239284, -0.01784086, -0.4797726, -0.6325378, 
    -0.1052918, 0.04680729, -0.02033138, 0.03407943, 0.3292291, 0.2770318, 
    0.3513646, 0.3931124, 0.40239, 0.4137506, 0.1095188, 0.05501032,
  -0.08079684, -0.2056017, -0.1544459, 0.03053117, 0.2494929, 0.2613906, 
    0.2154433, 0.2450984, 0.2632298, 0.1881484, 0.4797986, -0.02915311, 
    -0.4911973, -0.3087924, -0.2465191, -0.4734559, -0.8531103, -0.8875997, 
    -0.8383811, -0.5896664, -0.03558159, 0.03980923, -0.2277365, -0.2473006, 
    -0.2237983, -0.2158222, -0.2022972, -0.2581563, -0.2569361, -0.5987492, 
    -0.8569522, -1.308743, -1.027395, -0.4872097, -1.305455, -1.187389, 
    -1.004788, -0.8548204, -0.5725938, -0.6554877, -0.6154811, -0.7084174, 
    -0.6686876, -0.5750514, -0.6009306, -0.2154162, -0.0472188, -0.2674663, 
    -0.4268086, -0.401597, -0.1220398, 0.06957793, 0.1879699, 0.07839966, 
    0.09646606, 0.1058407, 0.1113741, -0.1313503, -0.3207386, -0.4354194, 
    -0.06645773, 0.07385796, -0.1432805, -0.3342798, -0.7307644, -0.6050155, 
    -0.92261, -1.028844, -1.038495, -1.376288, -1.612388, -1.652119, 
    -1.861852, -2.109215, -0.3996446, -0.1474147, -0.3651067, 0.2619758, 
    -0.4645691, -0.6033068, -0.07532787, -0.04414272, -0.4635286, -0.2991071, 
    -0.2229676, -0.1542339, -0.1066107, -0.01386976, 0.1661595, 0.1759089, 
    0.1393862, 0.1060691, -0.05763531, 0.1159484, -0.02122641, -0.1573105,
  0.09141982, 0.1135389, 0.3648901, 0.440134, 0.3821262, 0.1200332, 0.107875, 
    0.06078838, 0.1702935, 0.5447409, 0.6026338, -0.1657904, -0.1730495, 
    -0.1603379, -0.1796575, -0.1635447, -0.6848826, -0.6377134, -0.6044946, 
    -0.1997576, 0.2776661, -0.09775591, -0.4808292, -0.4211292, -0.1040225, 
    0.0153451, -0.04207659, -0.04664993, 0.05460334, 0.05269921, -0.161705, 
    -0.8929219, -0.9400742, -0.60692, -1.018508, -0.9199573, -1.010387, 
    -1.070282, -0.9190779, -1.119436, -1.391034, -1.534606, -1.318102, 
    -0.8296416, -0.4837754, -0.2763367, -0.4629738, -0.5726426, -0.2557154, 
    0.08079243, 0.5482402, 0.6973782, 0.5900536, 0.4076481, 0.4062805, 
    0.412221, 0.2028131, -0.174367, -0.2320006, -0.1103058, 0.07797551, 
    -0.1938829, -0.4088405, -0.6518419, -0.9714381, -1.100149, -1.670527, 
    -1.680048, -1.706318, -1.881106, -1.786608, -1.506611, -1.022757, 
    -1.481789, -1.581661, -1.30757, -0.8031101, -0.4866552, -0.5385599, 
    -0.3467636, -0.2370625, -0.2344594, -0.2824407, -0.2026715, -0.1645699, 
    -0.009361267, 0.0232563, 0.111326, 0.1656058, 0.1096653, -0.06818283, 
    0.1441224, 0.2458308, 0.2362117, 0.1404595, -0.01333272,
  0.3067356, 0.2111953, 0.2496555, 0.1785619, 0.07724333, -0.09839106, 
    0.1699362, 0.413002, 0.4514459, 0.5522758, 0.4893526, 0.2533827, 
    0.1081678, -0.08821905, -0.3248562, 0.05908012, 0.1084943, -0.07348824, 
    0.09646606, 0.4498343, 0.2029924, -0.5110695, -0.7532907, -0.350556, 
    0.2663224, 0.1954076, 0.09949279, 0.1902155, 0.2849583, 0.3264295, 
    0.1548477, -0.135403, -0.2995632, -0.216995, -0.3886585, -0.5773791, 
    -0.9849798, -1.251109, -1.36745, -1.541409, -1.704674, -1.33192, 
    -0.6129253, -0.1914253, -0.3042827, -0.677525, -0.7482285, -0.5443392, 
    -0.2114615, 0.04820728, 0.2462378, 0.1717257, 0.149168, 0.1795554, 
    0.1990213, 0.1575985, 0.03393316, -0.01881742, 0.1111798, 0.1483045, 
    -0.1265483, -0.6516297, -1.041848, -1.305569, -1.386982, -1.618557, 
    -1.628258, -1.302135, -1.213577, -0.3143907, 0.1394668, -0.07448179, 
    -0.6821316, -0.635777, -0.3425641, -0.296649, 0.03194809, -0.002313614, 
    -0.01364136, -0.02752447, -0.1074891, -0.08156157, -0.003078461, 
    0.02799273, 0.1463838, 0.1820455, 0.1969376, 0.4578753, 0.4392715, 
    0.4946756, 0.5236626, 0.977797, 0.8092585, 0.1665013, 0.1851536, 0.2510878,
  0.1094211, -0.4601092, -0.5724792, -0.2443542, -0.006577969, 0.3693337, 
    0.7175102, 0.8264459, 0.9996718, 0.7108047, 0.8628556, 0.7150202, 
    0.02314162, -0.2497911, -0.8409857, -0.5809761, 0.1319311, -0.04054594, 
    0.0940733, 0.1782036, -0.1376486, -0.2906113, -0.131155, 0.4770646, 
    0.4655898, 0.1025039, 0.009372368, -0.08961856, -0.001353502, 0.0113256, 
    0.1163874, 0.5046849, 0.9568007, 0.8061824, 0.02851295, -0.6331733, 
    -1.101679, -1.151289, -1.003388, -0.8498071, -0.6510112, -0.03600502, 
    0.3585587, 0.03476286, -0.2549834, -0.4639668, -0.3578796, -0.1976595, 
    -0.1378937, -0.05067062, -0.1016297, -0.140449, -0.01775932, 0.1007948, 
    0.01529694, -0.09484339, -0.06411457, 0.01902342, 0.04674196, 0.01510239, 
    -0.2320504, -0.5541205, -0.8263204, -1.039228, -1.001663, -0.7674507, 
    -0.06740174, -0.05965433, -0.3984564, 0.06578529, 0.09016657, -0.5681016, 
    -1.12536, -0.3004413, 0.4762678, 0.3109179, 0.1654439, 0.1647592, 
    0.1411276, -0.0638051, 0.02890301, -0.01943636, 0.02786255, 0.09083462, 
    0.06156921, 0.1018686, 0.2041965, 0.3170052, 0.3679824, 0.6249003, 
    0.6585755, 0.8098282, 0.3076797, -0.08667278, 0.05059969, 0.210414,
  -0.5038757, -0.9815938, -0.9004579, -0.5604024, -0.5257838, 0.1969218, 
    0.6480768, 0.7189916, 1.061976, 0.8629856, 1.067331, 0.8642877, 
    -0.1347846, -0.1042346, -0.2638209, -0.1978705, 0.1146294, -0.0997417, 
    0.0328424, 0.02628326, -0.05770129, -0.06150973, 0.2914525, 0.3914525, 
    0.1407851, 0.1127415, -0.09972595, -0.4142116, -0.01556182, 0.1211398, 
    0.1742818, 0.2307265, 0.3243788, 0.3974102, 0.1000955, -0.01512241, 
    -0.1398787, 0.06236768, 0.3112285, 0.3572569, 0.509552, 0.7509584, 
    0.643568, 0.1251774, 0.005075932, -0.05322456, -0.08986235, -0.03302574, 
    -0.1067739, -0.1469908, -0.2151399, -0.1736851, -0.1482449, -0.1391954, 
    -0.08735657, -0.05403948, -0.006838799, 0.001234531, 0.09537554, 
    0.1482401, 0.04954195, -0.01971245, -0.1890004, -0.3054553, -0.1200548, 
    0.3236302, 0.7626113, 0.4288711, 0.006556511, 0.2760553, -0.2595081, 
    -0.9193549, -0.5460639, 0.558217, 0.7159805, 0.5543275, 0.6318984, 
    0.5512505, 0.4698539, 0.247426, 0.1888642, 0.0463686, 0.1282525, 
    0.2170715, 0.1737123, 0.1942201, 0.09915066, 0.145391, 0.2562957, 
    0.3815732, 0.3476539, 0.327472, -0.04201126, -0.176289, -0.3819851, 
    -0.4612167,
  -0.6061385, -0.8101094, -0.7770691, -0.5287786, -0.3695011, 0.1792618, 
    0.5143366, 0.5052058, 0.7218887, 0.5155734, 0.4486465, 0.09322649, 
    -0.4063015, 0.04220128, 0.1676731, -0.006513059, 0.05684957, 0.02618551, 
    0.1243626, 0.2681125, 0.1863253, -0.1137071, -0.02671158, -0.0952332, 
    -0.112177, -0.06741801, -0.3389837, 0.04361701, 0.5114875, 0.1954889, 
    0.1982565, 0.2143035, 0.07006621, 0.156476, 0.216876, 0.4752908, 
    0.8027968, 1.026691, 0.8485653, 0.7776995, 1.006102, 0.9785786, 
    0.8531876, 0.6326962, 0.5186334, 0.3691545, 0.3169413, 0.1990862, 
    -0.1141133, -0.2142272, -0.2286973, -0.2304549, -0.1814156, -0.04248285, 
    0.07491589, 0.09137201, 0.134356, 0.1366997, 0.2397437, 0.2788057, 
    0.2733867, 0.2813451, 0.1224258, 0.1355117, 0.4704733, 0.6137023, 
    0.7602186, 0.322735, 0.182843, 0.09316182, -0.01989174, -0.02602768, 
    0.2309709, 0.6510234, 0.4776008, 0.5408502, 0.6705215, 0.4737434, 
    0.4336231, 0.2278779, 0.09111023, 0.04749036, 0.02958727, 0.02791119, 
    0.1156554, 0.1936331, 0.1084123, 0.1192846, -0.02422142, -0.07007074, 
    -0.04931831, -0.2006855, -0.1589708, -0.07998312, -0.2649278, -0.5024602,
  0.05099016, 0.01547599, -0.09642196, -0.2407739, -0.1133971, 0.0992322, 
    0.3388483, 0.604929, 0.5853164, 0.193666, 0.1361302, 0.05987692, 
    -0.01577425, 0.1027805, -0.05976832, -0.1975286, 0.03443742, 
    -0.006854892, -0.04842386, 0.2076795, 0.186179, -0.1551778, -0.2828801, 
    -0.4152532, -0.5157909, -0.6686218, -0.6382675, 0.2888973, 0.3609016, 
    -0.0070014, 0.03507233, -0.1137395, -0.2788439, -0.09448433, 0.06726694, 
    0.6364238, 1.091892, 1.261652, 1.12451, 1.1388, 1.199526, 1.013523, 
    0.9633117, 0.9156556, 0.8358052, 0.665004, 0.4445286, 0.1951146, 
    -0.0868845, -0.2240098, -0.31177, -0.3461127, -0.2773299, -0.1362169, 
    0.03919029, 0.1425431, 0.2301245, 0.2929018, 0.3282857, 0.2405577, 
    0.1882131, 0.2704239, 0.3075495, 0.382664, 0.3924782, 0.4162407, 
    0.1308405, 0.05020881, 0.08853865, -0.2603054, -0.271292, 0.03870165, 
    0.2342584, 0.3829076, 0.2715632, 0.2601534, 0.194268, 0.04905343, 
    0.01262766, -0.1002305, -0.1293646, -0.1394395, -0.1352403, -0.002004504, 
    0.1077285, 0.07356524, -0.03135014, -0.1181178, -0.326272, -0.4924011, 
    -0.6615741, -0.7077985, -0.4739604, -0.2427924, 0.03630921, 0.1004367,
  -0.3843777, -0.3787302, -0.2368357, 0.02376044, 0.4548315, 0.5834121, 
    0.7155569, 0.7185355, 0.1400039, -0.2359401, 0.01726627, 0.1572078, 
    -0.0990749, -0.2275256, -0.3311224, -0.3287787, -0.1090521, -0.07708585, 
    -0.00150001, 0.1611789, -0.07871389, -0.1279486, -0.08416605, -0.1251165, 
    0.04096413, 0.1374974, 0.3322728, 0.5775855, 0.1874161, -0.05241156, 
    -0.01924086, -0.2852728, -0.2743679, -0.1002141, 0.01044643, 0.2405734, 
    0.213116, 0.2335098, 0.6252254, 0.8989718, 0.8547009, 0.7190729, 
    0.7338028, 0.7638158, 0.7634739, 0.707289, 0.5147271, 0.2321263, 
    -0.08450776, -0.339, -0.4467311, -0.4057807, -0.3545437, -0.2674831, 
    -0.0791693, 0.04034567, 0.06082094, 0.1248834, 0.1796198, 0.1088679, 
    0.07859421, 0.1845677, 0.3210747, 0.2388639, 0.2939425, 0.2585748, 
    0.1895481, 0.1973444, 0.2625299, -0.07352152, -0.2397325, 0.01117903, 
    0.08391666, 0.08197969, 0.1264134, 0.1433079, 0.1774225, 0.1398411, 
    0.002764225, -0.160517, -0.1501164, -0.07376564, 0.02426493, 0.04286849, 
    -0.133629, -0.296959, -0.3610866, -0.4086452, -0.5213081, -0.6169951, 
    -0.726077, -0.7002958, -0.6118356, -0.4666857, 0.02310938, 0.0347631,
  -0.6378446, -0.7362003, -0.5041367, -0.2144883, 0.281589, 0.4193335, 
    0.2260064, -0.1470404, -0.3934271, -0.3271999, -0.2901556, -0.5874375, 
    -0.7983588, -0.6046574, -0.1147001, -0.3207873, -0.4016955, -0.1062689, 
    0.0366022, -0.1547064, -0.2861354, -0.09285736, 0.008395731, 0.03175192, 
    0.1529922, 0.1828263, 0.200681, 0.1228164, -0.1339056, -0.2247585, 
    -0.3292507, -0.446959, -0.2500514, -0.1462917, -0.148017, -0.1578478, 
    -0.1913764, -0.03515889, 0.1329076, 0.3489557, 0.5572727, 0.639304, 
    0.5506322, 0.4334606, 0.3156059, 0.1044734, -0.08331895, -0.2021503, 
    -0.2977078, -0.2781439, -0.1903834, -0.1990421, -0.2458353, -0.2210312, 
    -0.1661489, -0.1172225, 0.02856183, 0.1657852, 0.1422338, 0.03180075, 
    0.008672506, 0.05318755, 0.1789362, 0.2709122, 0.1544244, 0.2092422, 
    0.207289, 0.1511205, -0.1852076, -0.4626166, -0.3036159, 0.06054424, 
    0.1189264, 0.08225656, 0.1022598, 0.1358533, 0.2495579, 0.4499648, 
    0.4607074, 0.3197246, 0.234812, 0.2629371, 0.2613907, 0.1201146, 
    -0.1028841, -0.3294628, -0.5056505, -0.5266469, -0.5059925, -0.4111844, 
    -0.2634953, -0.277444, -0.2858261, 0.06003964, 0.4006484, -0.08561461,
  -0.4263211, -0.2489121, -0.1593615, -0.1178412, 0.01487367, 0.04960674, 
    -0.1336614, -0.3472846, -0.2376003, 0.008688748, -0.09681252, -0.4830593, 
    -0.6307806, -0.1864935, -0.03052026, -0.2517606, -0.2964871, 
    -0.002720729, 0.03157289, -0.1558946, -0.1623887, -0.08265236, 
    -0.06250262, -0.03494728, 0.007061243, -0.053388, -0.1311551, -0.2055691, 
    -0.2826523, -0.3837593, -0.5261743, -0.616132, -0.4482937, -0.2777698, 
    -0.1733916, 0.04111052, 0.2158827, 0.4324028, 0.3592584, 0.1929497, 
    0.2902154, 0.2786919, 0.1198385, 0.04205537, -0.1082869, -0.2739439, 
    -0.2946143, -0.2749534, -0.1868844, 0.002503395, 0.09208727, 0.1241999, 
    0.1533184, 0.1268859, 0.07929468, 0.06200886, 0.1234679, 0.1412091, 
    0.1172993, 0.06461382, -0.0653348, -0.1777207, -0.01805294, 0.1651341, 
    0.1201634, -0.05429951, -0.1516466, -0.2669458, -0.395136, -0.4285346, 
    -0.3089707, -0.1766301, -0.06242144, 0.09768605, 0.128334, 0.1905899, 
    0.2144506, 0.2446265, 0.1866841, 0.3052545, 0.4305801, 0.4704075, 
    0.3901832, 0.2650368, 0.1899066, 0.05878687, -0.03608608, 0.04939556, 
    0.1542137, 0.1852684, 0.1900532, 0.08139396, 0.03917408, 0.1698377, 
    0.1858697, -0.1497097,
  -0.001695514, -0.01284432, 0.1556773, 0.2014459, 0.04399151, -0.07962489, 
    -0.1441759, -0.1894231, -0.2065129, -0.2169459, -0.3770208, -0.5316597, 
    -0.4865261, -0.2724148, -0.2303737, -0.2227403, -0.1514349, -0.1026882, 
    -0.2479356, -0.3461289, -0.2281114, -0.1236029, -0.1148464, -0.05864522, 
    -0.03406841, -0.1209011, -0.2597194, -0.4701036, -0.6067734, -0.6750355, 
    -0.6699407, -0.5385606, -0.2573099, 0.02696681, 0.1615696, 0.2663548, 
    0.4063613, 0.7242005, 0.8928692, 0.8603008, 0.7660787, 0.7480605, 
    0.6729798, 0.522068, 0.336473, 0.2056785, 0.1342416, 0.02586031, 
    0.000436306, 0.0539031, 0.1661592, 0.3589654, 0.5143528, 0.5110812, 
    0.4840951, 0.4947567, 0.5094705, 0.4429173, 0.3050427, 0.1864071, 
    0.1225886, 0.09680772, 0.1146622, 0.08912492, -0.1283881, -0.2582382, 
    -0.3272974, -0.4295115, -0.4327996, -0.2401068, -0.04442012, 0.03155661, 
    0.1526339, 0.1742973, 0.1719537, 0.1821589, 0.1813123, 0.0737443, 
    0.04055691, 0.1985984, 0.223175, 0.3113251, 0.2902813, 0.3109999, 
    0.3337202, 0.348434, 0.3435035, 0.370863, 0.4078264, 0.4098606, 
    0.4352193, 0.4294734, 0.3355126, 0.3052552, 0.3478978, 0.209095,
  0.6234517, 0.5285463, 0.6384747, 0.5235658, 0.2969701, 0.2107396, 0.148109, 
    0.04607463, -0.006789923, 0.0022434, -0.1099473, -0.1550971, -0.01872027, 
    0.1025527, 0.05901426, -0.009508014, -0.08294547, -0.1798041, -0.3280299, 
    -0.3678737, -0.3045924, -0.2629584, -0.1868679, -0.1959825, -0.2830753, 
    -0.3367376, -0.3591337, -0.3479362, -0.2575061, -0.1782577, -0.03729129, 
    0.20755, 0.4987605, 0.5903946, 0.6638973, 0.7330053, 0.6623347, 
    0.5827451, 0.6845195, 0.9924293, 1.158266, 1.125616, 1.008168, 0.8525858, 
    0.6833639, 0.512465, 0.3336725, 0.179359, 0.1266251, 0.2080379, 
    0.4036922, 0.6257944, 0.7482553, 0.7257133, 0.689043, 0.7475395, 
    0.8310194, 0.7948866, 0.6609678, 0.5380344, 0.4775534, 0.3354139, 
    0.1106256, -0.1279812, -0.251744, -0.1750352, -0.04176641, 0.05613399, 
    0.1037416, 0.2333801, 0.3403618, 0.3006971, 0.2790664, 0.2877413, 
    0.3310846, 0.3395319, 0.2636528, 0.1776993, 0.1721163, 0.1430311, 
    0.03528452, 0.1184061, -0.01779175, 0.01850414, 0.05712605, 0.1828585, 
    0.2506967, 0.2553191, 0.3953581, 0.6000452, 0.7533498, 0.8811159, 
    0.94946, 0.9754376, 0.9965792, 0.876121,
  0.6042459, 0.555222, 0.3516095, 0.133754, 0.183217, 0.3617167, 0.3800924, 
    0.3063943, 0.431134, 0.6570125, 0.764711, 0.682403, 0.6238905, 0.549444, 
    0.3873998, 0.1619275, 0.05922604, 0.003724694, -0.03655863, -0.06736898, 
    -0.1205103, -0.1712102, -0.2123073, -0.23262, -0.2263536, -0.1612329, 
    -0.07418871, 0.03518629, 0.1021786, 0.1447239, 0.2622862, 0.5443661, 
    0.6993628, 0.5970674, 0.5703589, 0.6773736, 0.6737279, 0.6994275, 
    0.7601049, 0.9739883, 0.9646457, 0.62656, 0.3089817, 0.2544734, 
    0.2863255, 0.2593241, 0.2253561, 0.2042294, 0.2235003, 0.2866673, 
    0.4329567, 0.6018205, 0.6641412, 0.6639132, 0.6987276, 0.8337541, 
    0.924948, 0.8410776, 0.6526008, 0.4487278, 0.3136529, 0.1556289, 
    0.03038472, 0.02193761, 0.1396303, 0.2293437, 0.2870743, 0.3447733, 
    0.3933892, 0.4209771, 0.3969209, 0.3843397, 0.4965792, 0.658754, 
    0.7913716, 0.7082825, 0.5060039, 0.3306293, 0.209666, 0.1229796, 
    0.1112447, 0.07022905, 0.005304098, -0.1371932, -0.08463812, 0.1120744, 
    0.225421, 0.3023906, 0.4689918, 0.6358857, 0.7303677, 0.8630824, 
    0.9882784, 0.9458966, 0.7412248, 0.6047668,
  0.1454079, 0.1289041, -0.01242137, 0.05675173, 0.3035455, 0.67783, 
    0.7803853, 0.7342907, 0.7881806, 0.96126, 1.020489, 0.8743789, 0.6658662, 
    0.5584281, 0.4536754, 0.3977677, 0.3313614, 0.2161919, 0.1563449, 
    0.1724417, 0.2243464, 0.2472467, 0.2087541, 0.1475561, 0.09293365, 
    0.04700255, 0.06684303, 0.1017873, 0.1690727, 0.2929337, 0.4671855, 
    0.6161113, 0.5083308, 0.3555474, 0.352927, 0.5515273, 0.5658339, 
    0.3510227, 0.120196, -0.01219341, -0.1245632, -0.2376654, -0.2939479, 
    -0.2814479, -0.3534206, -0.4251328, -0.4191272, -0.2668645, -0.05705011, 
    0.1866348, 0.4283178, 0.609226, 0.7095841, 0.771921, 0.8057913, 0.852927, 
    0.8635389, 0.7601696, 0.5918756, 0.3914198, 0.2603652, 0.2462701, 
    0.3479466, 0.4121563, 0.3032038, 0.1916151, 0.1730441, 0.2626765, 
    0.3396944, 0.359942, 0.3408666, 0.4799126, 0.552146, 0.5614719, 
    0.4493468, 0.296824, 0.02198696, -0.1914897, -0.344696, -0.3374693, 
    -0.3405292, -0.2689474, -0.3600614, -0.5080916, -0.5592797, -0.5656934, 
    -0.503485, -0.3783221, -0.1620626, 0.03603268, 0.1332817, 0.21419, 
    0.2948868, 0.2566869, 0.1490047, 0.1251764,
  -0.3642441, -0.2316107, -0.1033554, 0.1359346, 0.3714001, 0.5796521, 
    0.5737926, 0.5565239, 0.5983859, 0.6646131, 0.674395, 0.5724421, 
    0.4212701, 0.2767714, 0.2207981, 0.2331353, 0.2579564, 0.3528292, 
    0.4141411, 0.4843233, 0.5086398, 0.477634, 0.4164035, 0.3730442, 
    0.3640924, 0.4031549, 0.3929009, 0.3883274, 0.4633601, 0.554327, 
    0.5807755, 0.5342422, 0.409714, 0.354001, 0.4312797, 0.5223932, 
    0.4348443, 0.1628392, -0.1449082, -0.2448759, -0.1712594, -0.06303978, 
    -0.03711203, -0.01562765, 0.01436913, 0.1050104, 0.2758924, 0.4376277, 
    0.5364721, 0.5986137, 0.66489, 0.7081517, 0.7340143, 0.7077774, 
    0.5629858, 0.4396133, 0.343145, 0.2255996, 0.1821914, 0.09750713, 
    0.1121067, 0.1702284, 0.2513485, 0.2056289, 0.04732788, -0.1046739, 
    -0.09103459, 0.1389296, 0.3763322, 0.3913711, 0.229099, -0.01956642, 
    -0.1678902, -0.3270044, -0.4692246, -0.5734401, -0.6072453, -0.5815781, 
    -0.5615748, -0.4834661, -0.3915227, -0.4130234, -0.5753608, -0.739049, 
    -0.6055854, -0.7723985, -0.8121771, -0.8248236, -0.8020045, -0.7864609, 
    -0.7994329, -0.7534696, -0.6159695, -0.4682971, -0.404967, -0.4046249,
  -0.2626328, -0.1665717, -0.02796495, 0.08582091, 0.1860976, 0.2849257, 
    0.3936172, 0.4745579, 0.578106, 0.6175104, 0.6035618, 0.5460422, 
    0.4344862, 0.3114231, 0.2592584, 0.2732558, 0.3460748, 0.4190729, 
    0.4964817, 0.5916477, 0.6176732, 0.5912245, 0.5479791, 0.5269179, 
    0.573565, 0.6684868, 0.6598606, 0.6283825, 0.6089492, 0.5676243, 
    0.5252905, 0.4761043, 0.420554, 0.3782688, 0.3561823, 0.3352838, 0.23211, 
    0.1310846, 0.05427796, 0.0978652, 0.142136, 0.1255182, 0.1241347, 
    0.2222305, 0.3822566, 0.6122695, 0.808168, 0.8919571, 0.9368302, 
    0.9703914, 0.900974, 0.7960261, 0.6805961, 0.5111952, 0.3388643, 
    0.2008436, 0.08391678, 0.04727918, 0.08141011, 0.1147109, 0.09065491, 
    0.02771546, 0.02034242, -0.02636983, -0.06704365, -0.05732686, 
    0.02752015, 0.1277155, 0.1585097, 0.004164159, -0.2242376, -0.3308131, 
    -0.2940944, -0.1650254, -0.1723334, -0.1719427, -0.1438015, -0.0631374, 
    -0.002541691, 0.01101625, -0.07918558, -0.1627632, -0.2776072, 
    -0.1980002, -0.2481954, -0.1483581, 0.0815568, -0.1099629, -0.2410996, 
    -0.4324901, -0.5700057, -0.6128285, -0.559394, -0.5018418, -0.4407253, 
    -0.3574408,
  -0.4869656, -0.4286485, -0.36011, -0.2415716, -0.06917582, 0.08696024, 
    0.2952448, 0.432761, 0.4244928, 0.3537084, 0.2592747, 0.1754043, 
    0.1093562, 0.1285293, 0.145554, 0.1937962, 0.2447566, 0.2942355, 
    0.3400689, 0.3577284, 0.3604954, 0.3571751, 0.3669407, 0.400095, 
    0.4751601, 0.6063775, 0.7031385, 0.7033339, 0.6512343, 0.6177382, 
    0.611716, 0.639483, 0.6758111, 0.6890272, 0.6086887, 0.6189101, 
    0.5692844, 0.4758762, 0.4361789, 0.3947564, 0.3664199, 0.3700331, 
    0.4253228, 0.5075006, 0.5718561, 0.5726537, 0.52197, 0.4114068, 
    0.3688776, 0.355222, 0.4040502, 0.4325819, 0.4161105, 0.4333472, 
    0.4047329, 0.3526013, 0.3206354, 0.3732558, 0.348614, 0.4758438, 
    0.4173963, 0.3429825, 0.18753, 0.07149816, 0.006654263, 0.0004042387, 
    0.01978901, -0.04347594, -0.1995795, -0.3502468, -0.4077012, -0.2457709, 
    -0.04108337, -0.0192572, 0.031638, -0.1148789, -0.140058, -0.1945827, 
    -0.1686062, -0.2414902, -0.1547227, -0.06211185, -0.08507681, 
    -0.06014204, -0.07954311, -0.02658176, -0.06872022, -0.1318712, 
    -0.07482362, 0.0114556, -0.02778566, -0.08387315, -0.1720406, -0.2868842, 
    -0.4095567, -0.4981471,
  -0.1139838, -0.22331, -0.2480822, -0.2082382, -0.138284, -0.06098902, 
    -0.03170842, -0.06640893, -0.1353217, -0.211819, -0.2319199, -0.2050157, 
    -0.1479193, -0.06426039, 0.0009739399, 0.03124735, 0.1072402, 0.1453099, 
    0.1978652, 0.2042617, 0.189776, 0.205401, 0.2851862, 0.3811009, 
    0.5095514, 0.6666966, 0.8017714, 0.855401, 0.8630182, 0.7964328, 0.75947, 
    0.7491509, 0.7195611, 0.7085748, 0.7024063, 0.7845678, 0.7898899, 
    0.7880833, 0.7241673, 0.7226211, 0.6385879, 0.6587865, 0.6177058, 
    0.6142552, 0.5667292, 0.4221491, 0.2334284, 0.07055408, -0.1487004, 
    -0.3975124, -0.5901397, -0.5958358, -0.5270207, -0.4159856, -0.3096867, 
    -0.2346547, -0.2630887, -0.3723824, -0.4660347, -0.4992378, -0.5203316, 
    -0.6009468, -0.568704, -0.356562, -0.3139511, -0.2893907, -0.287405, 
    -0.3058295, -0.2858262, -0.2883164, -0.1856797, -0.08968364, -0.04435486, 
    0.03363994, -0.003697276, -0.05866151, -0.06465107, -0.1976263, 
    -0.08250594, 0.04796267, 0.1435523, -0.01315308, -0.0411489, -0.1154976, 
    -0.1655462, -0.280504, -0.5101753, -0.5465035, -0.3893907, -0.2156601, 
    0.1112603, 0.1206517, 0.2150038, 0.1958957, 0.1303035, 0.02000058,
  0.07000077, 0.08450222, 0.0946424, 0.1379204, 0.1976047, 0.2456353, 
    0.2429334, 0.2309219, 0.2048478, 0.1484511, 0.1040012, 0.03700906, 
    0.02232808, -0.03690046, -0.04847276, -0.06806898, -0.02417254, 
    -0.01606709, -0.02684183, 0.006458938, 0.1341119, 0.2377578, 0.3738418, 
    0.5229141, 0.6769342, 0.8278131, 0.8703099, 0.9260228, 0.9089817, 
    0.8208308, 0.7613255, 0.5263808, 0.4744114, 0.5000951, 0.4805638, 
    0.4763807, 0.5131484, 0.4998347, 0.477862, 0.4875951, 0.4700332, 
    0.451625, 0.420261, 0.3952284, 0.3207005, 0.2291151, 0.1051568, 
    -0.006773472, -0.1098497, -0.1882349, -0.2305202, -0.2131373, -0.1872586, 
    -0.1505234, -0.157343, -0.1952988, -0.2708033, -0.3709826, -0.4320664, 
    -0.4914252, -0.5834336, -0.621487, -0.6624864, -0.6337267, -0.6496121, 
    -0.5824734, -0.5412461, -0.4813828, -0.4024278, -0.302558, -0.2076361, 
    -0.1228379, -0.1017116, -0.09769143, -0.1729844, -0.318655, -0.4915233, 
    -0.5072453, -0.1631699, -0.1532898, -0.2326679, -0.1982768, -0.09787059, 
    -0.01554632, -0.008335948, -0.1118517, -0.2144225, -0.205308, -0.1557477, 
    -0.1268737, -0.05436492, 0.04586339, -0.001500033, -0.08750254, 
    -0.05695254, 0.04340553,
  0.02473694, 0.02148163, 0.07815492, 0.132875, 0.2977186, 0.2723932, 
    0.224802, 0.09078503, 0.04828838, -0.007750034, -0.1241563, -0.2071478, 
    -0.2442897, -0.249433, -0.2893255, -0.3095241, -0.3595242, -0.2635444, 
    -0.229267, -0.1619167, -0.1351264, -0.1412461, -0.03852808, 0.05046934, 
    0.09425193, 0.2347142, 0.2313938, 0.2034641, 0.200453, 0.1838841, 
    0.1385065, 0.1074192, 0.1006321, 0.09592831, 0.08204484, 0.05626363, 
    0.03668356, 0.01879615, 0.01030004, -0.01190042, -0.03952086, 
    -0.08065033, -0.114, -0.1565131, -0.1854357, -0.228144, -0.2696642, 
    -0.3199246, -0.3684597, -0.4055203, -0.4360378, -0.4448432, -0.4456082, 
    -0.4446805, -0.4606798, -0.4633165, -0.475019, -0.482278, -0.4916368, 
    -0.49914, -0.4933946, -0.4769232, -0.4621446, -0.4593451, -0.4660508, 
    -0.4631537, -0.4480821, -0.4361355, -0.4192735, -0.3888535, -0.3459011, 
    -0.3190131, -0.3148952, -0.194241, -0.1787787, -0.1989124, -0.2166535, 
    -0.2309598, -0.2452173, -0.2254908, -0.1699734, -0.1023138, -0.02513278, 
    0.02856159, 0.03456783, -0.0001974106, -0.06268096, -0.1023946, 
    -0.127655, -0.1019235, -0.09455025, -0.07155204, 0.008688748, 
    -0.02964131, -0.004820347, -0.01539981,
  0.06295311, 0.133233, 0.1812637, 0.2090306, 0.2105931, 0.1836237, 
    0.1665175, 0.1390761, 0.1100071, 0.07003317, 0.01625712, -0.02667907, 
    -0.0729844, -0.1072617, -0.1434271, -0.1556179, -0.1631212, -0.1788601, 
    -0.1938177, -0.2077011, -0.2262722, -0.24053, -0.2809923, -0.3190294, 
    -0.3701036, -0.3950873, -0.4331407, -0.4867865, -0.5395046, -0.5961616, 
    -0.6406114, -0.7107612, -0.753437, -0.7783067, -0.7989285, -0.8063992, 
    -0.8202664, -0.8302924, -0.834101, -0.8394558, -0.8481635, -0.8583848, 
    -0.8612983, -0.8612494, -0.8534858, -0.8375841, -0.8117702, -0.7875026, 
    -0.7560247, -0.722545, -0.6869493, -0.6565619, -0.6313992, -0.6000352, 
    -0.5704779, -0.5430528, -0.5162136, -0.480097, -0.4567084, -0.4273952, 
    -0.3839707, -0.3472357, -0.316653, -0.2940456, -0.2652533, -0.2401231, 
    -0.209931, -0.1827989, -0.1544134, -0.1363145, -0.1229681, -0.1204942, 
    -0.1178738, -0.1337104, -0.1854031, -0.2153998, -0.2489609, -0.2998236, 
    -0.3004421, -0.3049668, -0.32025, -0.2837591, -0.2916692, -0.3094264, 
    -0.2950383, -0.2706243, -0.2533066, -0.3117539, -0.3274928, -0.3863634, 
    -0.3914089, -0.3817246, -0.3174994, -0.2177598, -0.1145371, -0.01443949,
  0.2740208, 0.3111465, 0.3539362, 0.3871393, 0.4090143, 0.4237929, 
    0.4307916, 0.431459, 0.423793, 0.4071588, 0.3795384, 0.3450332, 
    0.3012181, 0.2607721, 0.2167291, 0.1589166, 0.09408917, 0.0285618, 
    -0.0447129, -0.1196478, -0.1954128, -0.2683621, -0.3408066, -0.4045436, 
    -0.4668483, -0.5191271, -0.5698432, -0.6238634, -0.6681993, -0.7121934, 
    -0.7555203, -0.7947781, -0.8341661, -0.864586, -0.8822944, -0.8944362, 
    -0.9017931, -0.9018092, -0.8973984, -0.8966823, -0.8874213, -0.8768907, 
    -0.8632188, -0.8468125, -0.823489, -0.8039415, -0.7809923, -0.7523139, 
    -0.7254584, -0.6943223, -0.6586289, -0.6152859, -0.5738633, -0.5361354, 
    -0.5028184, -0.4579291, -0.4145371, -0.3764837, -0.3330267, -0.2951687, 
    -0.2627142, -0.2315944, -0.1959825, -0.1691433, -0.1428574, -0.1121771, 
    -0.08561461, -0.06479756, -0.04178324, -0.02348897, -0.01097269, 
    -0.009019554, -0.002525419, -0.0007350594, -0.01020771, -0.02228455, 
    -0.04440369, -0.05864521, -0.07921813, -0.1006862, -0.1161973, 
    -0.1248562, -0.1351426, -0.1408067, -0.1465033, -0.1481634, -0.1281602, 
    -0.1064805, -0.07733011, -0.0396348, -0.004804071, 0.0224583, 0.05859112, 
    0.1162246, 0.1750625, 0.2259576,
  -0.1340685, -0.1530304, -0.1718779, -0.1904655, -0.2088733, -0.2270047, 
    -0.2449897, -0.2620633, -0.2777371, -0.2915066, -0.302168, -0.3108265, 
    -0.3160841, -0.3182647, -0.3180046, -0.3159864, -0.3124382, -0.3083532, 
    -0.3022981, -0.2967958, -0.2901392, -0.2827339, -0.2739444, -0.2616067, 
    -0.2460961, -0.2251487, -0.1980977, -0.1654482, -0.1281929, -0.08672142, 
    -0.04269457, 0.002682686, 0.0484674, 0.09416986, 0.1383431, 0.1806774, 
    0.2206838, 0.2574999, 0.2907687, 0.3209771, 0.3473768, 0.3702772, 
    0.3899549, 0.4065561, 0.4200001, 0.4311495, 0.4421515, 0.4422655, 
    0.4448535, 0.4478326, 0.4488583, 0.4499335, 0.4592428, 0.5016913, 
    0.5082994, 0.5105453, 0.4963365, 0.477212, 0.5302391, 0.4750471, 
    0.4633613, 0.4923, 0.4475408, 0.4423652, 0.4367008, 0.4340806, 0.4302068, 
    0.4379215, 0.439239, 0.4221983, 0.4149227, 0.4068499, 0.4023738, 
    0.3781867, 0.3299942, 0.3422022, 0.2932754, 0.3063622, 0.3026514, 
    0.2785306, 0.2526031, 0.226903, 0.2004051, 0.1727524, 0.1433091, 
    0.1164212, 0.09073734, 0.0651679, 0.0394516, 0.01412582, -0.009603977, 
    -0.03213072, -0.05437994, -0.07570219, -0.09525013, -0.1149285,
  0.09163141, 0.07556689, 0.05557992, 0.03326546, 0.007858545, -0.01813427, 
    -0.04101843, -0.05761993, -0.06675082, -0.07041287, -0.07148713, 
    -0.07420522, -0.08312452, -0.09876579, -0.1177437, -0.1388048, 
    -0.1600783, -0.1793488, -0.1952342, -0.2066603, -0.2182159, -0.2301626, 
    -0.2427442, -0.2579625, -0.2789912, -0.3021836, -0.3274927, -0.3490734, 
    -0.3601742, -0.3578305, -0.3413262, -0.3111343, -0.2692399, -0.2172542, 
    -0.1575212, -0.09433746, -0.03081226, 0.02983189, 0.0831027, 0.1252244, 
    0.1618131, 0.1688124, 0.1623833, 0.1346653, 0.1150686, 0.07900071, 
    0.06674504, 0.06334305, 0.0421679, 0.02336955, -0.01325202, 0.0008273125, 
    0.009990215, -0.0059762, 0.003284693, -0.01521969, -0.009506702, 
    -0.003793716, 0.01401234, 0.02822113, 0.04739428, 0.07420063, 0.1026993, 
    0.1325977, 0.1647751, 0.1999807, 0.2332977, 0.2456515, 0.2648898, 
    0.2762017, 0.3154432, 0.3282525, 0.3203749, 0.3634087, 0.3022597, 
    0.3307101, 0.326869, 0.3352836, 0.3356254, 0.2614878, 0.3366182, 
    0.3625295, 0.3605111, 0.364336, 0.4388478, 0.4423151, 0.3997369, 
    0.3673153, 0.3274717, 0.2829237, 0.2396286, 0.198369, 0.1637342, 
    0.1379037, 0.1161913, 0.1022921,
  -0.06816721, -0.09207633, -0.1016141, -0.112812, -0.1253283, -0.1329292, 
    -0.131741, -0.1179227, -0.09149039, -0.05469026, -0.01898064, 
    -0.001858234, -0.006269217, -0.0334667, -0.08917952, -0.1645706, 
    -0.2472851, -0.3272977, -0.395885, -0.4398141, -0.4502149, -0.4193883, 
    -0.3464057, -0.260338, -0.2057319, -0.1988797, -0.2385125, -0.3086457, 
    -0.3863313, -0.4629264, -0.5272, -0.5767937, -0.5991726, -0.5846205, 
    -0.5358415, -0.4594584, -0.3655615, -0.266408, -0.1634293, -0.06235504, 
    0.0325346, 0.1482244, 0.179359, 0.1919887, 0.1218234, 0.09190804, 
    0.03684616, -0.01356071, -0.07168245, -0.1337756, -0.1883003, -0.224368, 
    -0.2323595, -0.2224799, -0.2092963, -0.1882842, -0.1695992, -0.1667184, 
    -0.1563178, -0.1265979, -0.08401966, -0.03927708, 0.001315355, 
    0.03798544, 0.07880586, 0.1192518, 0.1514946, 0.18377, 0.2271132, 
    0.2810519, 0.3359346, 0.3616346, 0.3503554, 0.354701, 0.3554823, 
    0.3634901, 0.358119, 0.44391, 0.4870903, 0.5425916, 0.5968069, 0.636927, 
    0.6302704, 0.5905567, 0.6542773, 0.684258, 0.6466606, 0.5841441, 
    0.506361, 0.4605277, 0.3182755, 0.2163224, 0.1199348, 0.03339505, 
    -0.01369119, -0.04715502,
  -0.4772162, -0.445771, -0.4010932, -0.3438349, -0.3071485, -0.2998402, 
    -0.3198762, -0.3481638, -0.3621775, -0.3461131, -0.2912468, -0.2207873, 
    -0.1523954, -0.0931831, -0.0550646, -0.06373973, -0.1446806, -0.2722203, 
    -0.3979039, -0.4808936, -0.5112648, -0.5031595, -0.4905295, -0.4604204, 
    -0.378795, -0.2714383, -0.2249539, -0.2318876, -0.2777209, -0.3469754, 
    -0.424075, -0.4931669, -0.554202, -0.6263051, -0.7013539, -0.7801623, 
    -0.8462107, -0.870151, -0.8516779, -0.8007832, -0.6985698, -0.5335464, 
    -0.3181653, -0.0695653, 0.08256507, 0.1026011, -0.1241894, -0.1147816, 
    -0.2076362, -0.2939969, -0.3480497, -0.3889676, -0.4183621, -0.4300483, 
    -0.4362983, -0.4711618, -0.6009145, -0.5371288, -0.5973012, -0.5792515, 
    -0.4990432, -0.4749377, -0.4192574, -0.3572297, -0.3353221, -0.2840846, 
    -0.2072453, -0.1232128, -0.02387953, 0.0518527, 0.1116827, 0.1783657, 
    0.244626, 0.3187957, 0.3741343, 0.4609505, 0.5057096, 0.47988, 0.4461073, 
    0.6241997, 0.6480767, 0.7148247, 0.7736951, 0.824867, 0.8485647, 
    0.8530407, 0.8230762, 0.7586395, 0.7593071, 0.677552, 0.4547329, 
    0.2270479, 0.08596802, -0.1673841, -0.370347, -0.4687195,
  -0.1379571, -0.1502619, -0.1212907, -0.04956198, -0.02575016, 0.03917503, 
    0.05344915, 0.02949047, -0.1411638, -0.08634567, -0.07472467, 
    -0.005372524, 0.06980658, 0.1016912, 0.1225228, 0.2176405, 0.2674615, 
    0.2424614, 0.2048801, 0.123955, -0.03900003, -0.01455212, 0.01865101, 
    -0.0221529, -0.1034679, -0.1439471, -0.1295595, -0.1186061, -0.130846, 
    -0.1809924, -0.2444208, -0.2754266, -0.2923539, -0.3003285, -0.3266309, 
    -0.3952668, -0.5064321, -0.636754, -0.7553902, -0.8319526, -0.8024768, 
    -0.6840525, -0.468981, -0.2196484, -0.009248137, 0.1101209, 0.009730101, 
    0.01298559, -0.03039008, -0.05799431, -0.06992459, -0.06618112, 
    -0.005308747, 0.03175181, -0.01136339, -0.09518507, -0.2715522, 
    -0.4985705, -0.6904812, -0.82012, -0.8538441, -0.8059272, -0.7100776, 
    -0.5834501, -0.495885, -0.4122097, -0.335322, -0.2872914, -0.2549187, 
    -0.19333, -0.2516961, -0.2114123, -0.1705269, -0.1060252, -0.06212878, 
    0.06173193, 0.15877, 0.2119927, 0.1708468, 0.2589653, 0.2794406, 
    0.3440239, 0.3900038, 0.4391574, 0.4768853, 0.5276177, 0.5956841, 
    0.6780568, 0.7438446, 0.7994599, 0.8567512, 0.7756476, 0.6137505, 
    0.4317036, 0.1865058, -0.08787584,
  0.3531218, 0.3651824, 0.1122689, 0.1479459, 0.1324999, 0.1274219, 
    0.07628298, 0.01853538, 0.04443073, 0.03186536, 0.0003547668, 
    -0.005455256, 0.05354691, 0.1030583, 0.05986118, 0.05144525, 0.1388314, 
    0.1494273, 0.1752411, 0.2235972, 0.04667664, 0.02698278, 0.05121899, 
    0.09998226, 0.05354691, 0.02092934, -0.009197235, -0.05273581, 
    -0.1306167, -0.2420588, -0.3542166, -0.4302421, -0.4333186, -0.3300467, 
    -0.203403, -0.1310568, -0.1332059, -0.198554, -0.2601104, -0.3420599, 
    -0.3761582, -0.3458042, -0.2609894, -0.174401, -0.03760064, 0.009648979, 
    0.04135466, 0.0744113, 0.1175103, 0.1650527, 0.2093723, 0.2707328, 
    0.3454888, 0.4238254, 0.4927543, 0.5426401, 0.5247529, 0.4068164, 
    0.2137338, 0.01374984, -0.1519235, -0.2747099, -0.3191762, -0.3118194, 
    -0.2743685, -0.2389842, -0.2107451, -0.1752961, -0.114212, -0.08979797, 
    -0.06772768, -0.03441036, -0.03152955, -0.02277291, 0.02270234, 
    0.04941142, 0.1187798, 0.1685845, 0.1859673, 0.1932427, 0.159372, 
    0.1611624, 0.1629367, 0.1624322, 0.1368788, 0.1220024, 0.1402316, 
    0.1581516, 0.2454888, 0.356703, 0.4641085, 0.5845187, 0.6476369, 
    0.6155405, 0.5533659, 0.4574833,
  0.7650852, 0.7475395, 0.7121066, 0.6310193, 0.5861138, 0.5740532, 
    0.6092257, 0.6264946, 0.6071424, 0.5762179, 0.5978651, 0.674395, 
    0.7554494, 0.7601043, 0.7008108, 0.6915985, 0.6986461, 0.6767873, 
    0.676462, 0.6985487, 0.6838676, 0.6402968, 0.5704559, 0.4499644, 
    0.4038055, 0.3314745, 0.2595344, 0.2250134, 0.2158823, 0.1707325, 
    0.1627898, 0.1639452, 0.1502247, -0.001516342, 0.074965, 0.1834929, 
    0.2509894, 0.3540332, 0.435137, 0.5326467, 0.5888314, 0.5857391, 
    0.5627081, 0.5418589, 0.5418429, 0.5395317, 0.5561496, 0.5003878, 
    0.4849416, 0.4914681, 0.5619925, 0.6332164, 0.6707971, 0.7805953, 
    0.8577113, 0.9723923, 1.092998, 1.162383, 1.142933, 1.006296, 0.8163869, 
    0.6285121, 0.4909956, 0.3848598, 0.3179653, 0.2788212, 0.2740035, 
    0.2974577, 0.3530564, 0.4715621, 0.486536, 0.4856737, 0.4401169, 
    0.4698858, 0.4191046, 0.3717086, 0.321367, 0.2591436, 0.1947067, 
    0.2750614, 0.3256638, 0.3722785, 0.4219203, 0.457516, 0.4580042, 
    0.4195766, 0.3647914, 0.3654749, 0.3942516, 0.4370738, 0.4974087, 
    0.5501108, 0.5823212, 0.6421194, 0.7064751, 0.7530571,
  0.9117482, 0.9551563, 0.9309373, 0.9093552, 0.9138479, 0.9588349, 
    0.9564424, 0.9297986, 0.883786, 0.8535452, 0.8950815, 1.020683, 1.188799, 
    1.324314, 1.468926, 1.478513, 1.489759, 1.496107, 1.521465, 1.571774, 
    1.583411, 1.539173, 1.46572, 1.437025, 1.462253, 1.495619, 1.504017, 
    1.503334, 1.498923, 1.509828, 1.574769, 1.688473, 1.945489, 2.088734, 
    2.261146, 1.920408, 1.536911, 1.474509, 1.353903, 1.355303, 1.506605, 
    1.731702, 1.959648, 2.243779, 2.303041, 2.297442, 2.275599, 2.10698, 
    1.766143, 1.509063, 1.385496, 1.327, 1.355613, 1.240932, 1.154506, 
    1.261912, 1.373419, 1.520994, 1.518243, 1.559454, 1.644871, 1.639369, 
    1.737432, 1.808738, 1.700047, 1.543617, 1.45672, 1.397605, 1.391388, 
    1.316746, 1.235073, 1.096043, 1.02547, 0.9789367, 1.097931, 1.23434, 
    1.468406, 1.602098, 1.793992, 1.819497, 1.797524, 1.721026, 1.488133, 
    1.156068, 0.9986627, 0.8925917, 0.7551727, 0.6086397, 0.5121067, 
    0.5431776, 0.6003878, 0.6259737, 0.6188774, 0.6369917, 0.7003057, 
    0.8169072,
  0.9749651, 1.089402, 1.190916, 1.300388, 1.463621, 1.525925, 1.49894, 
    1.634683, 1.750893, 1.949364, 1.985659, 2.184292, 2.427261, 2.527195, 
    2.925096, 3.147931, 3.220815, 3.321157, 3.405158, 3.52573, 3.26808, 
    2.911554, 2.621612, 2.504034, 2.309779, 2.181557, 2.07018, 2.025779, 
    2.242722, 2.356199, 2.340688, 2.354962, 2.34129, 2.363833, 2.297394, 
    2.188848, 2.094611, 2.004262, 1.895213, 1.838637, 1.937954, 2.215868, 
    2.558722, 2.833819, 2.97993, 3.022622, 2.986163, 2.914971, 2.852976, 
    2.818276, 2.825063, 2.821661, 2.767934, 2.680288, 2.578839, 2.50646, 
    2.430825, 2.377098, 2.379848, 2.383901, 2.290542, 2.129377, 1.995034, 
    1.978139, 1.933136, 1.76175, 1.509666, 1.331362, 1.26743, 1.251952, 
    1.250747, 1.232827, 1.140038, 1.051431, 1.090949, 1.277147, 1.479929, 
    1.518814, 1.412677, 1.322736, 1.362807, 1.424266, 1.36048, 1.333576, 
    1.470962, 1.807827, 1.90672, 1.570799, 1.037286, 0.8115864, 0.8159161, 
    0.7188778, 0.5790181, 0.5282044, 0.5908833, 0.7580872,
  1.937743, 1.864468, 1.986343, 2.080776, 1.997053, 2.002847, 2.028204, 
    1.90615, 1.87171, 1.787611, 1.613669, 1.494806, 1.48102, 1.587383, 
    1.7645, 1.861147, 1.927847, 1.998404, 2.076869, 2.15047, 2.376072, 
    2.556297, 2.586522, 2.559113, 2.469578, 2.184341, 2.091974, 2.072247, 
    2.081525, 2.077928, 1.984666, 1.811391, 1.63867, 1.563996, 1.582843, 
    1.683657, 1.915476, 2.17534, 2.309975, 2.314483, 2.294937, 2.275518, 
    2.252146, 2.307159, 2.502618, 2.680873, 2.743797, 2.798143, 2.920197, 
    3.145538, 3.366014, 3.452878, 3.320278, 3.074558, 2.896401, 2.81769, 
    2.671695, 2.420848, 2.181281, 2.048094, 1.951479, 1.774201, 1.648046, 
    1.664061, 1.713914, 1.698273, 1.642154, 1.528059, 1.336066, 1.169595, 
    1.110155, 1.090005, 1.069155, 1.05353, 1.080191, 1.095539, 1.095978, 
    1.165119, 1.108771, 0.9214177, 0.9902482, 1.110936, 1.207274, 1.18478, 
    1.123143, 1.184438, 1.397036, 1.58395, 1.80576, 1.687303, 1.744579, 
    1.922004, 1.963264, 1.905614, 1.87093, 1.812499,
  1.207924, 1.249396, 1.275437, 1.270148, 1.291144, 1.345392, 1.424688, 
    1.446385, 1.396564, 1.324429, 1.261049, 1.207614, 1.132549, 1.091127, 
    1.101234, 1.110739, 1.135104, 1.22957, 1.313571, 1.290801, 1.22573, 
    1.16813, 1.118959, 1.146222, 1.278155, 1.465247, 1.618877, 1.626512, 
    1.521352, 1.415507, 1.333477, 1.235202, 1.168682, 1.21126, 1.297638, 
    1.317331, 1.313896, 1.342217, 1.358429, 1.423582, 1.611993, 1.746808, 
    1.688946, 1.658949, 1.825454, 2.02114, 2.136164, 2.202831, 2.266438, 
    2.382437, 2.487466, 2.555907, 2.523028, 2.386294, 2.249363, 2.170376, 
    2.080125, 1.95869, 1.855516, 1.796906, 1.714972, 1.579767, 1.431314, 
    1.319237, 1.221239, 1.170002, 1.112254, 0.9855294, 0.8302879, 0.8369775, 
    0.9302554, 0.9475412, 0.8667464, 0.7818666, 0.7201481, 0.6037908, 
    0.4857078, 0.6207829, 0.7733383, 0.8828921, 0.8599596, 0.9281564, 
    1.085546, 1.201756, 1.216665, 1.210821, 1.23587, 1.299055, 1.350145, 
    1.382209, 1.376333, 1.322117, 1.278107, 1.267202, 1.240005, 1.193357,
  1.087678, 1.028204, 0.9607077, 0.8940086, 0.8718729, 0.898386, 0.8881006, 
    0.7554502, 0.5880184, 0.5288715, 0.5472803, 0.5144835, 0.4680967, 
    0.4441385, 0.4582491, 0.4721823, 0.4871063, 0.5834608, 0.679018, 0.73172, 
    0.8718729, 0.9452295, 0.8605289, 0.8064756, 0.8273582, 0.8239069, 
    0.8256655, 0.8546038, 0.9223108, 0.9525194, 0.8799295, 0.764451, 
    0.6766415, 0.6270647, 0.614419, 0.5878229, 0.5322399, 0.5251446, 
    0.5467091, 0.5231581, 0.6030579, 0.7237287, 0.7357564, 0.685008, 
    0.7252913, 0.7669415, 0.7359357, 0.7097478, 0.7655749, 0.9516587, 
    1.147199, 1.237742, 1.203807, 1.093228, 1.04269, 1.026415, 1.034943, 
    1.12311, 1.260122, 1.31092, 1.262108, 1.131151, 0.9960923, 0.8415022, 
    0.682209, 0.5860987, 0.5525699, 0.5000472, 0.4429507, 0.3921857, 
    0.4037747, 0.4383287, 0.3727202, 0.2543602, 0.2206693, 0.1605291, 
    0.01461267, -0.03221178, -0.05817223, -0.05665874, 0.1152816, 0.473176, 
    0.7857246, 0.9306788, 0.9722152, 1.007095, 1.085741, 1.129572, 1.108055, 
    1.154149, 1.252521, 1.301056, 1.280532, 1.220359, 1.160333, 1.126219,
  0.6687489, 0.614614, 0.5550766, 0.4786935, 0.401659, 0.3415675, 0.2971501, 
    0.1338363, -0.09274244, -0.1502132, -0.09311676, -0.02339029, 0.04449701, 
    0.1068182, 0.1770821, 0.228888, 0.2206697, 0.2815895, 0.3688622, 
    0.4233055, 0.6057434, 0.7328749, 0.6841936, 0.6646957, 0.6596498, 
    0.6437969, 0.5754375, 0.4195452, 0.2885227, 0.1762018, 0.03228951, 
    -0.03755093, -0.05639839, -0.1676302, -0.2320166, -0.1570997, -0.2332048, 
    -0.4226589, -0.4370298, -0.3967953, -0.3859882, -0.3370132, -0.2943048, 
    -0.2575049, -0.2068539, -0.1752291, -0.1315932, -0.259881, -0.3623061, 
    -0.3004575, -0.05883932, 0.05372572, -0.0561862, -0.2327981, -0.1931658, 
    0.07561684, 0.2765613, 0.3739734, 0.4650865, 0.5810046, 0.663898, 
    0.6458311, 0.5870748, 0.523273, 0.4229317, 0.3058414, 0.197557, 
    0.09168148, -0.04952955, -0.2844253, -0.4589696, -0.4106464, -0.3697772, 
    -0.4993181, -0.6386085, -0.670135, -0.6045918, -0.6466336, -0.7481952, 
    -0.7705588, -0.5382504, -0.1955581, 0.06453276, 0.2742496, 0.42202, 
    0.4288073, 0.4361315, 0.5145655, 0.607502, 0.7039862, 0.7993307, 
    0.8689928, 0.8510399, 0.7095361, 0.5914369, 0.6297674,
  0.2042956, 0.1360664, 0.05024242, -0.03439283, -0.06725407, -0.1579766, 
    -0.2281761, -0.1981959, -0.3115914, -0.4050157, -0.3357618, -0.2946968, 
    -0.277297, -0.2496109, -0.1807308, -0.09814596, -0.1766129, -0.2290869, 
    -0.1604505, -0.1519871, -0.09482574, -0.05957222, -0.086689, -0.06036949, 
    -0.03621674, 0.07338619, 0.1063299, -0.04077435, -0.1270704, -0.2292519, 
    -0.4206562, -0.6610694, -0.834393, -0.9260592, -1.017173, -0.9315605, 
    -0.8779964, -0.9690285, -0.9471374, -0.9279156, -0.9431987, -0.8392758, 
    -0.8109388, -0.8380389, -0.8934259, -1.016685, -1.04839, -1.037112, 
    -1.242906, -1.348374, -1.235647, -1.161721, -1.19079, -1.211363, 
    -1.137275, -0.9126329, -0.6776066, -0.4521508, -0.2682972, -0.07480717, 
    0.1088843, 0.1177382, 0.03572321, -0.05343676, -0.1833687, -0.2200871, 
    -0.2546248, -0.4109554, -0.5704284, -0.7366228, -0.8503113, -0.9995461, 
    -1.134507, -1.163853, -1.291278, -1.314439, -1.030667, -0.9659696, 
    -1.110061, -1.009492, -0.8241892, -0.8260124, -0.8145375, -0.8060086, 
    -0.6296418, -0.3276236, -0.1562207, 0.01098299, 0.1568003, 0.1974754, 
    0.2320461, 0.3144679, 0.3686504, 0.3062158, 0.2370753, 0.2281075,
  -0.5035996, -0.5465527, -0.5015333, -0.5151072, -0.4850457, -0.556383, 
    -0.6851428, -0.5534533, -0.5336291, -0.7437368, -0.8439647, -0.8954784, 
    -0.9946643, -1.025898, -1.066133, -1.056107, -1.128713, -1.256284, 
    -1.280373, -1.40311, -1.454087, -1.363478, -1.257, -1.109002, -1.05062, 
    -0.923439, -0.8601089, -0.8343439, -0.746079, -0.9529638, -1.165855, 
    -1.3001, -1.409573, -1.158759, -1.091311, -1.147366, -1.000149, 
    -0.771227, -0.6113474, -0.720185, -0.7078643, -0.5833361, -0.8757358, 
    -1.275915, -1.58109, -1.818314, -2.038609, -2.183173, -2.291555, 
    -2.380569, -2.203714, -2.041556, -1.958792, -1.772415, -1.618232, 
    -1.471032, -1.335045, -1.143347, -0.8881705, -0.7224805, -0.5781446, 
    -0.4922721, -0.4169142, -0.3885779, -0.5588737, -0.6714387, -0.7118196, 
    -0.7481153, -0.7463086, -0.8970411, -1.054691, -1.259313, -1.407522, 
    -1.308402, -1.284801, -1.089115, -0.5449409, -0.4131376, -0.926191, 
    -0.8713244, -0.7014188, -0.9230496, -1.026158, -1.253746, -1.218769, 
    -0.7386746, -0.4709012, -0.3459991, -0.245723, -0.2224157, -0.09414363, 
    0.04268885, 0.04783249, -0.05128765, -0.2245789, -0.3812366,
  -0.8268099, -0.9293323, -0.8185412, -0.715172, -0.5214871, -0.2416206, 
    -0.2637235, -0.3792671, -0.4600939, -0.8461291, -1.275833, -1.44582, 
    -1.614521, -1.486201, -1.463805, -1.566718, -1.547806, -1.742988, 
    -1.8668, -1.974775, -2.080309, -2.028828, -1.991344, -1.872268, 
    -1.820364, -1.629674, -1.406123, -1.276142, -1.132995, -1.191409, 
    -0.8952342, -0.6822293, -0.872187, -0.6273465, -0.4690295, -0.4381375, 
    -0.3789741, -0.4036161, -0.4923693, -0.7099637, -0.6094592, -0.5966174, 
    -1.08083, -1.446699, -1.779853, -2.069778, -2.407197, -2.755618, 
    -2.873717, -2.942695, -2.739244, -2.357816, -2.097138, -1.83153, 
    -1.587747, -1.374824, -1.304186, -1.349987, -1.286787, -1.295397, 
    -1.246585, -1.111803, -0.9557647, -0.7550161, -0.7227895, -0.6881378, 
    -0.7254425, -0.8461619, -0.8537954, -0.9620634, -0.9808297, -0.9561714, 
    -1.054641, -1.078258, -1.0522, -0.7912951, -0.2695991, -0.04373682, 
    -0.5577339, -0.5785999, -0.3497587, -0.5613308, -0.7165394, -0.8633331, 
    -1.03275, -0.8305203, -0.6834337, -0.5528836, -0.3830268, -0.4348499, 
    -0.5383493, -0.5692087, -0.613919, -0.6805696, -0.7857291, -0.7914745,
  -0.8085804, -0.8133982, -0.7051957, -0.6115913, -0.3754591, 0.104994, 
    0.1585747, -0.2145535, -0.286754, -0.4323928, -0.8597202, -1.078714, 
    -1.573977, -1.583759, -1.14976, -1.271878, -1.288741, -1.429642, 
    -1.485143, -1.504251, -1.653747, -1.691019, -1.698815, -1.609654, 
    -1.643818, -1.564, -1.391393, -1.275345, -1.049043, -0.8203644, 
    -0.2933295, -0.1384305, -0.48096, -0.4160513, -0.3876492, -0.3415716, 
    -0.2744981, -0.3665066, -0.5269071, -0.8446479, -0.8305368, -1.020934, 
    -1.482099, -1.506025, -1.647252, -1.933987, -2.18983, -2.530846, 
    -2.560192, -2.344615, -2.054837, -1.744225, -1.539098, -1.32375, 
    -1.08319, -0.9725451, -1.058792, -1.296861, -1.386005, -1.348245, 
    -1.2536, -1.055504, -0.8435738, -0.6929064, -0.7723985, -0.7519071, 
    -0.5955268, -0.6388866, -0.6576198, -0.6619657, -0.677119, -0.7681834, 
    -0.8363475, -0.7761425, -0.5535674, -0.2559272, -0.1830595, 0.2092582, 
    -0.0730496, -0.3070505, -0.02192658, -0.02290344, -0.3100617, -0.2885444, 
    -0.7391474, -0.9425654, -0.7216989, -0.5247263, -0.5575223, -0.5924181, 
    -0.7003771, -0.8489122, -0.9403998, -0.9768583, -0.9908556, -0.9223171,
  -0.5557644, -0.4330268, -0.3314154, -0.1436884, 0.1475396, 0.1627576, 
    -0.04147446, -0.2753286, -0.2180371, -0.3746126, -0.3939643, -0.01352859, 
    -0.8066924, -1.246795, -0.6314473, -0.7358747, -0.7926612, -0.8082862, 
    -0.8185234, -0.7914243, -0.9069839, -1.023309, -1.178908, -1.189146, 
    -1.182375, -1.078583, -0.9520369, -0.7898297, -0.5454779, -0.3320999, 
    0.05107141, 0.1534966, -0.1566598, -0.2192252, -0.278275, -0.3673213, 
    -0.2926624, -0.4802766, -0.6546905, -0.7997751, -0.830863, -0.9135275, 
    -1.170738, -1.225833, -1.273473, -1.428095, -1.480911, -1.505407, 
    -1.585582, -1.400003, -1.170429, -0.9562364, -0.8620796, -0.8710964, 
    -0.8188992, -0.9461455, -1.118688, -1.294258, -1.379414, -1.202168, 
    -1.001827, -0.7604203, -0.602412, -0.4893422, -0.5231476, -0.5873244, 
    -0.5033891, -0.4352405, -0.3433948, -0.3436713, -0.4111185, -0.4645042, 
    -0.4296408, -0.3197455, -0.1459169, 0.1325815, -0.05457687, 0.1994601, 
    0.2948375, -0.1517608, 0.1700005, 0.3874809, -0.008596659, -0.05817366, 
    -0.7158728, -1.018395, -0.7566435, -0.4365752, -0.6367381, -0.5766799, 
    -0.5675979, -0.5503452, -0.5734084, -0.6380725, -0.6864774, -0.7136748,
  -0.1599631, -0.1292992, 0.05844426, 0.3964816, 0.5080864, 0.05466843, 
    -0.1123894, -0.04370451, -0.1651888, -0.3890333, -0.3203969, 0.4491346, 
    0.08663461, -0.3872757, -0.04236937, -0.1093602, -0.07947731, -0.0655942, 
    -0.1437678, -0.2782893, -0.4323096, -0.4700046, -0.550343, -0.5722184, 
    -0.5667982, -0.5103207, -0.4553728, -0.3174329, -0.164536, -0.008743525, 
    0.2185029, 0.3417616, 0.0192349, -0.1678739, -0.1686873, -0.2142611, 
    -0.2571483, -0.4966664, -0.6066117, -0.6473651, -0.7514176, -0.8397317, 
    -0.7026057, -0.7470069, -0.7099295, -0.6419125, -0.6850762, -0.5702977, 
    -0.5957861, -0.4582863, -0.4527197, -0.5085301, -0.5592303, -0.7925963, 
    -0.9111185, -0.9984231, -1.004332, -0.9739933, -0.9492211, -0.8251162, 
    -0.7266304, -0.5886583, -0.4984078, -0.3223486, -0.2279811, -0.2378597, 
    -0.2225113, -0.2495294, -0.2025571, -0.1888523, -0.1579604, -0.1171241, 
    -0.1046238, 0.1058412, 0.1887679, 0.5566216, 0.4091118, 0.08891332, 
    0.1883271, -0.2070178, 0.07581103, 0.6504692, 0.484844, 0.2859509, 
    -0.4000523, -0.9464548, -0.6160827, -0.3671253, -0.5928731, -0.5312195, 
    -0.5702167, -0.5038428, -0.4834652, -0.4946957, -0.3929868, -0.3190608,
  0.08305454, 0.08238602, 0.1798472, 0.3953095, 0.5107068, -0.1168979, 
    -0.05905271, 0.197962, -0.07018542, -0.2788281, -0.4255245, 0.09443083, 
    0.1224582, -0.3794298, -0.2125177, -0.01336432, 0.1352358, 0.250145, 
    0.309617, 0.1812325, 0.05307388, 0.03517056, -0.004655838, -0.02233219, 
    -0.06687927, -0.05809069, 0.01899242, 0.0729804, 0.06671429, 0.1665492, 
    0.1639621, 0.2705538, 0.149395, -0.03581005, -0.1256704, -0.117466, 
    -0.3172708, -0.4105983, -0.4633317, -0.5554218, -0.6133966, -0.5326676, 
    -0.3530612, -0.3125992, -0.3078465, -0.0912776, 0.000128746, -0.08276558, 
    -0.2902522, -0.306756, -0.4699397, -0.7459812, -0.9030938, -0.9852881, 
    -0.9179702, -0.7567563, -0.6024265, -0.4237156, -0.3850598, -0.4617367, 
    -0.4763851, -0.3442564, -0.196909, 0.01070786, -0.05649567, -0.03724098, 
    -0.009815693, -0.00909996, 0.0144515, 0.03946781, 0.03121614, 0.08401537, 
    0.1085758, 0.2445951, 0.158771, 0.343259, 0.3553358, -0.0298208, 
    0.1873507, -0.1766792, -0.01424432, 0.4625295, 0.4429492, 0.5884733, 
    -0.1890652, -0.7700384, -0.4200535, -0.2571468, -0.5376968, -0.3690448, 
    -0.3320651, -0.2144384, -0.1239924, -0.03567839, 0.02781439, -0.003761292,
  0.2436817, 0.2164843, 0.07564831, 0.2936167, 0.6516411, 0.1267388, 
    0.05374038, 0.4103646, 0.09247708, -0.1809597, -0.3793979, -0.1157262, 
    -0.2344747, -0.5245948, -0.109458, 0.1454902, 0.2289701, 0.4754705, 
    0.5395489, 0.4869289, 0.3626604, 0.2828598, 0.255825, 0.2424302, 
    0.2402329, 0.1934233, 0.1764798, 0.1791492, 0.1237941, 0.2113419, 
    0.2305956, 0.2060518, 0.2443658, 0.1235975, -0.001955807, -0.007473707, 
    -0.1608086, -0.3568697, -0.1424499, -0.3703642, -0.5007176, -0.5233903, 
    -0.476336, -0.1784682, 0.1236477, 0.2853336, 0.3141427, 0.1821113, 
    -0.01399899, -0.3261895, -0.4400077, -0.3676772, -0.3596859, -0.2675633, 
    -0.1329117, -0.08226061, -0.03533697, 0.1058092, 0.07097816, -0.03229332, 
    -0.1000018, -0.04282379, -0.03029156, 0.0483222, 0.06892729, 0.1899886, 
    0.1310372, 0.2255192, 0.2025375, 0.2362289, 0.2186346, 0.2293768, 
    0.2747059, 0.1599746, 0.2266407, 0.09063852, 0.06427133, -0.09507112, 
    0.02891979, 0.02148161, 0.1346652, 0.2463351, 0.3028941, 0.7712531, 
    -0.008856773, -0.4818377, -0.2445326, 0.01948071, -0.0258317, 0.01603031, 
    0.04867983, 0.1288881, 0.1886864, 0.1874661, 0.1842108, 0.1852036,
  0.211797, 0.295033, 0.163132, 0.1090469, 0.5849741, 0.05196665, -0.1233426, 
    0.4724093, 0.3839972, -0.01383734, -0.2364936, -0.0672226, -0.3542333, 
    -0.4156432, -0.01901197, 0.009097099, 0.107306, 0.3153467, 0.3528471, 
    0.4853663, 0.5378566, 0.4744616, 0.3931952, 0.3248353, 0.3444643, 
    0.2416487, 0.2294416, 0.1895652, 0.1386051, 0.2186489, 0.3325815, 
    0.1539357, 0.0234828, -0.02020168, -0.08577824, -0.1290073, -0.1919284, 
    -0.2563839, -0.02417278, 0.01705408, -0.1500523, -0.1700859, -0.192287, 
    -0.2416358, 0.07361507, 0.2542629, -0.02091599, -0.3312187, -0.4061379, 
    -0.4171405, -0.4670749, -0.3650241, -0.2761736, -0.1455746, 0.05873871, 
    0.1607242, 0.2038722, 0.1865058, 0.02828598, 0.006541729, -0.1326189, 
    -0.07828903, 0.02337074, 0.1535468, 0.1917787, 0.2539697, 0.2318993, 
    0.3108711, 0.259748, 0.2824206, 0.2549953, 0.1460109, 0.2096481, 
    0.09688807, 0.2724093, 0.1358858, -0.01343049, -0.061575, 0.028285, 
    -0.01943636, 0.04366586, 0.1327609, 0.2904269, 0.2769825, 0.1934705, 
    -0.1569357, -0.2919784, 0.0264473, 0.1342106, 0.07114077, 0.1744123, 
    0.1638656, 0.2254057, 0.2276511, 0.2684221, 0.2476041,
  0.2450494, 0.3316541, 0.2603971, 0.1866837, 0.5392394, 0.01020229, 
    -0.3848009, 0.1932427, 0.2648084, 0.2995744, -0.160305, -0.1635451, 
    -0.1959171, -0.326776, -0.3095236, -0.0767107, 0.06803131, -0.0171566, 
    0.09259272, 0.06910658, 0.2352524, 0.3971338, 0.4563298, 0.4176908, 
    0.3506331, 0.2815905, 0.4262028, 0.2308885, 0.09846675, 0.3014777, 
    0.3810027, 0.2752085, -0.02233386, -0.2594435, -0.07016921, 0.03458309, 
    0.006067991, -0.06507438, 0.005026549, 0.003122211, 0.05232406, 
    0.1016243, 0.04430032, -0.3069861, -0.2969921, -0.1231637, -0.1995475, 
    -0.2877307, -0.2768257, 0.01741314, 0.2133441, 0.3194971, 0.4146795, 
    0.4156885, 0.4127259, 0.4375801, 0.4240708, 0.3043766, 0.1316552, 
    0.1169906, 0.09129095, 0.07638216, 0.07351732, 0.2409978, 0.2944813, 
    0.2232895, 0.2296858, 0.2248359, 0.3535628, 0.2505345, 0.172946, 
    0.157191, 0.1792122, 0.04283577, 0.01612675, -0.09292328, -0.1665066, 
    0.05427783, 0.01181364, -0.08265251, -0.01989207, 0.08031949, 0.01156914, 
    0.00764668, 0.1249967, 0.1145492, -0.2991395, 0.02462387, 0.1125798, 
    0.04376459, 0.1920881, 0.189549, 0.2869925, 0.2174609, 0.2371392, 
    0.1931446,
  0.3304823, 0.226885, 0.16222, 0.1759572, 0.2882293, 0.05367565, 
    -0.06500927, 0.01121143, 0.01384814, 0.6490527, 0.1345181, -0.2721387, 
    -0.1384795, -0.4126983, -0.7339061, -0.6576371, -0.5631216, -0.4790888, 
    -0.2517126, -0.3383825, -0.1261423, 0.02154589, 0.3593554, 0.4576302, 
    0.4992156, 0.4622364, 0.2830051, 0.08163792, 0.09351933, 0.1328908, 
    0.06936572, 0.04452848, -0.02243115, -0.03623331, 0.03110075, -0.0228706, 
    -0.0336779, -0.03330355, 0.005709529, 0.09400749, -0.07005572, 
    -0.1281281, -0.02072215, 0.1415985, 0.3267874, 0.7518525, 1.089157, 
    1.287335, 1.260317, 1.126773, 0.9506168, 0.8406725, 0.7941389, 0.6963201, 
    0.6166654, 0.5947738, 0.5148258, 0.3493471, 0.1580553, 0.03141117, 
    0.06163597, 0.03447104, 0.1372871, 0.1970849, 0.2592907, 0.1516738, 
    0.1280727, 0.1128061, 0.2205207, 0.1484995, 0.1585257, -0.0159207, 
    -0.1260933, -0.1776069, -0.1117218, 0.09273791, -0.09391552, 
    -0.003437012, 0.02748747, -0.120771, 0.02214894, -0.03519154, -0.1624703, 
    -0.04536462, 0.04796267, 0.1704407, 0.1025867, 0.3773422, 0.2919908, 
    0.2262678, 0.2545383, 0.2424777, 0.3149712, 0.2384405, 0.3161592, 
    0.3104465,
  0.2489386, 0.1523731, 0.1857066, 0.1256971, 0.08189833, 0.04863012, 
    0.04417042, -0.01448844, -0.002672017, 0.5842257, 0.4682262, -0.09352517, 
    -0.2042182, -0.2991076, -0.562991, -0.7728706, -0.804267, -0.97484, 
    -0.9589546, -0.8939481, -0.7364936, -0.6713569, -0.2345568, 0.01663136, 
    0.2673475, 0.3445611, 0.041924, -0.04907504, -0.13345, -0.3919787, 
    -0.1121938, 0.0132622, -0.01372347, 0.01663135, -0.2658721, -0.422106, 
    -0.1868029, 0.06562185, 0.1576467, 0.1604619, 0.08346045, 0.09931362, 
    0.2438124, 0.5321913, 0.8404756, 1.412253, 1.659144, 1.5506, 1.574591, 
    1.386717, 1.246401, 1.156672, 1.173469, 1.139679, 1.079849, 1.011359, 
    0.9410791, 0.8218246, 0.6584783, 0.5204902, 0.3854795, 0.2786756, 
    0.4013484, 0.3195772, 0.4349582, 0.3332164, 0.2790983, 0.2087698, 
    0.1187797, 0.1540499, 0.07709683, -0.185745, -0.03473639, -0.2893262, 
    -0.3688018, -0.03709614, -0.1384142, -0.008889496, 0.01653369, 
    -0.04879835, 0.01445031, 0.04125679, -0.3566926, 0.3383121, 0.2639141, 
    0.1859198, 0.3284812, 0.4920051, 0.3860807, 0.4012177, 0.3849741, 
    0.4428843, 0.5093071, 0.5980279, 0.5518038, 0.4027965,
  -0.06387031, -0.1038115, 0.04963887, 0.2096002, 0.2279106, 0.04420298, 
    0.09937875, 0.1044569, 0.1323214, 0.1446911, 0.1282687, 0.1584608, 
    -0.1899116, -0.2322782, -0.1140492, -0.2282417, -0.3843453, -0.83319, 
    -0.9896516, -1.190709, -1.270299, -0.9445833, -0.7410513, -0.3976915, 
    -0.1269885, -0.1355497, 0.02865946, -0.1213081, -0.4982287, -0.8269887, 
    -0.5522327, -0.06214476, 0.04669321, -0.0301137, -0.5792673, -0.6603383, 
    -0.3447944, 0.06414104, 0.2622205, 0.2635877, 0.1960584, 0.1061984, 
    0.1752251, 0.3342094, 0.5077609, 0.6418751, 0.4841602, 0.5424614, 
    0.67975, 0.5066862, 0.4678354, 0.4940071, 0.5526333, 0.4844532, 
    0.4732714, 0.5005338, 0.5640917, 0.4992478, 0.2946258, 0.1371388, 
    0.08738303, 0.03767598, -0.02594674, -0.1025743, -0.002834797, 
    -0.04715446, 0.03243536, -0.06961536, -0.1429715, 0.01869822, -0.1353548, 
    -0.2867546, -0.2121289, -0.7778502, -0.3467968, 0.06300181, 0.005449772, 
    0.3971652, 0.1823052, -0.2354846, -0.1107941, -0.03410101, -0.2931657, 
    -0.3183284, -0.2009306, -0.1776075, -0.04853821, 0.08347678, 0.05973035, 
    0.1224745, 0.137953, 0.180482, 0.08360696, 0.1996059, 0.07781303, 
    0.07063526,
  0.05094129, 0.2435842, 0.4787896, 0.6066216, 0.4478651, 0.332826, 
    0.5371717, 0.282175, 0.02218148, 0.1299452, 0.4739393, 0.4352349, 
    0.1675428, 0.2291476, 0.5174286, 0.1915822, -0.2504588, -0.646325, 
    -0.8889189, -1.044827, -0.895185, -0.7291535, -1.105814, -0.6057975, 
    -0.3522, -0.502477, -0.1787791, -0.1368355, -0.3901883, -0.5679067, 
    -0.4865754, -0.212503, -0.04909158, -0.214798, -0.8021516, -0.5835319, 
    -0.3840848, -0.12484, 0.1630181, 0.1993137, 0.2000298, 0.3382948, 
    0.5504855, 0.451576, 0.4396288, 0.345293, 0.2131152, 0.3191211, 
    0.1545541, -0.276793, -0.4193716, -0.3446474, -0.2519073, -0.3578153, 
    -0.2593613, -0.1973174, -0.1145535, -0.157002, -0.3520381, -0.5403187, 
    -0.673164, -0.8828967, -1.040107, -0.9064318, -0.7885607, -0.6177925, 
    -0.4119331, -0.532783, -0.3782745, -0.2577502, -0.3703315, -0.4131701, 
    -0.7710151, -1.297464, -0.1677762, 0.01308317, -0.09809875, 0.2695279, 
    -0.3149769, -0.7314305, -0.5063653, -0.259963, -0.5728045, -0.4366069, 
    -0.3417168, -0.2942233, -0.1441598, -0.07803059, -0.09930313, 
    -0.01896429, -0.07537735, 0.1329396, 0.1410773, 0.2817513, 0.1078098, 
    0.07439506,
  0.5203586, 0.5628716, 0.6318657, 0.459551, 0.1374156, 0.1732392, 0.3016572, 
    0.007923365, 0.1990858, 0.758884, 0.663246, 0.08705771, 0.1493461, 
    0.3558401, 0.7012016, 0.7964002, 0.3592092, 0.03243518, -0.1644726, 
    -0.03984714, -0.3576039, -0.9930366, -1.140888, -0.6853055, -0.4630887, 
    -0.1788114, 0.02830127, 0.04231495, -0.06556261, -0.06486279, 0.18766, 
    0.2960421, 0.02442765, -0.3870959, -0.7364777, -0.4603217, -0.285631, 
    -0.1231147, 0.2129041, 0.4804334, 0.7625461, 0.8099256, 0.6376436, 
    0.3135383, 0.2984836, 0.3766584, 0.4226055, 0.3624821, 0.2341294, 
    0.2018375, 0.2786765, 0.3571277, 0.3951316, 0.294188, 0.2409654, 
    0.1106591, 0.0720849, 0.01163578, -0.1713557, -0.3560247, -0.4307816, 
    -0.4721713, -0.5274451, -0.5209337, -0.5577013, -0.5063667, -0.6088406, 
    -0.5182645, -0.1784045, -0.09511995, -0.108271, -0.1324246, -0.3619659, 
    -0.6930696, -0.3362322, -0.3867369, -0.4361181, -0.5291529, -0.8671246, 
    -0.699091, -0.2785826, -0.2383313, -0.272625, -0.1711116, -0.02744293, 
    0.1751451, 0.2232733, 0.3065085, 0.3560843, 0.4325168, 0.4719373, 
    0.8993785, 0.8902642, 0.6011202, 0.3399875, 0.4002088,
  0.2005341, 0.006702662, 0.1099739, 0.1538219, 0.05139637, 0.01803112, 
    0.08464837, 0.2459764, 0.4894503, 0.6319796, 0.4045708, 0.1283826, 
    0.288799, -0.05194008, -0.2131702, 0.2224417, 0.3285942, 0.3444633, 
    0.4368788, 0.4051242, -0.200019, -0.6300483, -0.1036323, 0.2371879, 
    0.2262993, 0.3698052, 0.1945609, 0.1009731, -0.003779173, 0.2600393, 
    0.6509576, 0.461195, -0.0644238, -0.3972361, -0.385501, -0.3014517, 
    -0.1024773, 0.3581187, 0.6966115, 0.8181936, 0.8278615, 0.5765917, 
    0.3662243, 0.3313627, 0.4231267, 0.3267889, 0.1642728, 0.1960435, 
    0.2913723, 0.2705388, 0.2388978, 0.1959944, 0.1088686, 0.001039982, 
    -0.131577, -0.277606, -0.3194351, -0.3637547, -0.4536147, -0.5465188, 
    -0.5029473, -0.4683943, -0.4504747, -0.4442742, -0.5645707, -0.7763214, 
    -0.6579942, -0.04162061, 0.04570037, 0.05142957, 0.1551242, -0.01548129, 
    -0.415823, -0.4464066, 0.03766012, -0.08574343, -0.1498222, -0.1900902, 
    -0.2116389, -0.06847477, 0.02958822, -0.02890778, 0.06025219, 0.09723139, 
    0.2026839, 0.2887192, 0.2474918, 0.4443669, 0.5166326, 0.6855931, 
    0.8950486, 1.221384, 0.6279757, 0.2010061, 0.1905731, 0.2732229,
  0.03995466, -0.3018262, -0.296097, -0.1198926, -0.0555861, 0.1370409, 
    0.3390594, 0.495928, 0.6015598, 0.5780734, 0.7860484, 0.3717581, 
    -0.0364933, -0.2984891, -0.6518094, -0.5055044, -0.2405952, -0.3450548, 
    -0.2909044, -0.2030302, -0.1263862, 0.01825893, 0.393145, 0.7496223, 
    0.6352837, 0.2622206, -0.008889496, 0.1227511, -0.004397631, 0.06954467, 
    0.210886, -0.03667164, -0.1777849, -0.2201838, -0.003549576, 0.1234522, 
    0.2736793, 0.5072887, 0.5157354, 0.4368455, 0.3573213, 0.3606591, 
    0.5156074, 0.4905748, 0.3968406, 0.2896309, 0.2150702, 0.3145165, 
    0.2972636, 0.1867499, 0.2133126, 0.2919583, 0.2314115, 0.1369123, 
    -0.06684732, -0.2331395, -0.2245622, -0.2630553, -0.3437352, -0.3618178, 
    -0.3759785, -0.5196958, -0.4639668, -0.2306023, -0.1713088, -0.1791048, 
    0.2042289, 0.3869439, 0.02496469, 0.2194958, 0.1334932, -0.4256375, 
    -0.7907907, -0.5676138, -0.07758951, -0.0657897, -0.03872252, 0.1526022, 
    0.239419, 0.150373, 0.1839995, 0.2087226, 0.1772118, 0.1653957, 
    0.1784325, 0.2185693, 0.365428, 0.4977365, 0.5033841, 0.6930971, 
    0.7112284, 0.8529429, 0.1681443, -0.1195834, 0.09071922, 0.1824348,
  -0.2364125, -0.6657746, -0.7503128, -0.4577508, -0.3692741, 0.06026697, 
    0.405547, 0.3743293, 0.5946913, 0.5608534, 0.7135874, 0.4963835, 
    -0.07306647, -0.1710965, -0.4171903, -0.4236032, -0.3550483, -0.5749865, 
    -0.4925971, -0.1733426, 0.07677133, 0.03608125, 0.3639295, 0.3468885, 
    0.05242237, 0.02325571, -0.1166857, 0.02996135, 0.1081512, -0.01876926, 
    -0.05926418, -0.03550124, 0.09945965, 0.1771307, 0.2759748, 0.4832182, 
    0.6158023, 0.4390931, 0.2052398, 0.1389799, 0.3356428, 0.5130353, 
    0.4048328, 0.2533841, 0.2130032, 0.2613754, 0.4108543, 0.4451485, 
    0.2924466, 0.245718, 0.2106595, 0.05021, -0.222414, -0.4008317, 
    -0.6018405, -0.6948256, -0.5196142, -0.4038429, -0.3921561, -0.3766942, 
    -0.3049006, -0.2333841, -0.108808, 0.04972005, 0.3052216, 0.6500949, 
    0.8499159, 0.5074517, 0.2246386, 0.2404914, -0.3284695, -0.9437691, 
    -0.6822295, -0.2969093, -0.1492205, -0.1735206, 0.0675106, 0.2371721, 
    0.3235002, 0.4075816, 0.513978, 0.4502738, 0.3435521, 0.2929344, 
    0.2139297, 0.2063289, 0.2747378, 0.2899723, 0.2700667, 0.3176579, 
    0.2073388, 0.2376599, -0.1715851, -0.3525259, -0.2732613, -0.203356,
  -0.4550974, -0.6233597, -0.5048213, -0.1885612, -0.08325505, 0.2826304, 
    0.5191053, 0.3795871, 0.5173963, 0.3255832, 0.1767063, 0.1756154, 
    -0.08444285, -0.1011421, -0.1715034, -0.1762398, 0.03871799, -0.06256786, 
    -0.1633003, 0.09900415, 0.1033826, -0.1459991, 0.3332492, 0.1496066, 
    -0.04529929, 0.2489718, -0.07619119, 0.06710336, 0.363636, 0.08360672, 
    0.1549771, 0.257858, 0.265769, 0.3567367, 0.3542304, 0.4914699, 
    0.4202781, 0.1814923, 0.06012249, -0.09630728, 0.1238256, 0.353579, 
    0.1708636, 0.1276178, 0.3020649, 0.3464003, 0.3552389, 0.3125148, 
    0.2691069, 0.2710919, 0.1481919, -0.002328873, -0.2440286, -0.4601579, 
    -0.5849466, -0.5836773, -0.4507184, -0.3749371, -0.2864442, -0.119534, 
    0.04304695, 0.117233, 0.1808236, 0.3252577, 0.5741184, 0.6832327, 
    0.6567193, 0.6256318, 0.4277639, -0.1320671, -0.4619006, -0.3356965, 
    -0.08221149, -0.005520344, -0.07967472, -0.05177689, 0.07135153, 
    0.07408524, 0.01547527, -0.04770875, -0.1066442, -0.1811721, -0.1745479, 
    -0.1382358, -0.07832384, -0.03244162, -0.04515314, 0.02906585, 
    -0.03917909, -0.1443713, -0.2105656, -0.3085639, -0.3228056, -0.3367378, 
    -0.2269396, -0.2645867,
  -0.02392852, 0.195814, 0.2481414, 0.0738579, 0.01049483, 0.0393852, 
    0.1465304, 0.2245903, 0.4510227, 0.2169406, -0.05511338, -0.09531528, 
    -0.2364285, -0.0819038, -0.010631, -0.0835802, 0.03403044, 0.02434623, 
    -0.1683296, -0.01154244, -0.05975211, -0.2803257, -0.03802395, 
    -0.3249707, -0.4812369, -0.5094428, -0.6855321, 0.03331429, 0.1026497, 
    -0.2256864, 0.000859499, 0.1452441, 0.2358693, 0.45278, 0.3869433, 
    0.4365852, 0.3036752, 0.0983696, 0.1090956, 0.05178785, -0.01051784, 
    -0.1306348, -0.2775753, -0.1889679, -0.03206706, 0.1023407, 0.1440237, 
    0.1439424, 0.1575816, 0.05377293, -0.1275909, -0.300703, -0.4670278, 
    -0.5466174, -0.5963569, -0.6383979, -0.5848498, -0.501842, -0.3493518, 
    -0.03063464, 0.2844371, 0.4106089, 0.5300591, 0.6786431, 0.7403615, 
    0.6725559, 0.7345675, 0.770521, 0.312448, -0.419111, -0.4130561, 
    -0.1073271, -0.06338167, -0.009084821, 0.007614493, 0.09031224, 
    0.09285164, -0.02345729, -0.1748897, -0.2752308, -0.3559273, -0.5375679, 
    -0.6011746, -0.5014187, -0.3468614, -0.2243842, -0.1450873, -0.04883146, 
    -0.1299675, -0.1482129, -0.2157094, -0.4105499, -0.3962107, -0.3699574, 
    -0.1770535, -0.003388166,
  0.005319506, -0.07908805, -0.3199897, -0.4705106, -0.1067248, -0.1008491, 
    0.06449917, 0.3214002, 0.08790362, -0.181562, -0.2454129, -0.1687853, 
    -0.1706082, -0.1807972, -0.2121609, -0.2516792, -0.1511909, 0.03570688, 
    -0.08050407, -0.09272736, -0.04700828, 0.01545894, 0.1089817, 0.0949676, 
    0.1029427, 0.07004881, 0.233965, 0.4199353, -0.107002, -0.4069689, 
    -0.16457, -0.2530789, -0.1638536, -0.04502261, -0.2449572, -0.2569366, 
    -0.07697219, -0.05366487, -0.2003934, -0.2082549, -0.06999004, 
    -0.06481421, -0.02407539, 0.02151406, -0.0947293, -0.2390327, -0.398896, 
    -0.5433296, -0.7304227, -0.9329293, -1.019013, -1.035306, -1.020283, 
    -0.9094107, -0.8108594, -0.6620151, -0.3946486, -0.1239942, 0.05058289, 
    0.2155569, 0.3602836, 0.411016, 0.4676239, 0.5196587, 0.4693657, 
    0.5744113, 0.5740694, 0.5171522, 0.3418427, 0.0696913, -0.0184598, 
    -0.1229194, -0.1889839, -0.1216173, -0.08688429, -0.04591748, 0.05740283, 
    0.07561573, 0.1032036, 0.01288787, -0.156269, -0.3750842, -0.4358589, 
    -0.3074573, -0.1721544, -0.1102729, -0.0333198, -0.01048452, -0.04419222, 
    0.07693408, 0.02690157, -0.0119819, 0.07932663, -0.03825152, 0.09322643, 
    0.2273898,
  -0.2526557, -0.6803576, -0.9469591, -0.7960804, -0.4406115, -0.4720894, 
    -0.2818061, -0.2812364, -0.4861844, -0.5266303, -0.4894233, -0.5107449, 
    -0.6044461, -0.5600454, -0.3726107, -0.2684438, -0.05623657, 0.1360155, 
    0.09182668, 0.2704399, 0.645895, 0.4483859, 0.1214165, 0.1192355, 
    0.4251437, 0.3504366, 0.4714002, 0.3451145, -0.2472195, -0.4582872, 
    -0.428258, -0.4302114, -0.2646024, -0.2792997, -0.448066, -0.714635, 
    -0.6162952, -0.2635772, -0.2162306, -0.1805534, -0.001679778, 0.2007781, 
    0.3238416, 0.3358045, 0.2221975, 0.03083992, -0.2043977, -0.4410348, 
    -0.7528837, -1.060631, -1.156155, -1.127704, -1.029641, -0.9102235, 
    -0.7674661, -0.4677916, -0.147397, 0.08792114, 0.2594218, 0.4275208, 
    0.577976, 0.5822401, 0.433249, 0.2025363, 0.2124321, 0.3234185, 0.232826, 
    0.2628876, 0.2137501, 0.0347954, -0.1479683, -0.2042021, -0.117353, 
    -0.05480421, -0.0855664, -0.01689768, 0.02262092, -0.03826785, 0.0242641, 
    0.1733363, 0.3406382, 0.4269176, 0.3690884, 0.2743948, 0.1992483, 
    0.1247528, 0.09412098, 0.1300914, 0.2159312, 0.3467091, 0.4265754, 
    0.4623182, 0.4421197, 0.3563287, 0.3907036, 0.2348768,
  -0.3836128, -0.5511747, -0.4543325, -0.3083687, -0.3510933, -0.5252469, 
    -0.4776883, -0.4629585, -0.4945503, -0.2985542, -0.1631212, -0.2931505, 
    -0.2477079, -0.0234077, -0.008368969, 0.005628228, 0.07732439, 0.1465305, 
    0.1922498, 0.2484673, 0.3581027, -0.0117377, -0.2109566, -0.09329703, 
    -0.1314968, -0.3286324, -0.2463572, -0.2701693, -0.3979522, -0.4469596, 
    -0.4063344, -0.3720572, -0.523473, -0.7056179, -0.572659, -0.3216991, 
    -0.5679388, -0.6267915, -0.3397005, -0.2410021, -0.1114111, 0.1150694, 
    0.2955379, 0.334568, 0.2562318, 0.1091619, -0.002150059, -0.0916357, 
    -0.2765474, -0.4290218, -0.4725761, -0.5238461, -0.561883, -0.5091162, 
    -0.3952813, -0.2277036, -0.05577946, 0.1265936, 0.366209, 0.5184231, 
    0.5975246, 0.5566387, 0.3380501, 0.1402317, 0.2457981, 0.2727346, 
    0.2502085, 0.2336719, 0.08608103, -0.2243524, -0.3463898, -0.255358, 
    -0.07099915, -0.02715182, -0.07213879, -0.0279007, -0.06292629, 
    -0.08638024, -0.1448438, -0.08001614, 0.06026697, 0.2568977, 0.4256644, 
    0.5898409, 0.6900356, 0.6478162, 0.5487602, 0.4756963, 0.5067024, 
    0.589401, 0.6115038, 0.5922334, 0.5391078, 0.4335585, 0.2627739, 
    -0.03859323,
  -0.4923042, -0.4750841, -0.3621122, -0.2729357, -0.5197619, -0.6525908, 
    -0.4633495, -0.2285184, -0.2094755, -0.2244493, -0.3049181, -0.3510932, 
    -0.2053576, -0.09884715, -0.03751904, 0.06891, 0.2023735, 0.2070448, 
    0.09664437, 0.04098031, 0.06402719, -0.01037061, -0.06644157, 
    -0.03992787, -0.1563992, -0.2613801, -0.2583206, -0.3125355, -0.365335, 
    -0.3046091, -0.3646677, -0.4886589, -0.6005387, -0.6050973, -0.3390496, 
    -0.1619012, -0.3558784, -0.6251645, -0.6412125, -0.5217304, -0.4269547, 
    -0.3140478, -0.2328138, -0.1493506, -0.04425573, 0.04959154, 0.1332507, 
    0.1481919, 0.08193207, 0.0349431, 0.01583576, -0.06782341, -0.115447, 
    -0.02021694, 0.1557598, 0.2530575, 0.3164854, 0.4777164, 0.6130843, 
    0.6174955, 0.5945458, 0.5815415, 0.47874, 0.3070773, 0.2923312, 
    0.2435842, 0.1799779, 0.08502436, -0.1232762, -0.2627959, -0.2390659, 
    -0.2467477, -0.2642934, -0.1588087, -0.07654953, -0.08138299, 
    -0.09414351, -0.05128884, -0.08890319, -0.1442573, -0.2237983, 
    -0.2232442, -0.1094103, 0.1893044, 0.4339824, 0.507648, 0.4203434, 
    0.3409166, 0.3933253, 0.4774232, 0.4035463, 0.2859192, 0.1874332, 
    0.04897141, -0.1424994, -0.2991402,
  -0.4509959, -0.5100615, -0.450573, -0.3543813, -0.3441598, -0.2102406, 
    -0.06868792, -0.01160777, -0.01548135, -0.1201199, -0.3017117, 
    -0.3641792, -0.2599149, -0.1514839, -0.03214788, 0.1550916, 0.2426078, 
    0.154359, 0.02794302, 0.05780911, 0.0640105, -0.03678656, -0.160338, 
    -0.2794139, -0.3050816, -0.2418981, -0.2399774, -0.2748892, -0.2655306, 
    -0.2154977, -0.2910352, -0.3901064, -0.2375033, -0.1817579, -0.2700229, 
    -0.205162, -0.1581573, -0.2352736, -0.2513361, -0.2847185, -0.2705903, 
    -0.300571, -0.3172545, -0.2271175, -0.05185699, 0.1338525, 0.3482895, 
    0.5822411, 0.7438297, 0.8182111, 0.8499985, 0.8878565, 0.8855619, 
    0.8094382, 0.6935372, 0.6589499, 0.76092, 0.8633771, 0.817121, 0.6794744, 
    0.5689111, 0.4993293, 0.2812961, 0.1858533, 0.1270314, 0.09040999, 
    0.07299662, -0.0131855, -0.147902, -0.1750846, -0.1583204, -0.1528351, 
    -0.1203156, -0.04349279, -0.02269185, -0.05635047, -0.08398736, 
    -0.09341133, -0.08229482, -0.05299807, -0.01235676, -0.05071926, 
    -0.1376333, -0.05161285, 0.06533051, 0.1152983, 0.03176928, -0.03947115, 
    0.04584789, 0.1786766, 0.1835432, 0.04542494, -0.1827002, -0.3872905, 
    -0.4529161, -0.4382839,
  -0.8424025, -0.9365914, -0.737715, -0.5964386, -0.4438019, -0.2480662, 
    -0.07508445, 0.027601, 0.04788113, -0.03086233, -0.1490754, -0.1863149, 
    -0.09800112, -0.009231567, 0.01220405, 0.03251648, 0.04140258, 
    -0.003128529, -0.06432629, -0.06268215, -0.05403972, -0.1278031, 
    -0.1924677, -0.2053578, -0.2866566, -0.3084016, -0.3471062, -0.3633335, 
    -0.341198, -0.3213577, -0.3720899, -0.1925969, -0.03437829, 0.0391407, 
    0.0549283, 0.1273079, 0.2271938, 0.1807585, 0.2533998, 0.4942365, 
    0.6720178, 0.6577275, 0.4852183, 0.6446748, 0.7304814, 0.7990859, 
    0.8666804, 0.974607, 1.055092, 1.077342, 1.046402, 0.9952621, 0.8638167, 
    0.6838036, 0.5601382, 0.5792136, 0.6616359, 0.5988107, 0.3726387, 
    0.209177, 0.2745574, 0.3348443, 0.2966932, 0.2108696, 0.08546209, 
    -0.07697248, -0.1636586, -0.1763377, -0.08286476, -0.000670433, 
    0.03044951, 0.06977224, 0.1734669, 0.2466602, 0.1793101, 0.09128928, 
    0.01980495, -0.03188777, -0.05509734, 0.0287075, 0.110153, 0.02511072, 
    0.04721403, 0.08168745, 0.06791782, -0.03882027, -0.176743, -0.187078, 
    -0.04780436, 0.05245638, 0.003465176, -0.2087746, -0.5132017, -0.7431672, 
    -0.7711134, -0.81706,
  -1.105716, -0.9249706, -0.6848501, -0.4084501, -0.3168976, -0.2746942, 
    -0.193135, -0.06723964, -0.01124954, -0.009703636, -0.05114257, 
    0.003756762, 0.1009084, 0.1340137, 0.06039715, 0.01023459, 0.008020639, 
    0.03857064, 0.101429, 0.1613247, 0.1953905, 0.1721482, 0.1261034, 
    0.047328, -0.02287054, -0.07431984, -0.1056187, -0.04575491, 0.009551048, 
    0.03476214, 0.1846819, 0.2993307, 0.1908174, 0.147913, 0.1551723, 
    0.3071904, 0.3263638, 0.4681768, 0.9099419, 1.371937, 1.515459, 1.381019, 
    1.186488, 1.14474, 1.44487, 1.469219, 1.350258, 1.109063, 0.8620741, 
    0.6615858, 0.5272759, 0.4089164, 0.3051401, 0.2654266, 0.3046355, 
    0.3995576, 0.439857, 0.396856, 0.2971489, 0.2914196, 0.3722464, 0.363246, 
    0.224102, 0.04685569, -0.1216502, -0.1360707, -0.08232701, 0.03765976, 
    0.1956841, 0.2772923, 0.2505178, 0.3858366, 0.6118779, 0.8099411, 
    0.7604787, 0.4820933, 0.24806, 0.00701189, -0.0369339, 0.2329719, 
    0.1367643, 0.2055304, 0.1415329, -0.03504586, -0.2328482, -0.4517775, 
    -0.5868359, -0.5856805, -0.5497262, -0.5635126, -0.7172234, -0.9351761, 
    -1.131888, -1.234834, -1.216751, -1.090124,
  -0.5409375, -0.4584991, -0.313382, -0.167158, -0.01523769, 0.178447, 
    0.2519499, 0.2889132, 0.2165989, 0.1433402, 0.1327119, 0.1499484, 
    0.1547824, 0.1237766, 0.1310682, 0.1622853, 0.2510875, 0.3499806, 
    0.3568003, 0.3158166, 0.2270315, 0.1543264, 0.1255504, 0.1085584, 
    0.1081027, 0.1728977, 0.1711396, 0.1576304, 0.1361947, 0.1092577, 
    0.09706759, 0.1179333, 0.04351854, 0.04307961, 0.1283987, 0.2804494, 
    0.338913, 0.5351373, 0.7339654, 0.899232, 0.9588348, 0.8428355, 
    0.7356575, 0.6019177, 0.5221815, 0.4405569, 0.3809375, 0.3636525, 
    0.2650034, 0.09778309, -0.06780899, -0.1347848, -0.1045438, -0.03779566, 
    0.03918999, 0.2162082, 0.4084117, 0.4917613, 0.4548634, 0.2983208, 
    0.1833794, 0.06632215, -0.03126931, -0.07861638, -0.03135037, 0.1096164, 
    0.2627577, 0.3350233, 0.4358045, 0.5176243, 0.5401991, 0.5273899, 
    0.505287, 0.4024549, 0.264369, 0.1533176, 0.129994, 0.1958794, 0.2140107, 
    0.2210097, 0.1808727, 0.07201871, -0.0903185, -0.2066597, -0.2556017, 
    -0.5131701, -0.6414742, -0.6709177, -0.6875193, -0.7582549, -0.830488, 
    -0.8806508, -0.8801136, -0.8279002, -0.7122915, -0.6120474,
  0.3122206, 0.4882294, 0.611846, 0.6619105, 0.6717412, 0.6763479, 0.6193169, 
    0.4787083, 0.3540989, 0.3251599, 0.3498667, 0.4022757, 0.4072723, 
    0.4212372, 0.4433237, 0.4906708, 0.492559, 0.5010388, 0.3922985, 
    0.3126923, 0.2290497, 0.1657196, 0.1637993, 0.1468233, 0.1707979, 
    0.1974745, 0.2474093, 0.2650523, 0.2243621, 0.2967086, 0.3021454, 
    0.3225068, 0.3938775, 0.414662, 0.4363742, 0.4845676, 0.5107394, 
    0.5716118, 0.6157036, 0.6358209, 0.6814751, 0.534828, 0.355645, 
    0.1492485, 0.07040727, 0.1243787, 0.2531383, 0.3346163, 0.2463188, 
    -0.009345174, -0.2510444, -0.2971708, -0.1834989, -0.002639771, 
    0.1090624, 0.1206346, 0.07555008, 0.07312548, 0.1598604, 0.2440076, 
    0.1983208, 0.2631971, 0.3615858, 0.5172987, 0.6077446, 0.5930961, 
    0.5108371, 0.5205539, 0.5171034, 0.3994113, 0.1292615, -0.2142442, 
    -0.4505073, -0.4844754, -0.4056668, -0.1737981, 0.01218802, -0.07962516, 
    -0.1037788, -0.2275907, -0.2588732, -0.1232941, -0.1484087, 0.05569386, 
    -0.02275705, -0.06802106, 0.1926563, 0.2789681, 0.3786423, 0.3627574, 
    0.232744, 0.03925478, -0.1289741, -0.1829129, -0.08646119, 0.1064588,
  0.9225233, 0.9954075, 1.016387, 1.013181, 0.9902316, 0.9108534, 0.7997206, 
    0.6606092, 0.5497369, 0.4990044, 0.5055307, 0.5354462, 0.559258, 
    0.5892385, 0.628643, 0.5926405, 0.5413219, 0.4117156, 0.2710581, 
    0.1857554, 0.1736785, 0.136309, 0.1403131, 0.1359348, 0.1593559, 
    0.1253228, 0.1161916, 0.1640921, 0.2053353, 0.2035776, 0.2265272, 
    0.3042128, 0.4411757, 0.5470839, 0.5334445, 0.6780572, 0.8383433, 
    0.939955, 1.076087, 1.12669, 1.077845, 0.923858, 0.7907687, 0.652162, 
    0.6203748, 0.6765109, 0.6148248, 0.313897, -0.1289253, -0.4185575, 
    -0.657506, -0.4292185, -0.05006838, 0.4234829, 0.5002577, 0.4512339, 
    0.312757, 0.2092741, 0.2186007, 0.448386, 0.6090304, 0.6020963, 
    0.5262989, 0.4239227, 0.2758433, 0.1454881, 0.0112114, -0.1863309, 
    -0.4270046, -0.6430365, -0.8852892, -0.8656927, -0.7004747, -0.6024603, 
    -0.3337919, -0.423489, -0.3584989, -0.4215197, -0.5595242, -0.5754585, 
    -0.3048042, 0.1235156, 0.08053088, 0.1616828, 0.04431629, -0.09778953, 
    -0.1364774, -0.01592074, 0.144854, 0.1857069, 0.3175265, 0.3375133, 
    0.343682, 0.394382, 0.5729139, 0.7785291,
  0.4426728, 0.5022108, 0.5517714, 0.5940729, 0.6278782, 0.6463839, 0.64627, 
    0.625697, 0.5897758, 0.5789849, 0.6109185, 0.6781874, 0.7498345, 
    0.7898409, 0.7979138, 0.6188287, 0.5248019, 0.4242323, 0.315199, 
    0.2314425, 0.1801079, 0.1359673, 0.1687147, 0.2058403, 0.2112277, 
    0.1540011, 0.1194471, 0.07364631, 0.02960336, 0.08320034, 0.2325491, 
    0.4316376, 0.6545708, 0.8082327, 0.9887339, 1.211781, 1.43683, 1.581573, 
    1.387009, 1.329164, 1.061862, 0.8945122, 0.7003065, 0.5641736, 0.4552544, 
    0.3630343, 0.1561007, -0.1426134, -0.4924506, -0.8080106, -1.004479, 
    -0.9503611, -0.7282751, -0.4183629, -0.2729034, -0.2693715, -0.3622589, 
    -0.5186393, -0.5693715, -0.5722523, -0.5797887, -0.564424, -0.5542843, 
    -0.2794304, -0.3477407, -0.4546742, -0.5975454, -0.7452177, -0.8313016, 
    -0.819453, -0.7385769, -0.6000516, -0.5465196, -0.3304064, -0.3337592, 
    -0.3937691, -0.4575223, -0.7563992, -0.7185737, -0.5189155, -0.2212436, 
    -0.2667513, -0.123831, -0.2776077, -0.4507517, -0.572952, -0.7311878, 
    -0.7964387, -0.6471062, -0.5816276, -0.4865589, -0.2171578, -0.1615587, 
    -0.03074813, 0.1701957, 0.3438448,
  -0.04116511, 0.2138476, 0.4018035, 0.5316541, 0.5945935, 0.5917616, 
    0.4660778, 0.3816047, 0.3364389, 0.3266083, 0.2628547, 0.3619921, 
    0.4140267, 0.3951793, 0.3382783, 0.2481743, 0.1786593, 0.1573866, 
    0.1275688, 0.1412733, 0.1944797, 0.3018202, 0.4928358, 0.5696424, 
    0.6044569, 0.6770154, 0.7352837, 0.7948216, 0.8380669, 0.837481, 
    0.9060845, 0.8948377, 0.842852, 0.8051405, 0.7575493, 0.7100233, 
    0.6559868, 0.5980604, 0.5058241, 0.4371555, 0.3207492, 0.2040012, 
    0.08035207, -0.007343233, -0.05944282, -0.08118761, -0.1144233, 
    -0.1607612, -0.2152859, -0.2488472, -0.2527371, -0.2378609, -0.2005562, 
    -0.1627635, -0.1513053, -0.1434766, -0.1601433, -0.1997752, -0.2402213, 
    -0.2694204, -0.3304229, -0.3710643, -0.4383984, -0.4795603, -0.5691111, 
    -0.6914907, -0.6845896, -0.6542184, -0.5829129, -0.4840522, -0.369713, 
    -0.2196153, -0.1226753, -0.09822863, -0.05859649, -0.2530463, -0.4460315, 
    -0.4023149, 0.001966238, 0.0400033, -0.02684164, -0.13555, -0.2753611, 
    -0.3202993, -0.2627306, -0.3172882, -0.4683948, -0.5337095, -0.4581723, 
    -0.5195985, -0.5351431, -0.6105661, -0.5119007, -0.6071642, -0.5646186, 
    -0.4361518,
  -0.04370391, 0.01842141, 0.08206069, 0.1487275, 0.3883758, 0.3479624, 
    0.3474253, 0.207549, 0.2369601, 0.2925916, 0.3431776, 0.3811984, 
    0.3960095, 0.4017876, 0.3929985, 0.397572, 0.390899, 0.4144341, 
    0.4010714, 0.4255832, 0.478643, 0.5521945, 0.6648898, 0.7710747, 
    0.8294406, 0.7866184, 0.758298, 0.6970348, 0.6476535, 0.6063612, 
    0.5446261, 0.4560845, 0.3718397, 0.3048963, 0.242022, 0.1743136, 
    0.1145318, 0.08004284, 0.05393612, 0.03137743, 0.00678435, -0.01243767, 
    -0.04451773, -0.07360303, -0.1005562, -0.109687, -0.09306917, -0.079202, 
    -0.06282827, -0.04743117, -0.03234321, -0.03050405, -0.0420112, 
    -0.05757105, -0.06538361, -0.05218369, -0.07428658, -0.1151395, 
    -0.1719428, -0.2452013, -0.3014187, -0.341881, -0.3830593, -0.4057156, 
    -0.4123888, -0.4368353, -0.437991, -0.4311225, -0.3989285, -0.3369981, 
    -0.2268419, -0.1914579, -0.09489238, -0.08844686, 0.02245808, 0.07192075, 
    0.1202281, 0.1426077, 0.09376323, 0.01982141, -0.05771762, -0.1924181, 
    -0.2563342, -0.2735221, -0.2817581, -0.2451363, -0.2752953, -0.2478528, 
    -0.2277045, -0.1883008, -0.1655304, -0.2350942, -0.191051, -0.1972196, 
    -0.152786, -0.07944608,
  0.2375786, 0.268438, 0.3130506, 0.331996, 0.3370904, 0.3551568, 0.3618951, 
    0.3710259, 0.381231, 0.394024, 0.4045057, 0.4296522, 0.4631156, 
    0.4904758, 0.5090955, 0.5283175, 0.5503553, 0.5710585, 0.5951307, 
    0.6051078, 0.6182589, 0.6300102, 0.6382948, 0.6378552, 0.6161268, 
    0.5643202, 0.4980278, 0.4216769, 0.3398573, 0.2490044, 0.1826633, 
    0.1241346, 0.06827524, 0.01329476, -0.02654898, -0.06035432, -0.08445916, 
    -0.1017931, -0.1145047, -0.1247424, -0.1229845, -0.1201525, -0.1235868, 
    -0.1263537, -0.1270535, -0.1295275, -0.1454943, -0.1563179, -0.1740913, 
    -0.2042996, -0.2284207, -0.2399279, -0.2497912, -0.2664253, -0.3014839, 
    -0.3364285, -0.3659695, -0.3762397, -0.3885932, -0.3955757, -0.4001981, 
    -0.4011095, -0.3827176, -0.3502631, -0.3070991, -0.262226, -0.2130561, 
    -0.1703641, -0.1334988, -0.1006212, -0.06518829, -0.0306505, 
    -0.0004096031, -0.002102315, -0.03877228, -0.05379507, -0.08467072, 
    -0.1083198, -0.1169787, -0.09360626, -0.04940051, -0.04023719, 
    -0.07581663, -0.07462895, -0.008580804, 0.03396475, 0.05271482, 
    0.0305469, 0.03637385, -0.0102241, 0.004001141, 0.03197956, 0.05463594, 
    0.09417041, 0.1380506, 0.1846489,
  0.6043267, 0.5932915, 0.6053358, 0.5982883, 0.5976861, 0.5856417, 0.581589, 
    0.5783175, 0.5761203, 0.5769666, 0.5831352, 0.5776014, 0.5627414, 
    0.5694308, 0.5722466, 0.5639784, 0.5504041, 0.5308729, 0.5131482, 
    0.4894178, 0.4549451, 0.4113253, 0.3678195, 0.3178846, 0.2655571, 
    0.2086398, 0.1522108, 0.1007785, 0.03681365, -0.02698845, -0.08567984, 
    -0.1527534, -0.2145535, -0.276549, -0.3259793, -0.3702176, -0.4079129, 
    -0.4369656, -0.4604683, -0.4794787, -0.495299, -0.5099311, -0.5159696, 
    -0.5100288, -0.511217, -0.5246772, -0.5280952, -0.5189155, -0.5062528, 
    -0.4929227, -0.492353, -0.484215, -0.4759305, -0.4665555, -0.4609891, 
    -0.4518582, -0.4419461, -0.4323758, -0.4088244, -0.3856473, -0.3553413, 
    -0.326728, -0.2934598, -0.2568387, -0.2119982, -0.1623237, -0.1122912, 
    -0.06435822, -0.01323518, 0.03253303, 0.07196988, 0.1089165, 0.1428195, 
    0.1734999, 0.2047661, 0.2360812, 0.2619764, 0.2884412, 0.3207817, 
    0.3485975, 0.374981, 0.3971326, 0.4175591, 0.4399224, 0.4586886, 
    0.4762505, 0.4919569, 0.5048963, 0.5196261, 0.5330701, 0.5498833, 
    0.569675, 0.5769503, 0.5886691, 0.5915827, 0.6031548,
  -0.1608423, -0.1513534, -0.1397485, -0.1265161, -0.1119003, -0.09603116, 
    -0.08024339, -0.06522062, -0.05088151, -0.03950435, -0.03004813, 
    -0.02293527, -0.01954985, -0.01756406, -0.01885009, -0.02231669, 
    -0.02859926, -0.03779531, -0.04975867, -0.06260037, -0.07633734, 
    -0.08961868, -0.1007357, -0.108825, -0.116735, -0.1221552, -0.1247587, 
    -0.122545, -0.1184273, -0.1100776, -0.09959579, -0.08528852, -0.06772685, 
    -0.04796791, -0.02676022, -0.004868984, 0.01591539, 0.03490961, 
    0.05180413, 0.0660457, 0.07725978, 0.08438885, 0.08756268, 0.08824635, 
    0.08658624, 0.08100319, 0.07488275, 0.07104158, 0.06386399, 0.03687835, 
    0.04176188, 0.02743864, -0.004300117, 0.04304743, 0.05040359, 0.03792, 
    0.03785515, 0.05160809, 0.05068016, 0.05627966, 0.06288815, 0.08319974, 
    0.1116507, 0.1192677, 0.1297007, 0.1384244, 0.1476855, 0.1465135, 
    0.1541796, 0.1632779, 0.1651177, 0.1627576, 0.1514456, 0.1473284, 
    0.121856, 0.1215789, 0.09120822, 0.08450174, 0.07278323, 0.05116844, 
    0.03279352, 0.01350641, -0.006953239, -0.02791691, -0.0495801, 
    -0.07052755, -0.08996105, -0.107311, -0.123131, -0.1371615, -0.1492708, 
    -0.1591668, -0.1657259, -0.1696148, -0.1703148, -0.1667829,
  -0.4257349, -0.4167994, -0.3892766, -0.3430526, -0.2857935, -0.2219915, 
    -0.1606308, -0.1031764, -0.05089772, -0.008742809, 0.02514398, 
    0.05497795, 0.08183336, 0.1055476, 0.126739, 0.1441544, 0.1569961, 
    0.1676081, 0.1770808, 0.1849747, 0.188881, 0.1887834, 0.1855282, 
    0.1765277, 0.1613908, 0.1432595, 0.1191547, 0.08285856, 0.03971076, 
    -0.00524354, -0.04759407, -0.08011341, -0.09987259, -0.1056669, 
    -0.09904265, -0.08180618, -0.05724502, -0.02897358, 0.0002417564, 
    0.02631581, 0.04594475, 0.05497795, 0.04500073, 0.01166737, -0.01255119, 
    -0.02708578, -0.07521391, -0.1022971, -0.1343122, -0.1402042, -0.1559267, 
    -0.1710808, -0.1649764, -0.1738641, -0.1563827, -0.1891472, -0.1883497, 
    -0.1876659, -0.206579, -0.2138054, -0.2347357, -0.2364442, -0.2257185, 
    -0.1875672, -0.1300806, -0.05597579, 0.04369867, 0.1616023, 0.2718074, 
    0.3784969, 0.4567032, 0.5011855, 0.5082982, 0.5353001, 0.4633764, 
    0.4279597, 0.4001928, 0.3723444, 0.3235653, 0.3141576, 0.3462867, 
    0.3282202, 0.362058, 0.3422991, 0.355906, 0.3123837, 0.2634091, 
    0.1893206, 0.1044247, 0.01147223, -0.08161044, -0.1718612, -0.2535994, 
    -0.3232608, -0.3781437, -0.4127142,
  -0.2960636, -0.3344915, -0.3423528, -0.3311874, -0.313593, -0.2964706, 
    -0.2759465, -0.2502468, -0.2120305, -0.1712753, -0.1431829, -0.1339543, 
    -0.1336451, -0.1328313, -0.1349635, -0.1415225, -0.1555363, -0.1721213, 
    -0.1822126, -0.1795108, -0.1582379, -0.1208357, -0.06671786, 0.003464252, 
    0.08071038, 0.1554337, 0.2228491, 0.2774878, 0.3089982, 0.3179663, 
    0.3082008, 0.2842588, 0.2482882, 0.206768, 0.1652806, 0.1279917, 
    0.09721422, 0.07161188, 0.04985094, 0.04023123, 0.03899407, 0.04467511, 
    0.07380939, 0.08045006, 0.07138437, 0.05797267, 0.03049879, 
    -0.0005884469, -0.04393157, -0.0959335, -0.1374375, -0.1539902, 
    -0.1453477, -0.1335638, -0.1199406, -0.1136093, -0.1075547, -0.135875, 
    -0.1901392, -0.2646185, -0.3426621, -0.4217961, -0.4904322, -0.5214056, 
    -0.5064803, -0.4541854, -0.3725123, -0.2575871, -0.1271834, -0.004071534, 
    0.07966864, 0.1294408, 0.1621556, 0.1485489, 0.1293107, 0.1218399, 
    0.1466935, 0.2110326, 0.2445776, 0.3054336, 0.3728329, 0.4410132, 
    0.4814265, 0.523972, 0.5497372, 0.562937, 0.5337214, 0.5137833, 
    0.4460588, 0.3586891, 0.2543108, 0.1393206, 0.03370523, -0.06694579, 
    -0.1598494, -0.2401066,
  0.1121716, 0.01436877, -0.1123075, -0.2158062, -0.2894716, -0.3383811, 
    -0.3854027, -0.4333194, -0.4810407, -0.5143254, -0.5240583, -0.5104353, 
    -0.482343, -0.4418808, -0.4069036, -0.3841659, -0.3834499, -0.4253606, 
    -0.5012069, -0.6025251, -0.7049994, -0.7896185, -0.8300641, -0.8317406, 
    -0.7840683, -0.6961613, -0.57427, -0.4345891, -0.3045923, -0.2027205, 
    -0.1452336, -0.112177, -0.08161056, -0.03755128, 0.01362085, 0.05914474, 
    0.08193064, 0.06583333, 0.01389694, -0.03532171, -0.0622263, -0.07269144, 
    -0.02542639, 0.03243518, 0.0932107, 0.1288712, 0.02509534, -0.007017493, 
    -0.06990814, -0.1697291, -0.2838567, -0.39997, -0.4786159, -0.5047552, 
    -0.5030299, -0.4983912, -0.4819034, -0.4888533, -0.4683944, -0.4399924, 
    -0.4058943, -0.4728701, -0.5220075, -0.6344423, -0.7437034, -0.8023791, 
    -0.8373725, -0.8146517, -0.7686069, -0.682832, -0.5423861, -0.4110544, 
    -0.3098981, -0.1905458, -0.1162297, -0.04725182, 0.02245843, 0.1253881, 
    0.1682755, 0.2336889, 0.3725235, 0.3922338, 0.4136856, 0.4300593, 
    0.4572891, 0.4897436, 0.4940894, 0.4799129, 0.4399227, 0.3947242, 
    0.3297176, 0.3284318, 0.306036, 0.2945936, 0.2721, 0.213197,
  0.0721159, 0.06484079, 0.05911207, 0.06492233, -0.007261753, -0.03862572, 
    -0.1360378, -0.1987662, -0.3023138, -0.3397498, -0.3912635, -0.393363, 
    -0.3621292, -0.3163927, -0.2427268, -0.1736841, -0.1228053, -0.0966171, 
    -0.1000025, -0.1253767, -0.3011746, -0.4790392, -0.6869831, -0.8583531, 
    -0.9637558, -1.001386, -0.9692249, -0.8651721, -0.7557802, -0.6827822, 
    -0.6264834, -0.5660342, -0.5044293, -0.4316593, -0.3514671, -0.2790715, 
    -0.2299505, -0.2237493, -0.2464055, -0.2851751, -0.3135279, -0.3069198, 
    -0.2428899, -0.1333845, 0.01396227, 0.1304986, 0.1977677, 0.2847793, 
    0.3364232, 0.2795058, 0.1720352, 0.06122798, -0.01798752, -0.101386, 
    -0.1634953, -0.2196314, -0.2916366, -0.3955104, -0.4497422, -0.4649277, 
    -0.4677922, -0.4626164, -0.4340519, -0.3694196, -0.2757835, -0.1949731, 
    -0.1337914, -0.06486249, 0.03756261, 0.08077562, 0.00776124, 0.0753231, 
    0.118064, 0.1669084, 0.1963028, 0.2659481, 0.1778294, 0.2658828, 
    0.2838517, 0.3015763, 0.3001928, 0.3697566, 0.4362117, 0.5137833, 
    0.5704241, 0.5946917, 0.5620255, 0.4905575, 0.4757462, 0.452976, 
    0.3835912, 0.2123837, 0.150779, 0.06119514, 0.01038146, 0.06095052,
  0.3094373, 0.4054823, 0.1448219, 0.210007, 0.2379529, 0.2894015, 0.2951963, 
    0.2125628, 0.204555, 0.1335266, -0.042027, -0.145153, -0.149466, 
    -0.06048489, 0.01277399, 0.01887727, -0.02938056, -0.1103377, -0.1507511, 
    -0.1091821, -0.1724958, -0.1296744, 0.0009903908, -0.0007033348, 
    -0.08950567, -0.180326, -0.2401242, -0.3044629, -0.3831744, -0.4882193, 
    -0.5760126, -0.6092973, -0.5456905, -0.4271021, -0.2649765, -0.1452181, 
    -0.06243825, 0.004765987, 0.03101993, 0.03316832, 0.0368948, 0.02288198, 
    0.03614652, 0.0200659, 0.06671298, 0.1405411, 0.2062475, 0.3062963, 
    0.3484838, 0.3313614, 0.2593724, 0.1897598, 0.1282201, 0.09822339, 
    0.06552482, 0.03129625, 0.02358139, 0.05738688, 0.1166154, 0.1699357, 
    0.2058244, 0.1961727, 0.1954241, 0.2046362, 0.2612119, 0.3496883, 
    0.4515276, 0.5562965, 0.6261694, 0.686814, 0.7523577, 0.7586074, 
    0.7083308, 0.6321101, 0.563002, 0.5397599, 0.6030248, 0.6967748, 
    0.6306453, 0.7508601, 0.696905, 0.6823217, 0.682338, 0.7525854, 
    0.8321427, 0.8756486, 0.8435196, 0.7664526, 0.7244442, 0.7202125, 
    0.707338, 0.6868953, 0.6210915, 0.5110002, 0.3710427, 0.2923474,
  1.171547, 1.190248, 1.253969, 1.3006, 1.32005, 1.35571, 1.438393, 1.513572, 
    1.548809, 1.469464, 1.304018, 1.092836, 0.859275, 0.6813779, 0.6879201, 
    0.7731743, 0.804945, 0.6499976, 0.4506485, 0.3322891, 0.3816218, 
    0.5202286, 0.7055967, 0.8234515, 0.8471003, 0.8143206, 0.7556617, 
    0.6840307, 0.6026995, 0.4755023, 0.3609025, 0.2502744, 0.1478167, 
    0.01396203, 0.0554502, 0.1041317, 0.2120744, 0.3147762, 0.4281714, 
    0.5023903, 0.4775202, 0.4243464, 0.3280736, 0.2887833, 0.3626277, 
    0.5018041, 0.64378, 0.7530574, 0.8691056, 0.8645971, 0.7992001, 
    0.7727516, 0.7336076, 0.7595841, 0.6551245, 0.6209124, 0.5511695, 
    0.5264624, 0.5471169, 0.5901018, 0.626788, 0.6312802, 0.6116025, 
    0.5876117, 0.6365049, 0.7073219, 0.8790829, 0.9837542, 0.9976702, 
    1.038084, 1.011033, 1.00895, 1.054913, 1.132192, 1.057175, 0.924656, 
    0.9146623, 1.040688, 1.263718, 1.320326, 1.336244, 1.298565, 1.331785, 
    1.4506, 1.564402, 1.632794, 1.616762, 1.542527, 1.421742, 1.329538, 
    1.271124, 1.265736, 1.284975, 1.277064, 1.225941, 1.179701,
  1.468113, 1.490199, 1.553236, 1.592364, 1.619203, 1.671189, 1.757761, 
    1.882908, 2.051755, 2.223874, 2.366323, 2.390899, 2.197133, 1.946368, 
    1.789418, 1.805336, 1.849347, 1.879864, 1.76061, 1.576918, 1.499444, 
    1.547719, 1.647621, 1.788393, 1.881768, 1.936505, 1.966062, 1.992836, 
    2.019138, 1.982777, 2.010854, 2.051104, 2.039386, 1.910414, 1.766501, 
    1.571287, 1.445001, 1.362742, 1.377178, 1.50003, 1.5749, 1.625242, 
    1.631443, 1.667739, 1.693259, 1.784975, 1.916436, 2.008234, 2.113604, 
    2.204408, 2.229701, 2.200257, 2.134307, 2.049167, 2.028269, 1.953464, 
    1.813815, 1.693764, 1.516111, 1.393845, 1.406426, 1.39443, 1.344366, 
    1.329913, 1.236244, 1.213979, 1.323191, 1.389873, 1.443519, 1.472556, 
    1.562269, 1.649866, 1.76082, 1.927341, 2.05807, 2.092283, 2.064271, 
    2.108949, 2.26712, 2.465411, 2.596482, 2.628693, 2.755337, 2.751023, 
    2.624525, 2.40353, 2.235675, 2.180223, 2.064435, 1.909128, 1.749054, 
    1.650877, 1.67389, 1.700421, 1.645034, 1.540606,
  1.950404, 1.806101, 1.777423, 1.838978, 2.048126, 2.179962, 2.434682, 
    2.84251, 3.097035, 3.336862, 3.526755, 3.804587, 3.989173, 4.133639, 
    4.139743, 4.184909, 4.212741, 4.198581, 4.108525, 3.948874, 3.919951, 
    3.8561, 3.753415, 3.628675, 3.460609, 3.312627, 3.033802, 2.839694, 
    2.719414, 2.656653, 2.40343, 2.315475, 2.338522, 2.419626, 2.485413, 
    2.566728, 2.637252, 2.609778, 2.492917, 2.501689, 2.69513, 2.940394, 
    3.055481, 3.049622, 3.036845, 3.054179, 3.019756, 2.919853, 2.835169, 
    2.849557, 2.975892, 3.154114, 3.280319, 3.301283, 3.21585, 3.094561, 
    2.941387, 2.819349, 2.800469, 2.789694, 2.740572, 2.628073, 2.403007, 
    2.18403, 2.03556, 1.966956, 1.922344, 1.86476, 1.835203, 1.865069, 
    1.936065, 1.981833, 1.982468, 2.024883, 2.262253, 2.548484, 2.618877, 
    2.487123, 2.41406, 2.502553, 2.547263, 2.467639, 2.285836, 2.219967, 
    2.291174, 2.388978, 2.530953, 2.821741, 3.111715, 3.059437, 2.968454, 
    2.800941, 2.542951, 2.302863, 2.155206, 2.095571,
  2.018032, 1.764809, 1.54282, 1.523761, 1.470782, 1.476885, 1.597816, 
    1.822198, 2.090573, 2.327114, 2.551706, 2.798777, 3.052521, 3.335805, 
    3.585804, 3.730025, 3.806507, 3.796238, 3.597084, 3.276821, 3.087237, 
    3.013052, 2.856102, 2.726316, 2.664548, 2.597816, 2.5131, 2.430027, 
    2.367494, 2.313247, 2.276544, 2.23945, 2.190655, 2.119985, 2.114793, 
    2.289581, 2.616062, 2.894008, 2.961912, 2.961879, 2.997784, 3.068585, 
    3.181036, 3.272963, 3.323174, 3.402162, 3.459259, 3.384926, 3.236065, 
    3.125355, 3.19015, 3.378611, 3.547637, 3.694789, 3.740655, 3.715753, 
    3.625844, 3.536163, 3.476837, 3.35436, 3.1874, 3.07293, 2.959551, 
    2.809079, 2.676723, 2.606345, 2.579864, 2.513247, 2.347589, 2.12918, 
    1.967902, 1.899606, 1.831541, 1.693178, 1.61909, 1.617624, 1.546579, 
    1.426137, 1.41336, 1.543747, 1.858152, 1.993975, 1.998923, 1.941566, 
    1.87389, 1.873191, 1.977993, 2.11336, 2.163165, 2.181313, 2.161375, 
    2.152944, 2.133412, 2.127911, 2.229571, 2.189304,
  1.615509, 1.639466, 1.637936, 1.611976, 1.56108, 1.517282, 1.525387, 
    1.520065, 1.472898, 1.463344, 1.593015, 1.756866, 1.878692, 2.000535, 
    2.120489, 2.232094, 2.412075, 2.589694, 2.518243, 2.27516, 2.134894, 
    2.053025, 1.934226, 1.8909, 1.960317, 1.984616, 1.999102, 1.990541, 
    2.000014, 2.074395, 2.128904, 2.068536, 1.937986, 1.850567, 1.77726, 
    1.715964, 1.774574, 1.925892, 2.039792, 2.113555, 2.204066, 2.332012, 
    2.495195, 2.655286, 2.72026, 2.662138, 2.628708, 2.675616, 2.681313, 
    2.703138, 2.718927, 2.731671, 2.798012, 2.98377, 3.161276, 3.203171, 
    3.158005, 3.139385, 3.102992, 3.009844, 2.913148, 2.851398, 2.810007, 
    2.752325, 2.665411, 2.558527, 2.41712, 2.286798, 2.214239, 2.075469, 
    1.819968, 1.570601, 1.378936, 1.165883, 0.8866501, 0.5878067, 0.3248496, 
    0.3261695, 0.4602184, 0.6383924, 0.6527319, 0.6447401, 0.792933, 
    0.9690404, 0.9887996, 0.9724422, 1.065573, 1.217462, 1.3082, 1.371954, 
    1.457762, 1.50353, 1.462969, 1.434974, 1.470016, 1.540329,
  1.385478, 1.404506, 1.333981, 1.184194, 1.046482, 0.9118471, 0.8186655, 
    0.749135, 0.6862764, 0.6107712, 0.4643841, 0.2814569, 0.180253, 
    0.2112923, 0.3272419, 0.4408979, 0.5633926, 0.7554817, 0.9059057, 
    0.9801579, 1.113701, 1.193242, 1.070212, 0.938343, 0.939043, 0.9811821, 
    1.115345, 1.322002, 1.430336, 1.439158, 1.398402, 1.310658, 1.231378, 
    1.192835, 1.14347, 1.081849, 1.03001, 1.029523, 1.084519, 1.189337, 
    1.312578, 1.35317, 1.386617, 1.50221, 1.608249, 1.544935, 1.445896, 
    1.415167, 1.4027, 1.439744, 1.458624, 1.43307, 1.490232, 1.64059, 
    1.807729, 1.980873, 2.067689, 2.099119, 2.141518, 2.157761, 2.174281, 
    2.16546, 2.06528, 1.930108, 1.867104, 1.828904, 1.678595, 1.434096, 
    1.276267, 1.152732, 1.013539, 0.8984022, 0.7152805, 0.4611793, 0.2300596, 
    -0.06126642, -0.2888045, -0.4080606, -0.5496607, -0.8380241, -0.7993689, 
    -0.5575218, -0.4067078, -0.2966328, -0.1236849, -0.03058529, -0.07851791, 
    -0.01544857, 0.1889133, 0.4158835, 0.6671038, 0.8947568, 1.029733, 
    1.158721, 1.27944, 1.345407,
  0.4594049, 0.3989229, 0.2945938, 0.1581688, 0.0555315, -0.01439095, 
    -0.1343937, -0.3782744, -0.5882835, -0.6222029, -0.5550809, -0.4993834, 
    -0.4897156, -0.4836612, -0.4100285, -0.33708, -0.3463078, -0.3390331, 
    -0.2225618, -0.1131716, -0.009037018, 0.08023739, 0.007874489, 
    -0.07067299, -0.009620667, 0.09236336, 0.1909313, 0.2728643, 0.3536596, 
    0.4336882, 0.4166145, 0.3610153, 0.2997856, 0.1770325, 0.1266737, 
    0.1767073, 0.07800865, -0.1352396, -0.1954775, -0.214179, -0.2542667, 
    -0.222301, -0.1975298, -0.1369667, 0.01005602, 0.1057744, 0.1885056, 
    0.2350717, 0.2389774, 0.3766088, 0.5228491, 0.5209446, 0.5189099, 
    0.5449843, 0.6497045, 0.8613906, 0.9910617, 1.006524, 0.9661589, 
    0.920423, 0.9937625, 1.122783, 1.10955, 0.9861455, 0.7719526, 0.5456347, 
    0.3809209, 0.321692, 0.3238578, 0.2232885, 0.1109509, 0.1218238, 
    0.01500368, -0.2159042, -0.4535356, -0.7390499, -0.8331742, -0.9664903, 
    -1.383661, -1.671634, -1.410907, -0.9981971, -0.8785353, -0.9813514, 
    -0.933825, -0.843493, -0.8909216, -0.7826204, -0.5477405, -0.4260607, 
    -0.3016295, -0.1093121, 0.07935905, 0.284812, 0.4425917, 0.4895325,
  -0.572968, -0.6277542, -0.6600618, -0.7685585, -0.9734902, -1.121602, 
    -1.143786, -1.197073, -1.389163, -1.53275, -1.451337, -1.34232, 
    -1.289798, -1.245479, -1.222237, -1.180993, -1.168623, -1.191182, 
    -1.1363, -1.046112, -0.9615097, -0.8590517, -0.7901063, -0.7785845, 
    -0.7701516, -0.7355986, -0.7523127, -0.7559919, -0.6922069, -0.6304874, 
    -0.6070671, -0.6192255, -0.5959344, -0.6163611, -0.6780305, -0.6553411, 
    -0.7429876, -0.9318218, -1.022219, -1.111233, -1.373896, -1.331497, 
    -1.277232, -1.297382, -1.143085, -0.9788284, -0.7965045, -0.6566267, 
    -0.7860212, -0.7701373, -0.6581578, -0.6679072, -0.5902381, -0.4992385, 
    -0.4689651, -0.3951845, -0.3086939, -0.2239943, -0.1570663, -0.1611032, 
    -0.05099535, 0.01213932, 0.0259738, 0.08722067, 0.0529108, -0.08491468, 
    -0.2284365, -0.3579779, -0.3523135, -0.3732944, -0.5076361, -0.6159368, 
    -0.7920122, -0.8383813, -0.9759789, -1.255033, -1.101078, -1.18625, 
    -1.677639, -1.498505, -1.094273, -1.256806, -1.429447, -1.656416, 
    -1.802542, -1.629121, -1.501484, -1.369957, -1.151289, -0.9897819, 
    -0.801322, -0.6764035, -0.599678, -0.5377803, -0.5225129, -0.5344596,
  -1.169827, -1.205618, -1.244469, -1.394144, -1.629756, -1.982034, 
    -2.244224, -2.094566, -1.822415, -1.843297, -1.794795, -1.782946, 
    -1.916328, -1.981872, -1.998587, -1.970186, -1.861185, -1.775768, 
    -1.689846, -1.619599, -1.552835, -1.516897, -1.459378, -1.434817, 
    -1.485631, -1.424286, -1.387454, -1.318835, -1.221601, -1.335469, 
    -1.434589, -1.305748, -1.196943, -1.061347, -1.096047, -1.266506, 
    -1.121178, -0.9340682, -0.8902693, -1.002118, -1.221601, -1.251614, 
    -1.268932, -1.504186, -1.585876, -1.667712, -1.70609, -1.636348, 
    -1.692533, -1.709622, -1.613496, -1.598099, -1.577803, -1.502494, 
    -1.481009, -1.426794, -1.341637, -1.266003, -1.160745, -1.086266, 
    -1.038008, -1.027119, -1.032507, -0.9056025, -0.8551629, -0.8034534, 
    -0.7424343, -0.819469, -0.8723011, -0.98542, -1.099043, -1.213105, 
    -1.379821, -1.255781, -1.192532, -0.9883813, -0.1987656, -0.1010115, 
    -1.140367, -1.044729, -0.6633488, -1.034963, -1.052021, -1.249531, 
    -1.528225, -1.251321, -1.124254, -1.090612, -1.024189, -1.021683, 
    -1.006172, -1.093932, -1.145689, -1.200263, -1.220266, -1.14704,
  -1.10456, -1.110256, -1.137405, -1.108971, -0.7731797, -0.5717961, 
    -0.7484888, -0.8524928, -0.9019881, -1.292939, -1.618834, -1.73843, 
    -1.949351, -1.977883, -1.897691, -1.873977, -1.844208, -1.874661, 
    -1.909638, -1.917223, -1.825344, -1.809687, -1.777476, -1.677412, 
    -1.699547, -1.619045, -1.571552, -1.622382, -1.482831, -1.34538, 
    -1.083368, -0.8028183, -0.7835474, -0.7015324, -0.649677, -0.7127141, 
    -0.5847518, -0.5707545, -0.7069198, -0.8245956, -1.086282, -1.159377, 
    -1.244892, -1.524889, -1.804446, -2.097447, -2.292255, -2.33887, 
    -2.353225, -2.348293, -2.263788, -2.110029, -2.0279, -1.986575, 
    -1.960973, -1.915953, -1.845315, -1.869648, -1.828909, -1.700702, 
    -1.565286, -1.543167, -1.641116, -1.557164, -1.455569, -1.478713, 
    -1.470868, -1.41426, -1.343769, -1.397968, -1.408987, -1.437226, 
    -1.522903, -1.372773, -1.13065, -0.6545436, 0.135349, 0.3736794, 
    -0.3844914, -0.5077171, -0.308694, -0.4677595, -0.4256859, -0.4777856, 
    -0.733417, -0.6562361, -0.7388533, -0.8050806, -0.8391788, -0.9486514, 
    -1.08301, -1.309964, -1.400882, -1.433906, -1.35845, -1.152916,
  -0.7218937, -0.6246284, -0.5367539, -0.2716019, 0.1318336, 0.1771785, 
    0.07514393, -0.1321477, -0.3955753, -0.6047873, -0.9345727, -1.077151, 
    -1.255407, -1.375084, -1.214488, -1.259117, -1.37912, -1.476174, 
    -1.476321, -1.445234, -1.396568, -1.433857, -1.526272, -1.367011, 
    -1.322512, -1.24398, -1.096861, -1.046291, -0.9840845, -0.8387229, 
    -0.4886094, -0.3145207, -0.4378116, -0.5990419, -0.6432153, -0.5315455, 
    -0.3640325, -0.4980332, -0.601158, -0.540953, -0.9708518, -1.217157, 
    -1.48664, -1.777248, -1.898374, -2.008531, -2.131252, -2.214048, 
    -2.15552, -2.10954, -2.161314, -2.068671, -1.909899, -1.795592, 
    -1.724921, -1.795852, -1.793427, -1.76911, -1.817011, -1.866685, 
    -1.905748, -1.909263, -2.005797, -1.972545, -1.799091, -1.729446, 
    -1.74787, -1.76356, -1.669794, -1.580178, -1.371943, -1.247268, 
    -1.149661, -1.052737, -0.8151722, -0.3587915, -0.4201034, 0.0376929, 
    0.1071101, -0.3375187, -0.08808845, 0.1606258, 0.04373121, -0.02483976, 
    -0.4081242, -0.6148949, -0.5694684, -0.6578801, -0.8523787, -0.9322616, 
    -1.003062, -1.080162, -1.04735, -0.959052, -0.8789089, -0.7791691,
  -0.2480984, -0.12886, 0.0202117, 0.3476214, 0.4224746, 0.01939869, 
    -0.09704018, -0.1130881, -0.3529656, -0.4289579, -0.3257194, -0.1049502, 
    -0.3964872, -0.8067093, -0.6322618, -0.6411977, -0.756041, -0.8246934, 
    -0.8811064, -0.8739445, -0.8810248, -0.7962427, -0.8446798, -0.7599959, 
    -0.6674352, -0.6329613, -0.6196966, -0.5168324, -0.4607291, -0.3257511, 
    -0.077802, -0.12497, -0.265432, -0.3146355, -0.4767928, -0.342499, 
    -0.09441948, -0.3549829, -0.5341494, -0.5028182, -0.9227891, -1.062145, 
    -1.246878, -1.335143, -1.266914, -1.377185, -1.378324, -1.473392, 
    -1.513675, -1.461983, -1.535062, -1.619437, -1.572302, -1.496211, 
    -1.454642, -1.548051, -1.571358, -1.533401, -1.670266, -1.824758, 
    -2.03983, -2.063007, -1.98607, -1.903924, -1.768492, -1.609052, 
    -1.469257, -1.44613, -1.308207, -1.24683, -1.038366, -0.9361038, 
    -0.8045611, -0.6190782, -0.4437203, 0.1349261, -0.3404646, -0.005031824, 
    0.4475887, -0.4809268, -0.1804062, 0.2101374, 0.0196265, 0.1554989, 
    -0.4900577, -0.8390002, -0.5621772, -0.3165387, -0.2971702, -0.3347516, 
    -0.4420269, -0.3451688, -0.3183465, -0.3184767, -0.3226917, -0.3155308,
  -0.01224232, 0.09311199, 0.2269344, 0.5365536, 0.4185522, -0.07560456, 
    -0.07643473, -0.08084655, -0.2203643, -0.2623081, -0.1584177, 0.2315079, 
    0.199086, -0.4004915, -0.2542508, -0.07457972, -0.1170444, -0.1772823, 
    -0.4085321, -0.3818717, -0.3585162, -0.2251339, -0.2071652, -0.3007197, 
    -0.3249712, -0.17764, -0.1286006, -0.04258204, 0.03935242, 0.1089816, 
    0.2097957, 0.1956192, 0.3234349, 0.1290171, -0.1441107, -0.08745408, 
    0.02107501, -0.1299342, -0.5926619, -0.652216, -0.7316756, -0.7930212, 
    -0.6901078, -0.6367226, -0.5639358, -0.6840854, -0.6985388, -0.7997909, 
    -1.024238, -1.113479, -1.193818, -1.437681, -1.491865, -1.462096, 
    -1.391524, -1.333386, -1.410941, -1.443005, -1.554414, -1.588936, 
    -1.622334, -1.636739, -1.613822, -1.499401, -1.295772, -1.12502, 
    -1.058288, -1.114423, -0.9886909, -0.9218774, -0.7474799, -0.6077671, 
    -0.4914746, -0.1823106, -0.1268263, 0.3213353, -0.05981696, -0.02453041, 
    0.3654761, -0.1893253, -0.08050385, 0.1960587, 0.09026432, 0.3702939, 
    -0.05757046, -0.7018094, -0.3306341, -0.01318645, 0.0224576, 0.06947947, 
    -0.06725502, -0.0717802, -0.1545925, -0.1703477, -0.1275916, -0.07601261,
  0.1572404, 0.1594367, -0.002102017, 0.3286434, 0.4351375, 0.02262127, 
    0.2154597, 0.1797014, -0.1009636, -0.2754264, -0.4238153, -0.02641854, 
    0.4151667, -0.28, -0.3144894, -0.0101757, -0.0002465248, 0.1417947, 
    -0.02347231, -0.009345055, 0.09182692, 0.102211, 0.09185934, 0.1370096, 
    0.04534245, 0.1170535, 0.1940556, 0.1929164, 0.1347141, 0.2017388, 
    0.3248023, 0.5461074, 0.7235979, 0.5248184, 0.2686498, 0.1514778, 
    -0.1654329, -0.06631088, -0.2408066, -0.2339869, -0.2619176, -0.2185092, 
    -0.06906271, -0.1642451, -0.1746125, -0.3031287, -0.5047727, -0.6870642, 
    -1.026371, -1.246113, -1.263577, -1.402997, -1.436347, -1.347969, 
    -1.194925, -1.042744, -1.114245, -1.156775, -1.087276, -1.020983, 
    -0.9860387, -0.9516959, -0.946569, -0.8900089, -0.8236842, -0.7733097, 
    -0.695087, -0.5811224, -0.5371933, -0.5293808, -0.3879423, -0.2105341, 
    -0.1508985, -0.02109718, -0.07581711, 0.1690079, 0.2290176, 0.2054012, 
    0.4413386, -0.007196426, -0.07778573, 0.1228327, 0.1339656, 0.5356586, 
    0.3361788, -0.5178576, -0.2624545, 0.06461334, -0.09359074, 0.09958935, 
    0.08502293, 0.08523369, 0.09371376, 0.1207323, 0.1016726, 0.1601863,
  0.04215169, 0.1557918, -0.1151718, 0.1824683, 0.1564916, -0.1033716, 
    0.2666153, 0.2980118, 0.1800431, -0.2543163, -0.5597847, -0.3265328, 
    0.03158855, -0.2918496, -0.2735877, -0.02436876, -0.1202507, 0.1529751, 
    0.1908178, 0.1557918, 0.2645807, 0.3908663, 0.330759, 0.2677054, 
    0.1886854, 0.2442675, 0.2188277, 0.26126, 0.198678, 0.2118788, 0.3551733, 
    0.423142, 0.4698218, 0.5116026, 0.4678361, 0.3669083, 0.04215169, 
    0.2723932, 0.0234499, 0.06449938, 0.3023734, 0.08697605, 0.06602955, 
    -0.09235382, -0.1964054, -0.2863798, -0.414228, -0.5606647, -1.027868, 
    -1.344209, -1.158256, -0.9252148, -0.9332228, -0.8372917, -0.6956086, 
    -0.6078978, -0.5505242, -0.5994987, -0.5746779, -0.5901728, -0.5906124, 
    -0.5729189, -0.5672388, -0.5206404, -0.4762559, -0.3544621, -0.3045435, 
    -0.1819363, -0.2090683, -0.1334496, -0.09069252, -0.0926466, 0.001965523, 
    0.00624752, 0.05313897, 0.07138413, 0.02283278, -0.01736905, 0.07183993, 
    0.07245842, 0.03009188, 0.03696036, 0.07859451, 0.5452614, 0.4379854, 
    -0.3314323, -0.3186884, -0.001484871, 0.1175747, 0.1599083, 0.1497359, 
    0.2364874, 0.1942673, 0.1803513, 0.1422992, 0.1247368,
  0.1107397, 0.2568497, 0.05169016, 0.2742643, 0.2127419, -0.4191757, 
    -0.1569524, 0.07893631, 0.2308894, -0.1248884, -0.5647812, -0.4166861, 
    -0.5776069, -1.028747, -1.033792, -0.8652043, -0.5216341, -0.1614618, 
    0.1141238, 0.1699018, 0.07050419, 0.2662563, 0.3629684, 0.3218718, 
    0.2784958, 0.2651505, 0.2350388, 0.2406549, 0.2236457, 0.1255022, 
    0.1774714, 0.2499487, 0.04244541, 0.04919997, 0.05224356, 0.08744872, 
    0.2210915, 0.4524227, 0.06171632, -0.05666018, 0.4178038, 0.3907523, 
    0.3745415, 0.0430963, -0.3960967, -0.6007836, -0.7043478, -0.650279, 
    -0.7431185, -0.8715358, -0.788837, -0.6156116, -0.7402534, -0.6276731, 
    -0.4339228, -0.4306836, -0.3343301, -0.3853393, -0.4079299, -0.444665, 
    -0.4497094, -0.4046574, -0.3688173, -0.3081894, -0.3384628, -0.2107286, 
    -0.1366234, -0.07088566, -0.06505919, -0.05452824, -0.01030636, 
    -0.008433819, 0.03160477, -0.09598207, -0.02846931, -0.1998559, 
    -0.06650642, -0.01460212, -0.006415278, -0.03107347, -0.06484628, 
    -0.09443611, 0.03912508, 0.2299455, 0.3166471, 0.09397507, -0.2412624, 
    -0.1038775, 0.1965294, 0.06514931, 0.1609826, 0.1484013, 0.09955835, 
    0.2167773, 0.1399543, 0.1820774,
  0.1114721, 0.2078589, 0.1692035, 0.2921679, 0.5118623, -0.171324, 
    -0.06749928, 0.1223281, 0.2538875, 0.084975, -0.4422233, -0.4278841, 
    -0.4299347, -0.6506534, -0.94538, -0.9728701, -0.6236031, -0.3640494, 
    -0.09398127, 0.01651692, -0.03821945, 0.07561541, 0.2378058, 0.3410945, 
    0.31043, 0.2338834, 0.2383754, -0.03786063, 0.07984769, 0.3644832, 
    0.2444636, 0.2459122, -0.07575122, -0.1642766, 0.02605543, 0.08023834, 
    -0.05957288, 0.029392, 0.04863031, -0.02280533, 0.1259578, 0.2958798, 
    0.673728, 0.6722143, 0.4060196, 0.1322404, -0.03001547, 0.1126115, 
    0.1990373, 0.09919977, 0.0324676, 0.2025037, 0.2229786, 0.2724261, 
    0.3164687, 0.2558894, 0.1980429, 0.1841111, 0.0863409, -0.1581907, 
    -0.2550979, -0.2428908, -0.2377152, -0.2125196, -0.2593298, -0.2532263, 
    -0.1446972, -0.1523638, -0.06453705, -0.1657906, -0.1372266, -0.1758974, 
    -0.2395858, -0.187942, -0.1078802, -0.2330266, -0.1804551, 0.01596428, 
    0.000599701, -0.009719312, -0.01113532, -0.09025317, -0.1553574, 
    -0.06717384, 0.06768942, 0.3135219, -0.0734725, 0.08886385, 0.224721, 
    0.1188941, 0.2246232, 0.1339974, 0.1366014, 0.1126931, 0.05917728, 
    0.2037084,
  0.1630834, 0.1793265, 0.1521451, 0.1210099, 0.153627, 0.0289852, 
    -0.0007837564, -0.05042568, 0.05032301, 0.5183245, 0.2922335, -0.2626486, 
    0.02052188, 0.04461008, -0.1198105, -0.5229028, -0.7860215, -0.4800806, 
    -0.2610865, -0.08515871, 0.0833472, 0.07029378, 0.2821591, 0.3716611, 
    0.4196264, 0.4773738, 0.1041804, -0.1185898, 0.1108048, 0.2539362, 
    0.0166316, 0.02602288, -0.06813402, -0.1159856, -0.02353752, 0.0529272, 
    0.02061924, 0.003399186, 0.2092097, 0.4669572, 0.3012344, 0.2680964, 
    0.6475073, 1.064744, 1.301707, 1.45921, 1.730661, 1.916973, 1.583281, 
    1.354294, 1.228106, 1.081882, 0.9785943, 0.8875628, 0.7409306, 0.6180954, 
    0.504684, 0.4795537, 0.3446088, 0.2228317, 0.244072, 0.2441373, 
    0.1634245, 0.00548172, -0.01090717, -0.07217026, 0.01104879, -0.1046257, 
    -0.1090684, -0.1807802, -0.2188989, -0.3344914, -0.2986841, -0.2801782, 
    -0.2322453, -0.07026613, -0.1573267, 0.01311598, 0.02065179, 
    -0.002915919, -0.06657152, -0.3709661, -0.2507186, 0.01868248, 
    0.05136395, 0.400599, 0.3125615, 0.480515, 0.4537401, 0.3767383, 
    0.3198376, 0.3346658, 0.2889787, 0.1597632, 0.2517553, 0.2515599,
  0.1153297, -0.08903313, -0.2638693, 0.06959391, 0.0965144, 0.04591224, 
    0.007468194, 0.01847079, 0.2835587, 0.7428034, 0.6741996, 0.09501708, 
    0.1490211, 0.2555151, 0.1774063, -0.2048692, -0.4137394, -0.3022161, 
    -0.3598821, -0.2341008, -0.1515813, -0.2928247, -0.08252206, 0.06990308, 
    0.2448705, 0.5681291, -0.1103539, -0.1325383, 0.08811605, -0.3731959, 
    -0.2090032, 0.001071706, -0.0357447, -0.09365487, -0.1676131, 
    -0.07422113, 0.2996882, 0.5981258, 0.5822892, 0.5847143, 0.4775691, 
    0.4799128, 0.7128556, 0.9145971, 0.9556778, 1.073679, 1.39251, 1.400144, 
    1.194073, 1.191827, 1.316957, 1.20947, 1.1096, 1.025111, 0.9414039, 
    0.8571754, 0.7497697, 0.7300096, 0.7044568, 0.6691542, 0.6039686, 
    0.5216122, 0.4491506, 0.3853645, 0.3183236, 0.1683078, 0.1562641, 
    0.1122861, 0.0263648, -0.1056991, -0.2409693, -0.3419622, -0.244566, 
    -0.4605989, -0.3792672, -0.0948267, -0.1525904, -0.04069263, 0.09661207, 
    -0.08128506, -0.4074569, -0.1017603, -0.2616398, 0.1176562, -0.02555704, 
    0.1102991, 0.04666018, 0.1947238, 0.2178688, 0.2634904, 0.3502253, 
    0.3629532, 0.2465958, 0.190183, 0.1072242, -0.03270078,
  0.06659901, -0.05565023, 0.06604564, 0.2174454, 0.3532039, 0.2960912, 
    0.2577448, 0.2777807, 0.3053685, 0.1312638, 0.1210749, 0.2590797, 
    0.4206682, 0.5169892, 0.4701636, 0.2644831, 0.04970449, -0.2530136, 
    -0.4561871, -0.5420923, -0.6015323, -0.6821965, -0.8514347, -0.6526717, 
    -0.5618516, -0.2456568, -0.134703, -0.2009628, -0.4819195, -1.157945, 
    -0.7764837, -0.3389348, -0.2654972, -0.3244978, -0.7563502, -0.3607123, 
    0.2373021, 0.5373022, 0.4668919, 0.4038223, 0.4281876, 0.5850562, 
    0.67031, 0.5604142, 0.3680634, 0.04504871, -0.2866075, -0.4703155, 
    -0.4590359, -0.4143915, -0.3466334, -0.239814, -0.2026882, -0.3213406, 
    -0.3566601, -0.3951528, -0.4324088, -0.3994987, -0.3453484, -0.3259797, 
    -0.2071638, -0.08242416, -0.1172223, -0.1520858, -0.10552, 0.03092206, 
    0.09063888, 0.1817847, 0.1888484, 0.149379, 0.1197566, 0.06729889, 
    -0.07591397, -0.3630233, -0.1211936, 0.01489007, -0.1956403, -0.02008724, 
    0.04905348, -0.3919621, -0.2549503, -0.08773088, -0.2101436, -0.3982134, 
    -0.3376327, -0.2769394, -0.2188184, 0.07610345, 0.1036272, 0.2145647, 
    0.2422501, 0.07649487, 0.03080821, 0.1547503, 0.06791741, 0.004652441,
  0.05064854, 0.09548903, 0.1527807, 0.1806128, 0.2890925, 0.3304011, 
    0.4357399, 0.1455705, 0.04075268, 0.1431289, 0.1290827, 0.2897437, 
    0.6281878, 0.6823215, 0.6596816, 0.3069472, -0.06240463, -0.3393576, 
    -0.3907574, -0.3987654, -0.454169, -0.5987492, -0.8925164, -0.8026233, 
    -1.000328, -1.130538, -0.7946482, -0.4646021, -0.7529325, -0.9623563, 
    -0.7480005, -0.7105168, -0.1842961, -0.1910181, -0.5448919, 0.08520257, 
    0.5045711, 0.30545, 0.04369879, 0.1002254, 0.315964, 0.4946098, 
    0.5313933, 0.2688451, 0.1491022, -0.05750656, -0.2744665, -0.3106971, 
    -0.3335161, -0.4818234, -0.5049353, -0.5409055, -0.6822629, -0.9259315, 
    -0.9131546, -0.825736, -0.7465858, -0.6261101, -0.5133662, -0.4336624, 
    -0.4055853, -0.4590683, -0.5361521, -0.4340692, -0.2032092, 0.1949842, 
    0.320472, 0.5283337, 0.5633273, 0.5367482, 0.58722, 0.6196742, 0.1787734, 
    -0.3381705, -0.03688401, -0.06885016, -0.1339542, -0.2379904, -0.5453157, 
    -0.7047558, -0.5567083, -0.1770859, -0.2369003, -0.1438842, -0.007506847, 
    0.1238575, 0.3019333, 0.4486465, 0.5056937, 0.6353323, 0.6178197, 
    0.7715306, 0.7945291, 0.4609839, 0.2000788, 0.164239,
  -0.1296899, -0.2047875, -0.09167004, 0.1272764, 0.09093142, 0.01226902, 
    0.2319627, 0.009486675, 0.2916153, 0.585349, 0.1602515, -0.05887282, 
    0.1274393, 0.2970676, 0.5343881, 0.3965306, 0.1814425, 0.1862597, 
    0.138165, 0.3295875, 0.02188885, -0.4303257, -0.3200221, -0.4384136, 
    -0.5597196, -0.5009151, -0.4799504, -0.240042, -0.275393, -0.009540081, 
    0.1314754, -0.1371772, -0.105325, -0.257929, -0.2191105, 0.1534481, 
    0.3427706, 0.1345994, -0.1290073, -0.1012716, 0.0357399, 0.1150031, 
    0.2331185, 0.05377245, -0.129528, -0.2618842, -0.2034531, -0.0673852, 
    0.03736734, 0.07525778, 0.204587, 0.2011204, 0.1515436, 0.1681938, 
    0.3758936, 0.6019344, 0.6823702, 0.62918, 0.3317685, 0.09255838, 
    -0.1049023, -0.1961946, -0.1215529, 0.1237764, 0.3939257, 0.5413866, 
    0.3469374, 0.2783012, 0.2497041, 0.5957656, 0.9149873, 0.7882617, 
    0.0775857, -0.3832228, -0.08405304, -0.4993515, -0.8042836, -0.9834175, 
    -0.8138866, -0.6581898, -0.353241, -0.06147671, 0.02073193, 0.1449194, 
    0.3462543, 0.6097455, 0.7046676, 0.7647591, 0.8814917, 0.8452444, 
    0.891875, 1.214727, 0.6714005, 0.1903784, -0.1935894, -0.07400966,
  -0.3021181, -0.2930534, -0.0584507, 0.18294, 0.05154276, -0.1697454, 
    0.04501677, 0.3181779, 0.5771134, 0.5100398, 0.1372207, -0.2055202, 
    -0.1005726, 0.09784913, 0.05382252, 0.2448869, 0.3649063, 0.3533506, 
    0.210804, 0.3109019, 0.03845787, -0.2248232, -0.07825756, -0.2814322, 
    -0.0863955, 0.189841, -0.1484398, -0.2576845, -0.1859572, 0.1231091, 
    0.08682919, -0.02205753, 0.001347542, -0.1357121, -0.05247688, 0.2985482, 
    0.5791955, 0.2753386, -0.001077652, 0.1204715, 0.3814254, 0.340817, 
    0.2489061, -0.001695156, -0.1600447, -0.2092795, -0.08208275, -0.1116886, 
    -0.128356, -0.09791851, -0.01079273, 0.08539867, 0.2738419, 0.508997, 
    0.5921354, 0.5398731, 0.3233213, 0.08946705, -0.2057323, -0.3475122, 
    -0.3500023, -0.1897821, 0.01368427, 0.1671844, 0.2608862, 0.2589655, 
    0.1367652, -0.06928921, -0.1658064, 0.1005184, 0.3295548, 0.08486068, 
    -0.4219915, -0.31514, 0.1504374, -0.242321, -0.4334497, -0.3830752, 
    -0.2151718, -0.1067743, 0.08925438, 0.1602669, 0.3493295, 0.5567999, 
    0.6939907, 0.8075652, 0.8424282, 0.9355106, 0.8517218, 0.7332821, 
    0.7081027, 0.6835907, -0.09583569, -0.3899283, -0.2581902, -0.2549992,
  -0.4385602, -0.5598011, -0.6210644, -0.2936871, -0.3392274, -0.3133812, 
    -0.0396831, 0.2781878, 0.5477189, 0.5197729, 0.6310848, 0.06261158, 
    -0.273603, -0.03973222, -0.2730168, -0.2352562, 0.05136442, -0.01789045, 
    -0.06992483, -0.04137659, -0.0527041, -0.1184433, -0.2222356, 
    -0.08846283, 0.08990628, 0.08888096, -0.07760668, -0.1693547, 0.02013087, 
    0.2930964, 0.01622486, -0.1305537, -0.2860537, -0.08896828, 0.1627078, 
    0.3567357, 0.4274874, 0.08980894, -0.05316114, 0.08953094, 0.1771774, 
    0.06236601, -0.01795626, -0.17834, -0.1411328, -0.01678324, 0.1255507, 
    0.06713533, 0.0759902, 0.1553197, 0.1790004, 0.3393369, 0.472784, 
    0.5810184, 0.4925094, 0.3252249, 0.09174538, -0.1410828, -0.276907, 
    -0.2412453, -0.1997743, -0.1250525, 0.1112432, 0.2512507, 0.212399, 
    0.2087541, 0.2284968, 0.0838517, 0.00265038, 0.2654109, 0.1386695, 
    -0.13594, -0.4023787, -3.528595e-005, 0.4561496, 0.2812152, 0.3991013, 
    0.4099898, 0.3113747, 0.3008428, 0.4433732, 0.5000138, 0.5084448, 
    0.5633926, 0.6885872, 0.7340946, 0.7108035, 0.6054163, 0.4615688, 
    0.4413214, 0.4641089, 0.6075325, -0.03170848, -0.402916, -0.4224966, 
    -0.481415,
  -0.5782251, -0.87357, -1.097578, -0.8021183, -0.9384143, -0.5492699, 
    0.04441488, 0.0526017, 0.4079728, 0.3721655, 0.09208739, -0.2477405, 
    -0.3663435, -0.04809827, -0.1849472, -0.2196801, -0.1348331, -0.04575443, 
    -0.07034755, -0.1409854, -0.2412948, -0.2862004, -0.2195827, 0.03093824, 
    0.04478917, 0.05064845, -0.1051783, -0.5055853, -0.05521083, 0.20239, 
    -0.04642153, 0.009193659, -0.1213076, 0.04786444, 0.2988081, 0.1288385, 
    -0.07508469, -0.1650591, -0.1942091, -0.1838903, -0.2410846, -0.3684769, 
    -0.3561559, -0.3629103, -0.1768427, -0.05091476, -0.08315802, -0.1256218, 
    -0.006465435, 0.02786112, 0.008004189, 0.08853817, 0.01659822, 
    0.04578114, -0.07445002, -0.2791376, -0.4052119, -0.5471878, -0.6312046, 
    -0.6201043, -0.5070996, -0.288187, -0.07982063, -0.01959944, 0.04434943, 
    0.2346817, 0.4337703, 0.3032202, 0.1978654, 0.2133764, -0.09840745, 
    -0.3109401, -0.2510929, 0.04810905, 0.222312, 0.2199845, 0.4549289, 
    0.4641576, 0.4667449, 0.4460747, 0.3595512, 0.3267877, 0.3118458, 
    0.3816862, 0.3652642, 0.2780404, 0.1950822, 0.02888775, -0.2204938, 
    -0.5949092, -0.6753449, -0.2432966, -0.4917994, -0.8498564, -1.146015, 
    -1.036608,
  -0.9235054, -1.107343, -1.003957, -0.6074082, -0.6003932, -0.1202011, 
    0.08359124, -0.1223821, 0.1538223, -0.04023689, -0.4914739, -0.2767764, 
    0.02195388, 0.09166408, -0.08252206, -0.1590845, -0.03056896, 0.04736076, 
    -0.0430038, 0.02356517, 0.1361792, 0.02981532, 0.06803143, 0.01703858, 
    -0.005275846, 0.2298477, -0.04111564, -0.3108586, 0.1561816, 0.2617164, 
    -0.02168202, 0.09301543, 0.1189101, 0.1448207, 0.1648402, 0.02416658, 
    -0.2702336, -0.5528512, -0.7646022, -0.7476914, -0.6040883, -0.6046746, 
    -0.6501005, -0.6007352, -0.3831728, -0.2771838, -0.25137, -0.1343453, 
    -0.03592396, -0.008775473, 0.06210661, 0.111016, 0.06516647, 0.04324198, 
    -0.111722, -0.243525, -0.351305, -0.4880242, -0.4907088, -0.5838566, 
    -0.5746937, -0.4314487, -0.2924664, -0.09140885, 0.2193334, 0.34684, 
    0.2820288, 0.200616, 0.02371174, -0.03314054, -0.01028897, -0.0266788, 
    0.03206062, 0.06029987, -0.1446151, -0.08025932, 0.1744275, 0.08853936, 
    -0.1219425, -0.3048851, -0.347187, -0.2734072, -0.2571311, -0.2710636, 
    -0.3080268, -0.2407906, -0.2887237, -0.5319035, -0.8465035, -1.278827, 
    -1.546519, -1.698847, -1.456741, -0.8900577, -1.010061, -1.075491,
  -0.5049504, -0.4445338, -0.2560572, -0.2188827, -0.2731959, -0.2522648, 
    -0.1872583, -0.275442, -0.575865, -0.7432967, -0.4274114, 0.03059645, 
    0.05118561, -0.1744165, -0.2749862, -0.07972257, 0.01931715, -0.05599213, 
    -0.1556503, -0.02269125, -0.09676349, -0.2927759, -0.2161651, -0.360631, 
    -0.3405628, -0.3734083, -0.7588739, -0.4320826, 0.04677391, 0.190834, 
    0.2135719, 0.2426897, 0.242722, 0.3331351, 0.2027967, 0.1002095, 
    -0.1451364, -0.4162459, -0.5660179, -0.6638043, -0.7076032, -0.7368189, 
    -0.6806666, -0.5752956, -0.5025741, -0.5333033, -0.479332, -0.3613306, 
    -0.3116561, -0.2959823, -0.2254582, -0.1333358, -0.02636971, -0.05114184, 
    -0.2755233, -0.4423202, -0.6543808, -0.7986354, -0.7644883, -0.7855821, 
    -0.6757512, -0.4887233, -0.3202173, -0.07138932, 0.1340795, 0.1255509, 
    0.03741622, 0.06433666, 0.01725006, 0.01829177, 0.1130021, 0.07774806, 
    -0.09581959, -0.1835312, -0.4056177, -0.5976263, -0.5372095, -0.6047226, 
    -0.6882513, -0.6764022, -0.6568873, -0.7225448, -0.8432968, -0.9148787, 
    -0.9048202, -0.8056502, -0.843899, -0.9304387, -1.155732, -1.606415, 
    -1.999758, -2.295852, -2.099905, -1.535761, -0.9625514, -0.654983,
  -0.1133326, -0.04993725, -0.04614496, 0.2085102, 0.499835, 0.4670223, 
    0.4332331, 0.213051, -0.5067244, -0.5200709, 0.06873131, 0.08836007, 
    -0.1219264, -0.1683782, -0.02169847, 0.02947339, 0.002178475, 
    -0.07780199, -0.1802922, -0.2062851, -0.4082706, -0.2497091, -0.07088459, 
    0.02756882, -0.1940944, -0.3118029, -0.2929873, 0.2082495, 0.2384742, 
    0.1348445, 0.1438289, 0.1975886, 0.3075007, 0.4901342, 0.3148087, 
    0.2413224, 0.05575922, -0.1178899, -0.2001977, -0.2606794, -0.3220402, 
    -0.3608584, -0.3429232, -0.2903354, -0.2162304, -0.1678257, -0.10181, 
    -0.03390622, -0.04901052, -0.1210482, -0.1692085, -0.1911323, -0.2467966, 
    -0.4090683, -0.5991566, -0.7397983, -0.8243196, -0.7510939, -0.6876011, 
    -0.7236843, -0.6000512, -0.3937848, -0.1140647, 0.06384838, 0.009291109, 
    -0.0402531, 0.1098119, 0.305043, 0.3939588, 0.1916482, 0.06495512, 
    -0.04288989, -0.2243025, -0.3063665, -0.3340519, -0.4554712, -0.6778508, 
    -0.8477563, -0.8984236, -0.8510115, -0.8867537, -0.943785, -0.9554548, 
    -0.9929711, -1.079267, -1.221112, -1.260224, -1.144062, -1.273961, 
    -1.557196, -1.637812, -1.67707, -1.785224, -1.789537, -1.281318, 
    -0.3841008,
  -0.02571893, 0.03443742, 0.3461885, 0.8387673, 1.1381, 1.023826, 0.5443171, 
    0.3496557, 0.1310034, 0.2161433, 0.112058, -0.1227239, -0.07358649, 
    0.01445061, 0.1270158, 0.04234767, 0.03232172, -0.05423415, -0.1529484, 
    -0.0200057, 0.300909, 0.2103164, 0.1505509, 0.1177384, 0.2402807, 
    0.2096817, 0.3311172, 0.6373835, 0.5784155, 0.1801571, -0.00324142, 
    0.07400477, 0.06983793, 0.02520907, -0.1320176, -0.1404979, -0.1398787, 
    -0.1912787, -0.1865096, -0.04801798, -0.0004591942, -0.01808643, 
    0.09721327, 0.2795372, 0.3819461, 0.3981571, 0.3732715, 0.3882451, 
    0.4122686, 0.3770962, 0.2640104, 0.05071259, -0.2967157, -0.653584, 
    -0.8826861, -1.02349, -1.073814, -0.9987984, -0.9234891, -0.8202348, 
    -0.6586938, -0.4823275, -0.141881, 0.1333797, 0.03443754, 0.0590958, 
    0.1900202, 0.2999978, 0.3593717, 0.2876437, 0.07055426, -0.08017802, 
    -0.2194685, -0.366197, -0.4079123, -0.4069035, -0.4561384, -0.6791213, 
    -0.8329294, -0.8067091, -0.7364781, -0.6365106, -0.5765495, -0.6406934, 
    -0.7447784, -0.8633661, -0.9610548, -1.027754, -1.115416, -1.038577, 
    -0.9291208, -0.9568551, -0.8012724, -0.4212264, 0.07869215, 0.2000951,
  0.5526507, 0.7866189, 1.086977, 0.9683731, 0.7946752, 0.7529597, 0.8209448, 
    0.7386042, 0.6157364, 0.5443171, 0.2802221, 0.3006486, 0.3837052, 
    0.2856095, 0.1609839, 0.05735433, -0.04458249, -0.08592373, -0.04988858, 
    0.02299553, 0.04120833, -0.1815455, -0.2400091, 0.0451147, 0.1729467, 
    0.06472731, 0.01617551, -0.04850531, -0.08543539, -0.2048697, -0.1160026, 
    0.03280973, -0.0229845, -0.1810417, -0.1730826, -0.1335971, -0.02721739, 
    0.01646805, -0.01409769, 0.04296637, 0.08028793, 0.1700821, 0.2717581, 
    0.3451138, 0.4355278, 0.578577, 0.6699505, 0.7324352, 0.8214164, 
    0.8360977, 0.6949844, 0.4209614, 0.1042128, -0.1614609, -0.431807, 
    -0.6691279, -0.7253613, -0.6233759, -0.5493851, -0.4468136, -0.3674679, 
    -0.2388382, 0.01399517, 0.1853653, 0.2155087, 0.2311664, 0.257647, 
    0.1527319, 0.1834273, 0.0964818, -0.2185419, -0.4094267, -0.3470247, 
    -0.3108594, -0.435257, -0.4887724, -0.328486, -0.2549024, -0.3369007, 
    -0.425036, -0.3871446, -0.2045441, -0.05589533, -0.04733372, -0.1240263, 
    -0.2378278, -0.2859397, -0.3389025, -0.3721051, -0.295022, -0.1926298, 
    0.009681702, 0.3790503, 0.5846982, 0.563702, 0.5767877,
  1.201771, 0.9403783, 0.9955704, 0.9007623, 0.7691218, 1.102878, 1.380792, 
    1.091127, 0.7873836, 0.6673803, 0.5998021, 0.6475561, 0.5025365, 
    0.09776767, -0.07366788, -0.1057968, -0.1640487, -0.08937427, 
    -0.007082641, -0.07916918, -0.1062525, -0.1014022, -0.1337753, 
    -0.1177271, -0.08066659, -0.01230717, -0.05680561, -0.2087429, -0.211282, 
    -0.05195642, 0.08355808, 0.1795874, 0.1624975, 0.1466446, 0.1779752, 
    0.1121068, 0.04701805, 0.1635227, 0.132874, 0.1280737, 0.2731724, 
    0.4394169, 0.50348, 0.5269661, 0.6011515, 0.6946583, 0.7513304, 
    0.7930632, 0.80509, 0.7474413, 0.6360321, 0.5107718, 0.3594213, 
    0.1780567, -0.03455639, -0.1548862, -0.09695864, 0.00530386, 0.001135826, 
    -0.04446936, -0.0174675, 0.06471014, 0.2620578, 0.3893529, 0.3502743, 
    0.2380674, 0.1476212, 0.2206345, 0.3131638, 0.1257625, -0.04601526, 
    -0.05809188, -0.03854465, 0.01342511, -0.1508976, -0.274921, -0.2515486, 
    -0.186542, -0.2231958, -0.1928086, -0.02042866, 0.085886, 0.088099, 
    0.07820415, 0.03666639, -0.08548546, -0.1495156, -0.106514, -0.0494504, 
    0.06173134, 0.3305793, 0.8063931, 1.220065, 1.356573, 1.50501, 1.496205,
  1.474054, 1.483998, 1.802732, 1.729929, 1.550909, 1.71821, 1.694676, 
    1.242136, 0.9073706, 0.8301569, 0.6661108, 0.4580704, 0.23906, 
    -0.03699794, -0.2084009, -0.2175155, -0.1827662, -0.227151, -0.3593125, 
    -0.4376328, -0.3771996, -0.3041855, -0.3035995, -0.350507, -0.2852085, 
    -0.2000034, -0.1765819, -0.2384791, -0.1507516, 0.07504606, -0.04979157, 
    0.09791422, 0.1196423, 0.1106575, 0.2111464, 0.2468238, 0.2786431, 
    0.07553434, -0.1182151, 0.06223679, 0.3703914, 0.6004686, 0.7455368, 
    0.929863, 1.072799, 1.051999, 1.059127, 1.17301, 1.168421, 0.9637499, 
    0.7756801, 0.6670208, 0.5409145, 0.3670864, 0.2456999, 0.2140589, 
    0.2535286, 0.2842412, 0.3641567, 0.5385542, 0.6921353, 0.6650529, 
    0.5143367, 0.5314265, 0.6435523, 0.4943979, 0.3723111, 0.4313602, 
    0.4386044, 0.2863896, 0.173907, 0.1008766, -0.004396915, -0.07186115, 
    -0.06870365, -0.1210474, -0.181806, -0.1013858, 0.06352293, 0.1239558, 
    0.1906059, 0.01998472, 0.06664777, 0.1423802, 0.1416306, 0.02830124, 
    -0.1010766, -0.1201196, -0.006382465, 0.1823368, 0.4947066, 0.8941374, 
    1.185463, 1.433705, 1.706426, 1.759795,
  2.115362, 2.49308, 2.253025, 1.852146, 1.706231, 1.831605, 1.744594, 
    1.253513, 0.8615537, 0.7067521, 0.5229306, 0.3088516, 0.167071, 
    0.04734445, -0.1170273, -0.2027205, -0.2407413, -0.2721052, -0.3175652, 
    -0.3515332, -0.3984733, -0.4606955, -0.3789899, -0.1506705, 0.08725238, 
    0.01046228, 0.1031218, 0.1033659, 0.04205394, 0.1258759, 0.09809256, 
    0.1811333, 0.2699838, 0.3612444, 0.4046679, 0.4412241, 0.2779589, 
    -0.2314324, -0.2555037, 0.2362924, 0.7591116, 0.9263648, 0.8686012, 
    1.158038, 1.480857, 1.666746, 1.658477, 1.522002, 1.348158, 1.130743, 
    0.9287736, 0.7091286, 0.4349263, 0.2668266, 0.301446, 0.4652319, 
    0.7037396, 0.9074683, 1.104083, 1.211993, 1.070001, 0.7405249, 0.5136694, 
    0.6243627, 0.7311013, 0.5785449, 0.4291806, 0.4682915, 0.4581032, 
    0.3401181, 0.2422989, 0.2479794, 0.218536, 0.1786435, 0.2812641, 
    0.4637673, 0.5830219, 0.4601864, 0.4004533, 0.3385556, 0.309063, 
    0.2321582, 0.4689746, 0.6167781, 0.5695605, 0.3834767, 0.2302709, 
    0.1913548, 0.273663, 0.4502902, 0.7905574, 1.240313, 1.658314, 1.841062, 
    1.828709, 1.942234,
  1.996938, 1.917103, 1.577878, 1.127618, 1.097231, 1.320114, 1.188067, 
    0.7498346, 0.387351, 0.2685847, 0.204457, 0.08813226, -0.01237226, 
    -0.08138275, -0.06982684, 0.002536654, 0.06171632, 0.163718, 0.2234998, 
    0.2793593, 0.284893, 0.2464974, 0.2991829, 0.4105768, 0.4147592, 
    0.2814267, 0.2056291, 0.2017715, 0.2444313, 0.1471493, 0.1956353, 
    0.3251429, 0.376039, 0.4274871, 0.4373991, 0.3679981, 0.1327286, 
    0.07255507, 0.2408664, 0.7689591, 1.095603, 1.056735, 0.7033179, 
    0.7392392, 1.076934, 1.262888, 1.299493, 1.25475, 1.247312, 1.259959, 
    1.15169, 0.8609024, 0.5335424, 0.3616511, 0.3951147, 0.5601537, 
    0.7387019, 0.9088842, 1.04238, 1.046889, 0.876609, 0.6196589, 0.6224421, 
    0.5373348, 0.3651017, 0.3042618, 0.4771135, 0.648142, 0.5568334, 
    0.3396621, 0.2372208, 0.3802224, 0.639353, 0.9358375, 1.161228, 1.251707, 
    1.018357, 0.5601377, 0.2028623, 0.112643, 0.1424608, 0.5393198, 
    0.7643368, 0.7396624, 0.627553, 0.524395, 0.5418596, 0.6917622, 
    0.9005511, 1.075209, 1.250681, 1.480955, 1.738849, 1.90353, 1.935072, 
    1.891095,
  0.3115535, 0.2577123, 0.2276668, 0.3053685, 0.3420873, 0.194659, 
    0.07971752, -0.05662689, -0.1444198, -0.1320501, -0.1906112, -0.2985865, 
    -0.3479517, -0.3172877, -0.2290716, -0.08584237, 0.02573001, 0.1209773, 
    0.1983702, 0.3233376, 0.4807105, 0.4619118, 0.3844702, 0.338474, 
    0.2520646, 0.2336238, 0.2987932, 0.3431128, 0.3397763, 0.2505186, 
    0.4255178, 0.4932427, 0.4963186, 0.4278779, 0.336977, 0.1813617, 
    0.07760179, 0.1402644, 0.2262995, 0.3933733, 0.3123186, 0.3701475, 
    0.3542293, 0.3303523, 0.3520973, 0.4799619, 0.6234834, 1.050436, 
    1.104457, 0.8696098, 0.4325495, 0.02856207, -0.2245629, -0.2542502, 
    -0.1714377, -0.01209545, 0.07314229, 0.2129695, 0.2982397, 0.2966936, 
    0.2834772, 0.2591772, 0.2932754, 0.2114234, 0.1682266, 0.3198217, 
    0.5619768, 0.5597143, 0.5033665, 0.4225072, 0.5301896, 0.8088679, 
    1.090378, 1.173874, 1.099167, 0.9622534, 0.6567032, 0.2954076, 
    0.03370512, -0.02718341, 0.06570399, 0.153985, 0.06931716, -0.137763, 
    -0.1427597, -0.1956568, -0.08312428, 0.1447729, 0.3889949, 0.6597306, 
    0.8143692, 0.8899063, 0.982875, 1.027813, 0.8721655, 0.5629206,
  -0.7625188, -0.7033228, -0.4987655, -0.3169459, -0.2857609, -0.4348495, 
    -0.5003931, -0.4735864, -0.4756047, -0.5776067, -0.7554062, -0.799205, 
    -0.6982936, -0.5017929, -0.3631047, -0.2538437, -0.1862655, -0.07959223, 
    0.1102355, 0.2986467, 0.4710426, 0.4757789, 0.3966446, 0.3293106, 
    0.3447402, 0.4096004, 0.5344703, 0.5579728, 0.5666313, 0.6461728, 
    0.5267061, 0.4221818, 0.3957496, 0.2775691, 0.1240209, 0.1019994, 
    0.264353, 0.2966935, 0.3051245, 0.2249324, 0.1534805, 0.1850723, 
    0.2519343, 0.2884089, 0.2900041, 0.3040178, 0.3789039, 0.3928199, 
    0.1975563, -0.1868187, -0.5714705, -0.6644716, -0.5373561, -0.3008168, 
    -0.175719, -0.0938499, -0.04188061, 0.1235163, 0.2957169, 0.3660131, 
    0.2675593, 0.1008276, 0.04242912, 0.1463517, 0.3705216, 0.5301245, 
    0.6346818, 0.642185, 0.6057429, 0.5516577, 0.4785782, 0.3700171, 
    0.1386694, -0.02068935, -0.2405136, -0.2947129, -0.2651718, -0.09977466, 
    -0.1476099, -0.211412, -0.3157903, -0.2632837, -0.2280464, -0.09694338, 
    -0.104804, -0.02653337, -0.02962518, 0.1466763, 0.391485, 0.6661429, 
    0.8215954, 0.7531227, 0.6385554, 0.3211238, -0.1077662, -0.5350448,
  -0.6989281, -0.7809921, -0.8587102, -0.9540716, -1.040367, -0.9779485, 
    -0.9115422, -0.8511255, -0.913886, -1.010029, -1.09595, -1.326516, 
    -1.105032, -0.7929225, -0.4473495, -0.3082056, -0.1796086, -0.04847252, 
    0.03476357, 0.1573383, 0.2706031, 0.3598119, 0.4123511, 0.4683081, 
    0.5475398, 0.6212378, 0.648517, 0.5807593, 0.4571917, 0.2829893, 
    0.1519182, 0.1461239, 0.229506, 0.2684219, 0.3493789, 0.3758926, 
    0.4476538, 0.3733699, 0.4380672, 0.4554664, 0.4758441, 0.3867489, 
    0.3888809, 0.2923965, 0.1982397, 0.1567195, 0.004099041, -0.3761906, 
    -0.8525578, -1.233873, -1.608189, -1.652118, -1.425523, -0.4245954, 
    -0.0802443, 0.004310846, 0.0887183, 0.1669083, 0.2174616, 0.09273833, 
    0.01879627, -0.009963393, 0.01700604, 0.2006159, 0.3261044, 0.4788874, 
    0.5906225, 0.568308, 0.4538875, 0.2225398, 0.008867919, -0.1471868, 
    -0.2157903, -0.450328, -0.2227402, -0.1249212, -0.1869329, -0.2008488, 
    -0.4431829, -0.6521022, -0.7286972, -0.6045601, -0.2681344, -0.1865258, 
    -0.2140489, -0.2974467, -0.3032578, -0.2125351, -0.05232999, 0.156752, 
    0.3416966, 0.3665503, 0.2336076, -0.05026305, -0.3321639, -0.5634302,
  -0.7208846, -0.7289738, -0.7611353, -0.8020694, -0.8096053, -0.7912947, 
    -0.7630883, -0.7490097, -0.7832546, -0.8261256, -0.8012557, -0.676744, 
    -0.4331243, -0.1890162, -0.03690034, 0.03186597, 0.2948543, 0.3174779, 
    0.2188452, 0.04143628, 0.05886793, 0.1549617, 0.238116, 0.3503556, 
    0.4544734, 0.5075336, 0.4756813, 0.3575823, 0.2570615, 0.2159318, 
    0.2253394, 0.3705217, 0.545831, 0.6414526, 0.6093888, 0.5188453, 
    0.3738908, 0.2369115, 0.1590795, 0.1690567, 0.1328588, 0.1630183, 
    0.1089981, 0.02418369, -0.03976488, -0.05024664, -0.07466072, -0.1661809, 
    -0.3457057, -0.5683618, -0.7586287, -0.8018744, -0.7071159, -0.5409043, 
    -0.4448273, -0.4113472, -0.4549019, -0.5670927, -0.6571641, -0.6715033, 
    -0.5809109, -0.3514514, -0.06723928, 0.03879976, 0.1904111, 0.263523, 
    0.2331356, 0.1138321, -0.0518254, -0.3694361, -0.4057643, -0.4533553, 
    -0.5725774, -0.446015, -0.3966172, -0.3908066, -0.4229355, -0.715302, 
    -0.7744655, -1.002688, -1.088089, -0.455374, -0.2609246, -0.22528, 
    -0.3061222, -0.4444035, -0.7011914, -0.8565626, -0.7361355, -0.6096714, 
    -0.4784203, -0.414065, -0.6408716, -0.7712265, -0.800979, -0.7394553,
  -0.9266463, -0.6913596, -0.5131049, -0.3276885, -0.1663277, -0.1610541, 
    -0.2722039, -0.5588076, -0.7587106, -0.8356799, -0.9286976, -0.8923364, 
    -0.8190942, -0.6443222, -0.486184, -0.452037, -0.4358585, -0.4144232, 
    -0.3405624, -0.2578313, -0.1239772, 0.01804757, 0.1471003, 0.3024226, 
    0.3816219, 0.2769018, 0.2696427, 0.1927384, 0.1301895, 0.104864, 
    0.2199356, 0.3007137, 0.3645971, 0.368715, 0.2976375, 0.1440893, 
    0.02892002, -0.01784116, -0.006708264, -0.00714761, 0.00481528, 
    0.01251382, -0.01356053, -0.07609308, -0.1433619, -0.1841985, -0.1890975, 
    -0.1676133, -0.1429062, -0.1314477, -0.1633162, -0.2025089, -0.2353537, 
    -0.2593122, -0.2717471, -0.2665875, -0.2494977, -0.2288435, -0.1842144, 
    -0.1350285, -0.07996666, -0.02550697, 0.01036537, 0.0561173, 0.03494215, 
    -0.2452661, -0.370429, -0.4883488, -0.5857121, -0.652916, -0.6837429, 
    -0.6272324, -0.6042506, -0.5546575, -0.5132675, -0.6195013, -0.5907576, 
    -0.6009626, -0.5008821, -0.3698111, -0.173831, -0.08183861, -0.06790638, 
    -0.05644774, -0.02078702, 0.009047031, -0.02085304, -0.0233593, 
    0.008477211, 0.003968716, -0.1011584, -0.251158, -0.39136, -0.5501815, 
    -0.7585149, -1.012242,
  -0.1382512, -0.08279872, 0.01386476, 0.009681821, 0.1037736, 0.09679115, 
    0.06742918, -0.04064369, -0.1099797, -0.1944524, -0.2581729, -0.3053572, 
    -0.3094588, -0.2787133, -0.2301456, -0.1550318, -0.07746017, -0.01160735, 
    0.03263092, 0.07073319, 0.1104467, 0.1447729, 0.1725397, 0.1724095, 
    0.201674, 0.05756581, 0.04080141, 0.07252347, 0.07299554, 0.070131, 
    0.0731746, 0.1111466, 0.1203751, 0.1288712, 0.1186661, 0.1003067, 
    0.07778069, 0.05927485, 0.03912508, 0.02727613, 0.01604566, 0.002064556, 
    -0.01499274, -0.03634691, -0.075149, -0.1112005, -0.1274602, -0.1282415, 
    -0.1330592, -0.1462753, -0.1630885, -0.1795761, -0.1880396, -0.1858913, 
    -0.1832871, -0.1747584, -0.1544622, -0.1370794, -0.1330104, -0.1485214, 
    -0.1684759, -0.2108424, -0.256871, -0.3156113, -0.3788111, -0.4280624, 
    -0.4573105, -0.4783229, -0.4711776, -0.4549178, -0.4075708, -0.3278996, 
    -0.2971216, -0.2381372, -0.2051456, -0.2018741, -0.2106956, -0.1943707, 
    -0.2291689, -0.2280623, -0.2195827, -0.2444524, -0.2711775, -0.2984233, 
    -0.311657, -0.2795119, -0.3103056, -0.3056178, -0.300312, -0.2487988, 
    -0.1784852, -0.148033, -0.1939154, -0.2154322, -0.2128443, -0.1802109,
  0.09970453, 0.1512508, 0.2000626, 0.2334448, 0.2362442, 0.239711, 
    0.2354141, 0.2363907, 0.2418757, 0.2479792, 0.2589167, 0.2811986, 
    0.3047012, 0.3241349, 0.3470352, 0.3600561, 0.3639624, 0.3501765, 
    0.3310357, 0.3010879, 0.2562963, 0.209698, 0.1630834, 0.1298966, 
    0.09630281, 0.08360752, 0.08302158, 0.08495843, 0.08228916, 0.08241937, 
    0.08977614, 0.09928133, 0.107338, 0.1052709, 0.09052483, 0.05850986, 
    0.01918694, -0.0224309, -0.06595303, -0.1058782, -0.1344426, -0.1524276, 
    -0.1654647, -0.1717798, -0.1680364, -0.1805364, -0.1869329, -0.1926783, 
    -0.1987981, -0.2050318, -0.2201197, -0.2436874, -0.2709498, -0.2938827, 
    -0.3261256, -0.3551783, -0.378274, -0.393248, -0.4036158, -0.396845, 
    -0.3746933, -0.3518254, -0.3257024, -0.3040065, -0.2781438, -0.2419948, 
    -0.1998398, -0.1592962, -0.1274602, -0.1092636, -0.09987217, -0.09896076, 
    -0.1034529, -0.1072454, -0.1292018, -0.1660833, -0.1925644, -0.2198105, 
    -0.2008651, -0.2149602, -0.2148626, -0.2236841, -0.2978215, -0.3391463, 
    -0.2693057, -0.2559106, -0.2915715, -0.3188176, -0.2770531, -0.2807155, 
    -0.2439479, -0.1978541, -0.1286483, -0.06273037, -0.001434803, 0.05077873,
  0.2922501, 0.3205379, 0.3731095, 0.3974096, 0.4110327, 0.4215144, 
    0.4221818, 0.4286759, 0.4292618, 0.4331681, 0.4354956, 0.4279272, 
    0.4157039, 0.4141088, 0.3998185, 0.3770646, 0.3614396, 0.3439591, 
    0.3206193, 0.2847957, 0.2586401, 0.2360977, 0.2112768, 0.1838842, 
    0.1550268, 0.1237931, 0.1041316, 0.08567457, 0.05933993, 0.0381648, 
    0.01659904, -0.007440671, -0.02493741, -0.05262294, -0.07394457, 
    -0.1017766, -0.1277694, -0.1545761, -0.1866887, -0.2221216, -0.251565, 
    -0.2808293, -0.3060084, -0.3220077, -0.3376327, -0.3549992, -0.3716007, 
    -0.3862004, -0.3972193, -0.4019719, -0.4063176, -0.4058781, -0.4032902, 
    -0.3982772, -0.3934921, -0.3801457, -0.3718775, -0.3605331, -0.3471868, 
    -0.3389348, -0.3232121, -0.3096054, -0.3082056, -0.3033065, -0.2894882, 
    -0.2802759, -0.270315, -0.2607121, -0.2568547, -0.2618189, -0.2626653, 
    -0.2719263, -0.2772486, -0.2758814, -0.2833196, -0.2871607, -0.2848333, 
    -0.2829127, -0.2782415, -0.2719589, -0.2594426, -0.2394882, -0.2227401, 
    -0.2025741, -0.1805201, -0.1518417, -0.1211614, -0.08590746, -0.05342048, 
    -0.01994067, 0.02392328, 0.06921948, 0.1160457, 0.1679662, 0.2086563, 
    0.2490372,
  -0.06305695, -0.05047584, -0.03963602, -0.03179091, -0.02635473, 
    -0.02433646, -0.02588269, -0.03042371, -0.03696668, -0.04552794, 
    -0.05641657, -0.06912816, -0.07920301, -0.08488333, -0.08751988, 
    -0.08681989, -0.08063507, -0.06999016, -0.05371428, -0.03117204, 
    -0.003128529, 0.02751923, 0.0588994, 0.09047532, 0.1214485, 0.1485481, 
    0.1731083, 0.1925745, 0.2089157, 0.2216275, 0.2326953, 0.2414191, 
    0.2477341, 0.2517542, 0.2539352, 0.2553836, 0.2567344, 0.2589643, 
    0.2632287, 0.26873, 0.2750451, 0.283183, 0.2932905, 0.3039513, 0.3148239, 
    0.3248339, 0.3308233, 0.3368781, 0.3458626, 0.3437142, 0.3588831, 
    0.3619759, 0.3211069, 0.3437626, 0.3533003, 0.3402796, 0.3438766, 
    0.3388474, 0.3211718, 0.2992153, 0.2741666, 0.2789843, 0.2449348, 
    0.2195929, 0.1890265, 0.1557745, 0.120488, 0.08380175, 0.04156542, 
    0.0001591444, -0.03904986, -0.07466173, -0.103096, -0.1180865, 
    -0.1549841, -0.190889, -0.2032751, -0.2217484, -0.2480341, -0.2634475, 
    -0.2710972, -0.2757033, -0.2745314, -0.2719274, -0.264766, -0.2540724, 
    -0.2413771, -0.2251823, -0.2075553, -0.1884475, -0.1686232, -0.1494011, 
    -0.1305699, -0.1114944, -0.09391642, -0.07760763,
  -0.2621132, -0.247774, -0.2283892, -0.2039263, -0.1831744, -0.1663775, 
    -0.1581744, -0.1592323, -0.1685585, -0.1836464, -0.2005897, -0.2140175, 
    -0.2223508, -0.2248898, -0.2205279, -0.2127316, -0.2018593, -0.188106, 
    -0.1749224, -0.1633339, -0.1493039, -0.1283404, -0.1004107, -0.06728899, 
    -0.03433001, -0.00283587, 0.03590131, 0.07957006, 0.1247199, 0.1677215, 
    0.2030079, 0.234225, 0.2555957, 0.2644987, 0.260283, 0.2453414, 
    0.2226201, 0.1953087, 0.1695761, 0.1521609, 0.1374474, 0.1390099, 
    0.1396772, 0.1764936, 0.2061974, 0.1989545, 0.2793256, 0.3204554, 
    0.3462367, 0.3258265, 0.3560349, 0.4139615, 0.3263962, 0.3913541, 
    0.2450483, 0.5042121, 0.5109992, 0.4946581, 0.486227, 0.4808069, 
    0.4890912, 0.4998984, 0.4995731, 0.4856082, 0.4809857, 0.4875613, 
    0.4737104, 0.4463179, 0.4163048, 0.3678347, 0.3248172, 0.2696902, 
    0.2136844, 0.1778934, 0.1321577, 0.100338, 0.07585883, 0.06487253, 
    0.05725533, 0.04952419, 0.06239855, 0.067379, 0.07011336, 0.06529564, 
    0.06495386, 0.04841757, 0.02652627, -0.0003944039, -0.03579479, 
    -0.07681048, -0.1208046, -0.1658404, -0.201843, -0.2307492, -0.2544797, 
    -0.2649778,
  -0.1969276, -0.1873736, -0.1439817, -0.07313202, 0.004146576, 0.07655871, 
    0.1247195, 0.145553, 0.1523889, 0.1478318, 0.1348269, 0.1066856, 
    0.06739527, 0.02799094, 0.003837377, -0.001582548, 0.00894804, 
    0.02206653, 0.03385037, 0.03744739, 0.03507107, 0.03567326, 0.03534776, 
    0.02566352, 0.01135689, -0.0009152293, -0.009378731, -0.0209673, 
    -0.03263736, -0.03760147, -0.0266149, -0.006839514, 0.01252913, 
    0.03285813, 0.05002928, 0.05541682, 0.04568338, 0.01238275, -0.04113293, 
    -0.1104528, -0.1759475, -0.2170286, -0.2238644, -0.2171751, -0.1800005, 
    -0.172009, -0.1303749, -0.0848345, -0.05026424, -0.01937234, 0.02086192, 
    0.06023383, 0.09831977, 0.1428999, 0.178935, 0.1924441, 0.1933718, 
    0.1951784, 0.1811811, 0.1451948, 0.1060346, 0.07133409, 0.05608347, 
    0.05207954, 0.04270454, 0.02821887, 0.02410105, 0.00976184, -0.01439181, 
    -0.03958711, -0.06120169, -0.07796603, -0.06810275, -0.04310274, 
    -0.02848686, -0.0219439, -0.0353879, 0.002714336, -0.00825578, 
    -0.007848978, -0.001436234, 0.0139122, 0.03030217, 0.06872988, 0.1195111, 
    0.1498822, 0.1686323, 0.1705202, 0.1553834, 0.129358, 0.09148395, 
    0.039433, -0.01836306, -0.08096087, -0.1365761, -0.1791054,
  0.1220503, 0.07449186, 0.0177536, -0.01990891, -0.03074861, -0.01276374, 
    0.02167606, 0.05823219, 0.1007289, 0.1365036, 0.1650516, 0.1702598, 
    0.1524864, 0.1171837, 0.07670516, 0.04376251, 0.01872994, -0.008402228, 
    -0.03688529, -0.06642634, -0.08405328, -0.06836319, -0.0300982, 
    0.01218694, 0.02779569, 0.007743597, -0.03006566, -0.05876046, 
    -0.08945698, -0.131026, -0.1687863, -0.1951861, -0.2116249, -0.2236851, 
    -0.2263218, -0.2160842, -0.2112176, -0.2340364, -0.2799025, -0.3339877, 
    -0.3740106, -0.3834181, -0.3543491, -0.2837926, -0.2478876, -0.2867389, 
    -0.3199257, -0.3078814, -0.2902544, -0.2525754, -0.1572466, -0.06491264, 
    0.04635038, 0.1591434, 0.2185183, 0.2364057, 0.2398562, 0.2314253, 
    0.2417768, 0.1866986, 0.129342, 0.08399713, 0.05505824, 0.05813444, 
    0.06843722, 0.0944953, 0.1235969, 0.1211066, 0.1114225, 0.09828758, 
    0.08145809, 0.06220341, 0.04211879, 0.01527953, 0.03289032, 0.07724261, 
    0.0735153, 0.05102146, 0.02387309, -0.04770887, -0.1139198, -0.1768104, 
    -0.2161822, -0.2310746, -0.2233598, -0.1916703, -0.1348343, -0.06336617, 
    0.01759088, 0.04696882, 0.1129029, 0.1653932, 0.1995241, 0.2250938, 
    0.2122684, 0.1717734,
  0.1066693, 0.1285771, 0.09316039, 0.1017382, 0.07729125, 0.06933236, 
    0.07097626, 0.08565736, 0.1433721, 0.1196253, 0.1356089, 0.1533499, 
    0.1653128, 0.1559865, 0.1151984, 0.03266263, -0.04331422, -0.0904007, 
    -0.1683466, -0.2316117, -0.4011264, -0.5687861, -0.6811395, -0.6769404, 
    -0.5990596, -0.4968948, -0.4325229, -0.3904659, -0.3420933, -0.2934444, 
    -0.2586136, -0.2643266, -0.2851924, -0.2922724, -0.2959674, -0.3039101, 
    -0.3293658, -0.370593, -0.4087766, -0.4345253, -0.4230832, -0.3801958, 
    -0.3008502, -0.1981646, -0.1137245, -0.0868853, -0.2091021, -0.3105344, 
    -0.4284869, -0.4860553, -0.4932655, -0.4301307, -0.2879432, -0.119828, 
    0.01809517, 0.1435509, 0.2665164, 0.3261355, 0.3644168, 0.3615522, 
    0.3217084, 0.2773563, 0.2256637, 0.2054324, 0.2258916, 0.258818, 
    0.3215133, 0.4017055, 0.4747359, 0.5359179, 0.4907519, 0.4172002, 
    0.3133591, 0.1881149, 0.09356749, 0.03484344, -0.006237268, 0.04547161, 
    0.1397097, 0.1648561, 0.1340131, 0.09604114, 0.05513945, 0.05308867, 
    0.0431765, 0.03744733, 0.03637302, 0.01205695, -0.02578473, -0.0505569, 
    -0.02886105, -0.1039586, -0.04848993, 0.005807042, 0.06431901, 0.09066999,
  0.2163866, 0.237643, 0.1767542, 0.1847783, 0.1535283, 0.1257128, 
    0.08997023, 0.0161097, -0.04590201, -0.07497096, -0.0885452, -0.09451854, 
    -0.07897496, -0.0226922, 0.03336263, 0.05266595, 0.02779603, 0.03721976, 
    0.08956349, 0.02530539, -0.04350948, -0.2400098, -0.4817257, -0.6242061, 
    -0.636251, -0.5593629, -0.463757, -0.3848348, -0.2882361, -0.1946163, 
    -0.1484573, -0.1179562, -0.1039259, -0.07254577, 0.0205369, 0.09615517, 
    0.09161448, 0.05273104, 0.000305891, -0.03670597, -0.04795277, 
    -0.03704774, -0.002314806, 0.02263641, 0.05328393, 0.07870716, 0.1035281, 
    0.0375125, -0.05604219, -0.1947466, -0.2865109, -0.2690142, -0.1582232, 
    -0.03703183, 0.06173122, 0.1853315, 0.3210248, 0.4390588, 0.524394, 
    0.5873172, 0.6414838, 0.6723758, 0.6605268, 0.6354942, 0.6111616, 
    0.5882612, 0.5960574, 0.6717247, 0.785771, 0.8346479, 0.8451948, 
    0.8040978, 0.6908816, 0.5344038, 0.3918094, 0.320439, 0.3200157, 
    0.3444949, 0.3480756, 0.4955366, 0.5054976, 0.4846804, 0.4234337, 
    0.3870893, 0.3858035, 0.3925255, 0.4059044, 0.4155722, 0.4080528, 
    0.3699994, 0.306474, 0.2097621, 0.1059698, 0.04143524, 0.05831385, 
    0.1334276,
  0.6766075, 0.7531701, 0.7386032, 0.6870245, 0.5556933, 0.3963345, 
    0.2283005, 0.1826137, 0.2059209, 0.2338181, 0.2712367, 0.3096808, 
    0.3350713, 0.3606412, 0.4269171, 0.480628, 0.4957974, 0.5098109, 
    0.5872524, 0.681914, 0.7013963, 0.5954393, 0.448076, 0.2630501, 
    0.1800258, 0.1008105, 0.04893875, 0.02271795, 0.04939437, 0.06013656, 
    0.07288098, 0.1120572, 0.2234342, 0.3248177, 0.4412074, 0.5208626, 
    0.5144823, 0.5399543, 0.4689256, 0.4308559, 0.4206182, 0.4170864, 
    0.4242963, 0.4485315, 0.4863406, 0.5411746, 0.6592247, 0.7074018, 
    0.6898399, 0.5887332, 0.5242637, 0.5264611, 0.5537884, 0.6113406, 
    0.6567019, 0.6599737, 0.6518681, 0.6431605, 0.7090622, 0.8263962, 
    0.9021285, 1.143665, 1.446921, 1.671432, 1.757532, 1.806051, 1.822539, 
    1.921709, 1.943502, 1.872929, 1.76847, 1.707435, 1.745228, 1.751836, 
    1.598987, 1.327584, 1.129554, 1.00527, 0.9673302, 0.9563439, 0.8856082, 
    0.9421999, 1.012561, 1.035201, 0.9770958, 0.8623497, 0.8052371, 
    0.8706668, 0.9962364, 1.125973, 1.169934, 1.063538, 0.8836713, 0.7099082, 
    0.6327274, 0.6171024,
  1.097587, 1.093177, 1.146578, 1.188489, 1.204456, 1.139563, 1.139775, 
    1.204293, 1.202519, 1.17275, 1.060413, 0.9186975, 0.84902, 0.8597133, 
    0.9585903, 1.061455, 1.080091, 0.9542117, 0.8106732, 0.7322553, 0.768144, 
    0.9028607, 0.973157, 0.9773725, 1.049899, 1.172115, 1.206149, 1.227226, 
    1.267167, 1.442542, 1.715052, 1.99303, 2.158379, 2.22052, 2.163554, 
    2.066565, 1.965979, 1.888717, 1.76344, 1.64054, 1.536585, 1.457369, 
    1.388489, 1.291093, 1.193567, 1.12843, 1.110478, 1.114254, 1.087708, 
    1.036064, 0.9906701, 1.011048, 1.130319, 1.285153, 1.408558, 1.520081, 
    1.596009, 1.631962, 1.577259, 1.521237, 1.515996, 1.566077, 1.747766, 
    1.986308, 2.146741, 2.234746, 2.299313, 2.380823, 2.500273, 2.573727, 
    2.557386, 2.534762, 2.536438, 2.45719, 2.370813, 2.327242, 2.276331, 
    2.202291, 2.083118, 1.904765, 1.764954, 1.711878, 1.782207, 1.924345, 
    2.020814, 2.010967, 1.923385, 1.87944, 1.838847, 1.798336, 1.792233, 
    1.76388, 1.62944, 1.406686, 1.22166, 1.131149,
  1.833737, 1.772995, 1.845342, 2.061846, 2.368811, 2.631116, 2.809485, 
    2.987269, 3.07874, 3.026673, 2.867331, 2.712643, 2.610966, 2.586064, 
    2.593812, 2.6165, 2.593486, 2.513961, 2.372522, 2.204261, 2.125989, 
    2.093095, 2.153089, 2.278887, 2.399297, 2.54041, 2.630807, 2.641305, 
    2.554814, 2.53831, 2.733134, 3.10973, 3.389108, 3.464238, 3.426836, 
    3.390312, 3.422685, 3.402568, 3.256035, 2.97957, 2.741663, 2.633411, 
    2.612789, 2.588294, 2.547278, 2.464677, 2.375371, 2.279277, 2.135722, 
    1.95802, 1.837041, 1.800647, 1.824296, 1.90929, 2.018144, 2.093828, 
    2.172132, 2.251966, 2.319837, 2.331653, 2.181588, 1.99775, 1.987382, 
    2.128381, 2.251526, 2.320015, 2.453853, 2.655708, 2.797733, 2.847489, 
    2.915816, 2.988098, 2.962414, 2.928365, 3.016891, 3.231506, 3.328918, 
    3.223254, 3.148156, 3.136666, 3.006424, 2.72581, 2.506393, 2.47415, 
    2.549394, 2.659843, 2.812806, 2.837171, 2.715166, 2.643584, 2.678675, 
    2.727991, 2.603626, 2.356751, 2.155042, 2.008346,
  2.36733, 2.369706, 2.380839, 2.457873, 2.596643, 2.763684, 2.984892, 
    3.217476, 3.468795, 3.708833, 3.710851, 3.53997, 3.393762, 3.378088, 
    3.39246, 3.384517, 3.370064, 3.347701, 3.322066, 3.244771, 3.141923, 
    3.032076, 2.877909, 2.776281, 2.763407, 2.82065, 2.985949, 3.151314, 
    3.204748, 3.138619, 3.074735, 3.155757, 3.373173, 3.575777, 3.756034, 
    3.96261, 4.225679, 4.406083, 4.409778, 4.216711, 3.946415, 3.70203, 
    3.618192, 3.714449, 3.804976, 3.70758, 3.492834, 3.191385, 2.926363, 
    2.718013, 2.51274, 2.317932, 2.169088, 2.051802, 1.958817, 1.963375, 
    2.09508, 2.291532, 2.438911, 2.517281, 2.415458, 2.238163, 2.136047, 
    2.169055, 2.219121, 2.204227, 2.268274, 2.456848, 2.605481, 2.653105, 
    2.692672, 2.812707, 2.869185, 2.838619, 2.851136, 2.779781, 2.532418, 
    2.334306, 2.465979, 2.812902, 3.100354, 3.117639, 3.022733, 2.962398, 
    2.831897, 2.717867, 2.745129, 2.802567, 2.89189, 3.047961, 3.126217, 
    3.046431, 2.875679, 2.697489, 2.527356, 2.405155,
  2.727438, 2.712301, 2.667346, 2.573255, 2.457939, 2.44705, 2.515068, 
    2.604554, 2.773727, 3.063831, 3.245586, 3.258818, 3.217786, 3.151885, 
    3.123255, 3.160755, 3.250175, 3.297246, 3.249492, 3.136927, 3.115817, 
    3.063864, 2.908476, 2.787692, 2.772913, 2.821855, 2.92594, 3.076347, 
    3.216777, 3.339499, 3.351543, 3.220943, 3.251999, 3.478252, 3.625729, 
    3.713602, 3.875648, 4.034192, 4.117118, 4.155464, 4.071415, 3.784485, 
    3.53883, 3.456897, 3.366679, 3.223417, 3.086389, 2.991744, 2.927063, 
    2.876542, 2.738017, 2.464807, 2.183183, 2.032889, 1.956083, 1.9144, 
    1.907352, 1.90592, 1.905432, 1.909257, 1.847115, 1.763554, 1.645993, 
    1.649215, 1.747067, 1.824736, 1.84233, 1.909111, 2.032581, 2.175176, 
    2.232321, 2.196888, 2.110169, 2.093144, 2.052503, 1.752617, 1.378658, 
    1.474361, 1.900126, 2.149297, 2.111129, 2.093372, 2.205221, 2.331686, 
    2.403577, 2.450371, 2.45286, 2.378317, 2.397572, 2.597408, 2.795618, 
    2.841077, 2.825273, 2.808541, 2.777259, 2.726249,
  1.931637, 1.866142, 1.815702, 1.746009, 1.636975, 1.558606, 1.591044, 
    1.655123, 1.732922, 1.813717, 1.865507, 1.949377, 2.034208, 2.058003, 
    2.102454, 2.169414, 2.197864, 2.212497, 2.221383, 2.256214, 2.352617, 
    2.389042, 2.278723, 2.148385, 2.083671, 1.999866, 1.893844, 1.841387, 
    1.853431, 1.966224, 2.124849, 2.141809, 2.153853, 2.295227, 2.344413, 
    2.354554, 2.45732, 2.537984, 2.613929, 2.768535, 2.870602, 2.813082, 
    2.598417, 2.218974, 1.925534, 1.924329, 2.008069, 2.156832, 2.297147, 
    2.471773, 2.570601, 2.423368, 2.271529, 2.24788, 2.216386, 2.101965, 
    1.856946, 1.528381, 1.275713, 1.129814, 1.074736, 1.044902, 0.8945928, 
    0.7171516, 0.6801233, 0.684062, 0.7168255, 0.8109012, 1.001803, 1.200729, 
    1.398043, 1.505188, 1.473434, 1.454798, 1.407207, 0.9551072, 0.4411583, 
    0.3491173, 0.4582314, 0.2952437, 0.3843875, 0.7696738, 1.030123, 
    1.132158, 1.293095, 1.49137, 1.581018, 1.537854, 1.478333, 1.539384, 
    1.726135, 1.922799, 2.046187, 2.054651, 2.020308, 1.983363,
  1.068029, 1.002925, 0.9168901, 0.8195276, 0.7035599, 0.6077271, 0.5241985, 
    0.4047155, 0.3072386, 0.3004189, 0.327014, 0.3998499, 0.5347614, 
    0.6803188, 0.8349085, 0.9758587, 1.063976, 1.152633, 1.222766, 1.246822, 
    1.235186, 1.183785, 1.049735, 0.8323526, 0.6147261, 0.4096622, 0.169982, 
    0.01018333, -0.08517742, -0.1254282, -0.07386589, -0.07770634, 
    -0.1037483, -0.02594757, 0.1143837, 0.3643513, 0.4845829, 0.4887486, 
    0.7701292, 1.015345, 0.9666305, 0.9418907, 1.083444, 1.077356, 0.9299283, 
    0.8437791, 0.7630005, 0.7055135, 0.8170204, 1.081897, 1.302926, 1.331083, 
    1.32288, 1.282792, 1.201103, 1.125924, 0.9758911, 0.8338175, 0.6713986, 
    0.4195766, 0.2485967, 0.2419558, 0.1917443, 0.07704687, -0.02847052, 
    -0.09665108, -0.1119342, -0.04572344, 0.07091141, 0.1109343, 0.1823859, 
    0.4339323, 0.4503384, 0.2256799, 0.06187773, -0.1670933, -0.3774776, 
    -0.6464391, -1.121748, -1.349678, -1.05985, -0.7127476, -0.5518589, 
    -0.4383011, -0.3017941, -0.186039, -0.05239677, 0.1928353, 0.4638629, 
    0.5815883, 0.7073693, 0.9480915, 1.12625, 1.218258, 1.241321, 1.167346,
  0.0742631, -0.03774834, -0.1920452, -0.3524127, -0.6156616, -0.8834672, 
    -1.035306, -1.155668, -1.313302, -1.355294, -1.172953, -0.9556847, 
    -0.8116741, -0.7032919, -0.6213908, -0.4728231, -0.2760782, -0.1514206, 
    -0.1657915, -0.2480507, -0.2952194, -0.3482466, -0.3843956, -0.5285521, 
    -0.7122602, -0.8330774, -1.140759, -1.4981, -1.692176, -1.90627, 
    -2.108923, -2.297839, -2.34823, -2.181515, -2.030749, -1.755342, 
    -1.515986, -1.402819, -1.099711, -0.7980342, -0.8784051, -0.7799349, 
    -0.594193, -0.5644727, -0.6118202, -0.621016, -0.5252314, -0.4858594, 
    -0.5516634, -0.4364295, -0.2456741, -0.09801769, 0.01661444, -0.0182004, 
    -0.08538771, -0.07680988, -0.05130625, -0.008320808, 0.01096582, 
    -0.0883832, -0.2442913, -0.3286176, -0.4295449, -0.5412965, -0.6408572, 
    -0.6969762, -0.7436233, -0.8553095, -0.8411822, -0.7880244, -0.8702998, 
    -0.8890662, -0.8639846, -0.8023472, -0.9285841, -1.187471, -0.9235384, 
    -0.8919632, -1.559004, -1.552722, -1.041492, -1.293949, -1.473897, 
    -1.487894, -1.577493, -1.443347, -1.231431, -0.9399605, -0.6508007, 
    -0.4663448, -0.2808304, -0.1385293, -0.06885099, 0.05398369, 0.1660771, 
    0.1286583,
  -0.8297234, -0.8505726, -0.9443064, -1.194746, -1.624417, -2.066687, 
    -2.423767, -2.366263, -2.136511, -2.167988, -2.174043, -2.142125, 
    -2.096096, -2.03747, -2.013268, -1.87943, -1.743721, -1.654821, 
    -1.580977, -1.572904, -1.524141, -1.487878, -1.439408, -1.456531, 
    -1.602966, -1.670756, -1.852071, -2.145299, -2.410892, -2.943443, 
    -3.50054, -3.933792, -4.026745, -3.555782, -3.323653, -3.154952, 
    -2.529853, -1.6703, -1.150378, -1.324548, -1.395544, -1.059021, 
    -1.011446, -1.227933, -1.432441, -1.618183, -1.695071, -1.806253, 
    -1.906448, -1.816166, -1.698587, -1.654887, -1.567224, -1.423978, 
    -1.239717, -1.073881, -0.8717971, -0.6317418, -0.5466995, -0.6065459, 
    -0.7570672, -0.9267774, -1.016117, -1.057621, -1.198636, -1.33586, 
    -1.384688, -1.436527, -1.398522, -1.412113, -1.461966, -1.517988, 
    -1.645723, -1.443981, -1.228812, -1.044421, -0.2227739, -0.02521491, 
    -1.165564, -1.145528, -0.6929072, -1.229626, -1.437487, -1.817826, 
    -2.047546, -1.663578, -1.424092, -1.253177, -1.104007, -1.072432, 
    -1.029056, -1.012942, -1.045869, -1.010192, -0.9715528, -0.9237175,
  -1.140531, -1.140352, -1.08446, -1.056319, -0.8093951, -0.6378944, 
    -0.9277707, -1.108142, -0.8983925, -1.343672, -1.950427, -2.273392, 
    -2.361755, -2.290385, -2.245056, -2.126534, -2.058728, -1.96475, 
    -1.732913, -1.629251, -1.521081, -1.459134, -1.482116, -1.45946, 
    -1.559151, -1.665824, -1.814847, -2.086739, -2.361544, -2.654154, 
    -2.447204, -2.387064, -2.451663, -1.978975, -1.764164, -1.68586, 
    -1.568461, -1.244275, -0.8738482, -1.234916, -1.505147, -1.133777, 
    -1.175834, -1.417745, -1.683288, -2.075394, -2.44823, -2.664294, 
    -2.681628, -2.609363, -2.59294, -2.499352, -2.277478, -2.07668, 
    -1.712667, -1.359411, -1.200769, -0.9502154, -0.8065794, -0.8353065, 
    -0.9127316, -1.012243, -1.171391, -1.299402, -1.35754, -1.449353, 
    -1.591784, -1.686836, -1.644958, -1.660941, -1.552445, -1.372237, 
    -1.470202, -1.48586, -1.191768, -0.6575071, 0.2345828, 0.5077603, 
    -0.428438, -0.5412145, -0.3079951, -0.7846389, -0.9526887, -1.252738, 
    -1.56501, -1.28892, -1.215629, -1.170349, -1.167321, -1.142142, -1.13791, 
    -1.159867, -1.191051, -1.194095, -1.107979, -1.095462,
  -1.009313, -0.9281936, -0.7444048, -0.338171, 0.1542281, 0.2390262, 
    -0.03281635, -0.3450884, -0.4188349, -0.5529494, -1.056091, -1.550215, 
    -1.737634, -1.650834, -1.428031, -1.360322, -1.343493, -1.264441, 
    -1.107035, -1.019649, -0.9896032, -1.002803, -1.132897, -1.141035, 
    -1.168786, -1.255586, -1.244095, -1.329919, -1.326973, -1.075964, 
    -0.5460488, -0.7883013, -1.393249, -1.26457, -1.344697, -1.090824, 
    -0.8377643, -0.983272, -0.8261268, -0.9168007, -1.166166, -1.072822, 
    -1.271276, -1.544258, -1.719519, -1.808744, -1.92279, -2.083793, 
    -2.209802, -2.233549, -2.17961, -2.177526, -2.038936, -1.908467, 
    -1.611315, -1.176142, -1.066849, -1.055635, -0.9370153, -0.9119339, 
    -1.075508, -1.175264, -1.334558, -1.44224, -1.439017, -1.458272, 
    -1.532767, -1.692239, -1.631872, -1.617288, -1.581237, -1.445657, 
    -1.187129, -1.030276, -0.7139196, -0.232816, -0.2448117, 0.2742479, 
    0.1411583, -0.2878127, -0.08991265, -0.04891312, -0.1272334, -0.2905473, 
    -0.8738806, -1.244079, -0.9946975, -0.9389524, -1.271423, -1.288073, 
    -1.302152, -1.264848, -1.18682, -1.176713, -1.111804, -1.03542,
  -0.5640502, -0.3495483, -0.07503605, 0.5141568, 0.6445925, -0.04551136, 
    -0.3088902, -0.5264522, -0.5610385, -0.1641796, -0.09573913, -0.1167514, 
    -0.4136264, -0.6646037, -0.6934609, -0.7724319, -0.7554886, -0.6369333, 
    -0.5634472, -0.5269887, -0.6003129, -0.6352091, -0.6501503, -0.6810913, 
    -0.5854211, -0.5460491, -0.4941444, -0.3722863, -0.05098009, 0.482044, 
    0.7812298, 0.2581505, -0.5233757, -0.5778193, -0.8682973, -0.8727245, 
    -0.5150751, -0.4947627, -0.3722366, -0.6207067, -1.115563, -1.15002, 
    -1.056286, -0.9533081, -0.9095583, -0.8843141, -0.9192424, -1.053845, 
    -1.150997, -1.202413, -1.229529, -1.377462, -1.354464, -1.208777, 
    -1.280277, -1.297921, -1.266264, -1.222107, -1.113741, -1.054285, 
    -1.210893, -1.316427, -1.389637, -1.301404, -1.270333, -1.322481, 
    -1.331385, -1.447725, -1.432263, -1.443119, -1.208272, -1.105229, 
    -0.8313026, -0.5086794, -0.1585655, 0.319577, -0.3976275, 0.08894503, 
    0.5256146, -0.4490435, -0.2201698, 0.06122661, -0.08175802, -0.03703177, 
    -0.5182327, -1.138399, -1.127624, -0.9307002, -1.275541, -1.314391, 
    -1.37017, -1.232637, -1.083842, -0.9544635, -0.8490109, -0.7581744,
  -0.1648479, 0.03562498, 0.1131477, 0.5307907, 0.9499639, 0.2570928, 
    0.04747367, -0.1590853, -0.4991734, -0.2669468, -0.06294298, 0.3217736, 
    0.1964643, -0.2926791, -0.4227734, -0.3420935, -0.3979049, -0.461267, 
    -0.3951044, -0.2630892, -0.2362504, -0.2324581, -0.2084513, -0.1968141, 
    -0.05192471, 0.07193661, 0.1350713, 0.3102341, 0.5694141, 0.7407191, 
    0.8446577, 0.7268354, 0.3278936, -0.1935258, -0.3795123, -0.3821812, 
    -0.2472529, -0.03273493, -0.2597365, -0.6763055, -0.7865925, -0.7494993, 
    -0.4161339, -0.1734738, 0.05544901, 0.1278119, 0.1013799, -0.08864307, 
    -0.4320998, -0.7611527, -0.8624387, -0.9125528, -1.18184, -1.351615, 
    -1.473458, -1.494438, -1.395854, -1.271635, -1.196798, -1.10002, 
    -1.010111, -0.8580608, -0.8817582, -0.8993692, -0.9313183, -0.9141965, 
    -0.9633822, -1.045805, -0.9798379, -1.01527, -0.7519894, -0.6349645, 
    -0.3984413, -0.02786827, 0.0751586, 0.3515587, -0.05290091, 0.1279423, 
    0.3064415, -0.3628128, -0.4367714, -0.3382523, -0.3760782, -0.3425494, 
    -0.3345739, -1.059281, -1.102738, -0.8393428, -1.037601, -0.9681189, 
    -1.012569, -0.8686399, -0.7927284, -0.568933, -0.4073606, -0.3168173,
  0.1290331, 0.2206836, 0.01803029, -0.06240594, 0.4008104, 0.194381, 
    0.1580529, 0.233639, -0.06924152, -0.3927116, -0.4792678, 0.02325463, 
    0.2421674, -0.02454782, -0.003209591, 0.1648726, 0.02916288, -0.1580276, 
    -0.06735373, 0.03342724, 0.2009239, 0.1582971, 0.08966112, 0.2380662, 
    0.2563276, 0.3498821, 0.4315557, 0.4870734, 0.5910449, 0.6852016, 
    0.6267378, 0.8574018, 0.9378871, 0.5349897, 0.3308393, 0.2447069, 
    0.1680961, 0.3723106, 0.1547983, -0.1843133, 0.06780195, 0.4747357, 
    0.6498008, 0.6097455, 0.8718553, 0.7936163, 0.4938602, 0.3023891, 
    -0.0293498, -0.3916383, -0.7235718, -0.8846555, -1.074646, -1.303829, 
    -1.27629, -1.081661, -1.060681, -0.9970417, -0.8701372, -0.699955, 
    -0.6043658, -0.5158238, -0.5290723, -0.5248246, -0.5819211, -0.5175333, 
    -0.4842978, -0.4935417, -0.5406127, -0.5067415, -0.445837, -0.3049192, 
    -0.1092162, 0.02209854, 0.02377558, 0.2692345, 0.468144, 0.3873177, 
    0.1385704, 0.003430367, -0.2817909, -0.5204628, -0.3636105, -0.2749872, 
    -0.2891963, -1.083158, -0.9593954, -0.5762081, -0.8542032, -0.6008019, 
    -0.5616407, -0.4229856, -0.2872758, -0.1965532, -0.1078811, 0.0243125,
  0.1705368, 0.2206668, 0.1592085, -0.05709982, 0.1376593, 0.2367963, 
    0.2214643, 0.391435, 0.3481081, -0.05566764, -0.5182486, -0.3151886, 
    0.0858686, 0.03536463, 0.259876, 0.5902476, 0.5050907, 0.1994591, 
    0.1267867, 0.2133427, 0.3796024, 0.4285932, 0.3147745, 0.30164, 0.353219, 
    0.4896121, 0.491663, 0.5072563, 0.4559209, 0.4915326, 0.5075808, 
    0.5054163, 0.5877736, 0.6414838, 0.6077437, 0.4944137, 0.3185349, 
    0.5668256, 0.6334281, 0.3040004, 0.5581834, 0.8120251, 0.9530566, 
    0.9592578, 1.049541, 1.367103, 1.090687, 1.03058, 0.847018, 0.5021617, 
    -0.09609747, -0.7140172, -0.8383992, -0.6580443, -0.5777225, -0.5645714, 
    -0.4613967, -0.2975788, -0.2535515, -0.1949906, -0.2540727, -0.2799034, 
    -0.3349156, -0.2541213, -0.259655, -0.2380729, -0.3090854, -0.2153363, 
    -0.2752643, -0.2012405, -0.2655959, -0.1629267, -0.1244345, -0.1179073, 
    0.1449994, 0.165377, 0.1925256, 0.03199491, -0.02612683, 0.02597278, 
    -0.08581107, -0.2655473, -0.3639524, -0.2824908, -0.1612178, -0.8502159, 
    -0.5626011, -0.1058307, -0.2665563, -0.1404333, -0.1411819, 
    -0.0006217957, 0.01920176, 0.07540274, 0.1712203, 0.1896291,
  0.1655886, 0.1012006, 0.08887982, 0.04215169, 0.1383431, 0.01197565, 
    -0.1369016, -0.03309315, 0.1422488, -0.0567584, -0.4018099, -0.3196166, 
    -0.255928, -0.6016148, -0.2670608, 0.1774218, 0.5756476, 0.4476039, 
    0.2827439, 0.3835568, 0.4531217, 0.6238408, 0.5819302, 0.4200974, 
    0.4227018, 0.450078, 0.3415008, 0.3412398, 0.3551231, 0.1376752, 
    0.05338216, 0.06558943, -0.08196974, 0.08585286, 0.374492, 0.4448047, 
    0.5020307, 0.2757776, 0.225159, 0.1337366, 0.7059696, 0.8042121, 
    1.146578, 1.290035, 0.8940392, 1.426054, 1.251233, 1.085429, 0.9470502, 
    0.5919883, 0.2388475, -0.2930861, -0.9106483, -0.8893917, -0.6270547, 
    -0.5534711, -0.3651404, -0.1399937, -0.0363965, 0.01707029, -0.167696, 
    -0.170414, -0.2071486, -0.1491246, -0.2329788, -0.1343951, -0.2013054, 
    -0.1054397, -0.1509638, -0.1862674, -0.1609249, -0.1688023, -0.1971717, 
    -0.1710811, -0.1013547, -0.1768591, -0.1021848, -0.1018592, -0.04831107, 
    -0.1346229, -0.1900755, -0.1858273, -0.2959186, -0.4698931, -0.3227901, 
    -0.3274448, -0.3954141, -0.1400104, 0.02530527, 0.06042957, 0.1081014, 
    0.2067022, 0.1328745, 0.2393525, 0.1616666, 0.1958297,
  0.01978785, -0.1218623, -0.153584, -0.05524421, 0.1350229, -0.05819011, 
    -0.06722397, -0.00753963, 0.141256, -0.1014034, -0.3257196, -0.5631869, 
    -0.7423049, -0.5009478, -0.2322792, -0.1739784, 0.3276167, 0.36165, 
    0.2279103, 0.0635221, 0.2094529, 0.5028286, 0.6471319, 0.5062304, 
    0.310348, 0.3753543, 0.3324506, -0.2248898, -0.1618527, -0.06981158, 
    -0.2826855, -0.3174024, -0.3806839, -0.2767289, 0.2142543, 0.3345178, 
    0.3798139, 0.04792917, -0.03302787, 0.1304324, 0.7171187, 0.7399213, 
    1.110755, 1.473141, 1.151233, 1.236097, 0.9948693, 0.9407676, 0.9166465, 
    0.6611128, 0.4877895, 0.5817187, 0.2004528, 0.1404586, 0.250843, 
    0.3493776, 0.3717575, 0.4758101, 0.5473924, 0.6049771, 0.5091925, 
    0.4125943, 0.141777, 0.1422162, 0.02244091, -0.01833057, -0.05895519, 
    -0.03755283, -0.04889679, -0.08131886, -0.1190298, -0.1831574, 
    -0.2686396, -0.2086464, -0.2029009, 0.05206323, -0.1215208, -0.07555716, 
    -0.03003308, -0.02571994, -0.07165092, -0.1492551, -0.157263, -0.363871, 
    -0.2833043, 0.07201791, -0.1055374, 0.001704693, 0.2768524, 0.419642, 
    0.4091115, 0.3535609, 0.3736784, 0.3711554, 0.1141402, 0.1635705,
  -0.07156932, -0.1257684, -0.08877301, 0.01506782, 0.002877355, -0.0514037, 
    -0.04700899, -0.0903521, 0.1344038, 0.2331182, 0.1958137, -0.3115107, 
    -0.6560743, -0.2298868, 0.1684369, 0.485185, 0.5365847, 0.2237755, 
    0.2447065, -0.007360578, 0.132532, 0.3683556, 0.5894656, 0.4813601, 
    0.3236454, 0.2954224, 0.4023074, -0.05058971, -0.1631385, -0.107344, 
    -0.04578847, -0.11252, -0.04850639, -0.007946491, 0.1968223, 0.1028607, 
    0.05181912, 0.03552681, 0.03049751, 0.3214155, 0.2846316, 0.03655221, 
    0.1833296, 0.5190555, 0.7190717, 0.7178022, 0.8053023, 0.9298468, 
    0.8518686, 0.9061821, 0.650892, 0.7246222, 0.6480923, 0.7829232, 
    0.7811975, 0.9204226, 0.9132943, 1.051038, 0.97472, 0.8536582, 0.8152471, 
    0.7970834, 0.6301885, 0.5460901, 0.4382615, 0.3888965, 0.3831511, 
    0.3597465, 0.2572718, 0.226608, 0.03432238, 0.03754503, -0.1283404, 
    -0.2637244, -0.3324904, 0.08635712, 0.03316677, 0.05216093, 
    -0.0008013099, -0.008809119, 0.01606068, -0.3949909, -0.2105669, 
    -0.2286006, -0.214798, -0.05973673, -0.08154726, 0.2067354, 0.3471646, 
    0.4935021, 0.4338343, 0.4545046, 0.4357221, 0.4431603, 0.3103152, 
    0.2001752,
  -0.03231156, -0.141377, -0.2813022, 0.01931584, 0.01449817, -0.02161837, 
    -0.03411837, 0.0188927, 0.3772423, 0.2586066, 0.3623662, 0.2254689, 
    -0.07223654, 0.2232065, 0.621725, 0.9124637, 0.6993289, 0.3349082, 
    0.5026329, 0.3109503, 0.3296515, 0.4262009, 0.5483035, 0.3006961, 
    0.3937137, 0.1389613, 0.03507096, -0.1916867, -0.4916865, -0.5258827, 
    -0.06305717, -0.03903373, -0.02585014, 0.09073517, 0.004048947, 
    0.1563764, 0.1169233, 0.09937769, 0.005660117, 0.1437788, -0.08748734, 
    -0.2880895, -0.2316277, -0.1512725, 0.01160121, -0.08319044, -0.1773798, 
    -0.1111853, -0.05924845, 0.1988082, 0.1058235, 0.1711068, 0.1048784, 
    0.2587523, 0.3220015, 0.5370083, 0.5685024, 0.7675095, 0.7967415, 
    0.8849897, 0.7459602, 0.5980759, 0.5169563, 0.5208137, 0.4911916, 
    0.4826298, 0.4382288, 0.4805303, 0.4118619, 0.4593874, 0.2675906, 
    0.2348595, 0.1104293, -0.02580142, -0.2193553, 0.1925743, 0.3033001, 
    -0.1173378, 0.1189741, 0.02320588, -0.2577021, -0.193298, -0.4119011, 
    -0.4062696, -0.5384479, -0.3381877, -0.1820512, -1.978874e-005, 
    0.04019809, 0.2285122, 0.1951784, 0.1987917, 0.1247032, 0.3111615, 
    0.2375289, 0.071383,
  0.000272911, -0.1003456, 0.06555605, 0.02335232, 0.183183, 0.1892703, 
    0.1537234, 0.2413698, 0.1644656, -0.001826704, 0.09462512, 0.3185513, 
    0.3132942, 0.3551884, 0.7118454, 0.8971646, 0.8533335, 0.9347627, 
    1.125128, 1.02249, 1.003822, 0.6618459, 0.6956506, 0.4447563, 0.6101527, 
    0.3355433, 0.09550405, -0.3774127, -0.4572959, -0.4165244, -0.1824577, 
    -0.2747923, -0.2663286, -0.3573767, -0.549906, -0.02127635, -0.08673811, 
    -0.1941767, -0.2310908, -0.1721551, -0.1290884, -0.1681676, -0.1325235, 
    -0.06128263, -0.09565783, -0.2147498, -0.4405632, -0.4118037, -0.4350462, 
    -0.6052933, -0.7355995, -0.6786008, -0.8246455, -0.8617225, -0.9877639, 
    -1.009396, -0.9519248, -0.9242387, -0.9518762, -0.7906942, -0.7168336, 
    -0.5587931, -0.4690628, -0.2614293, -0.1688187, -0.02829123, 0.09128928, 
    0.3044403, 0.3192837, 0.3886523, 0.2447228, 0.1587366, 0.0957973, 
    0.1166141, 0.07222962, 0.1789513, 0.4949837, -0.261055, 0.2353803, 
    -0.2814977, -0.4908726, -0.4372759, -0.3990107, -0.4703975, -0.4372592, 
    -0.08992863, 0.05038691, 0.1835737, 0.1980109, 0.3551724, 0.2580044, 
    0.2821088, 0.4398563, 0.4808067, 0.07556588, 0.01313099,
  -0.05708385, -0.1041051, -0.06686544, 0.04001927, 0.1539513, 0.2002078, 
    0.2200973, 0.08123004, 0.02851184, 0.2304161, 0.1627891, 0.2257615, 
    0.3272429, 0.07462168, 0.4713993, 0.7941046, 0.8026662, 0.9613414, 
    1.105906, 1.119333, 1.058428, 0.2529593, 0.3948855, 0.6317663, 0.484664, 
    0.5426879, 0.5675259, -0.1732295, -0.1157432, -0.2377152, -0.2562213, 
    -0.04554415, 0.113652, -0.07487357, -0.06842804, 0.08536458, -0.2189817, 
    -0.197432, -0.03315783, 0.05846024, -0.07982111, -0.2059121, -0.1526732, 
    0.01729727, -0.1421261, -0.1197958, -0.11973, 0.0009069443, 0.06158447, 
    -0.01142979, -0.02407646, -0.07436848, -0.1643915, -0.2640343, 
    -0.3400106, -0.4144573, -0.4351282, -0.4614458, -0.4769897, -0.3963094, 
    -0.4041705, -0.2721882, -0.2870803, -0.1269407, -0.2182488, -0.04902697, 
    0.1367798, 0.4974737, 0.6762991, 0.8101039, 1.105123, 1.412317, 
    0.8330207, 0.1027799, 0.1301557, 0.2908816, 0.2091924, -0.2927928, 
    -0.3117547, -0.906498, -0.9002476, -0.4754438, -0.3804722, -0.08042336, 
    0.02927637, 0.2949023, 0.4317832, 0.6468062, 0.6894817, 0.797246, 
    0.7852666, 0.9532026, 1.066337, 0.4776818, 0.1008265, 0.06889284,
  -0.2634799, -0.301924, -0.2150264, -0.07659793, -0.1200886, -0.08789372, 
    0.04307938, 0.03490853, 0.1786583, 0.466549, 0.202389, -0.01450551, 
    0.04500008, 0.04975224, 0.3675261, 0.4837852, 0.5042281, 0.6347461, 
    0.6716118, 0.7252407, 0.8461226, 0.365557, 0.7573862, 0.9996219, 0.57651, 
    1.097425, 0.9747038, 0.3630176, 0.1608202, 0.1460903, 0.4058723, 
    0.5964479, 0.4863734, 0.005856037, 0.2627077, 0.2908978, 0.3103156, 
    0.4023724, 0.2465615, 0.317574, 0.1430135, 0.1387825, 0.2215128, 
    0.3181601, 0.1587038, 0.07561398, 0.1145144, 0.3001099, 0.4708929, 
    0.5385208, 0.4838982, 0.3932896, 0.3820105, 0.26614, 0.3694935, 
    0.5380487, 0.6127548, 0.5742788, 0.4109812, 0.3815384, 0.2522745, 
    0.1797647, 0.2187462, 0.3136358, 0.2770472, 0.3203249, 0.2493453, 
    0.6054819, 0.885169, 1.150436, 1.52, 1.508363, 0.69679, 0.2666144, 
    0.9119749, 0.7501087, 0.3315058, -0.1854706, -0.6038771, -0.5433793, 
    -0.3472862, -0.2110229, -0.08260441, -0.05579758, 0.05891562, 0.3873172, 
    0.5623336, 0.6761999, 0.7337041, 0.8125291, 0.9396777, 0.9812467, 
    0.5008104, 0.1983693, -0.08421564, -0.0516634,
  -0.4015656, -0.4141476, -0.2187047, 0.0005497932, -0.1516638, -0.2516475, 
    -0.0357461, 0.2073371, 0.3138146, 0.5211713, 0.3883751, 0.04110944, 
    -0.04878235, 0.06910443, 0.2145633, 0.3197885, 0.3368611, 0.337822, 
    0.3290653, 0.4517221, 0.4981574, 0.1096482, 0.4599898, 0.5252409, 
    0.4301074, 0.8794559, 0.2982874, 0.1204717, 0.1481571, 0.3839972, 
    0.5960252, 0.6334763, 1.000257, 0.5365691, 0.4586229, 0.4590778, 
    0.5681767, 0.5848756, 0.3824177, 0.4145145, 0.4191527, 0.5354939, 
    0.4692836, 0.3783646, 0.2689571, 0.2536745, 0.3911419, 0.5213499, 
    0.58079, 0.6880331, 0.7879515, 0.7842073, 0.8093386, 0.8312769, 
    0.9261351, 0.9477644, 0.7625113, 0.6122341, 0.5116653, 0.4521914, 
    0.3856392, 0.3413534, 0.3045535, 0.2150192, 0.276494, 0.1999149, 
    0.09153295, 0.2630827, 0.124362, 0.1720502, 0.2634401, 0.001819134, 
    0.1144331, 0.7544079, 1.060966, 0.6647906, 0.2534304, -0.0399456, 
    -0.2276244, -0.2411661, -0.3993201, -0.4174676, -0.2919965, -0.201582, 
    0.1348271, 0.3605108, 0.6393838, 0.8938107, 1.063602, 1.05942, 1.093844, 
    1.026331, 0.2821581, 0.07564688, -0.04557633, -0.228617,
  -0.1644893, -0.4249873, -0.5465691, -0.2785516, -0.3345091, -0.2648308, 
    -0.05976892, 0.1584604, 0.2906375, 0.4596967, 0.6340134, 0.1933885, 
    -0.1725297, 0.02559841, 0.1567345, -0.04543024, -0.09248352, 0.03782177, 
    0.0003547668, -0.1684127, -0.1413443, -0.02938202, 0.04429954, 
    -0.1183957, -0.2007525, 0.03847277, -0.01076224, 0.0983035, -0.06945372, 
    -0.08250707, -0.04123068, -0.1177931, 0.2015915, 0.3073201, 0.4830852, 
    0.5109172, 0.3726854, 0.3457484, 0.3639288, 0.3528605, 0.3131962, 
    0.3284302, 0.4146442, 0.545536, 0.5064092, 0.531148, 0.6297321, 0.690393, 
    0.8214478, 1.07008, 1.234924, 1.317476, 1.523531, 1.729081, 1.660884, 
    1.512203, 1.214954, 0.9358034, 0.8276148, 0.6757755, 0.5261517, 
    0.4399538, 0.3450642, 0.2789674, 0.3352671, 0.3245738, 0.4992806, 
    0.3974087, 0.05164003, 0.1197392, 0.1665165, 0.1688927, 0.5844526, 
    1.029587, 0.7560511, 0.5072556, 0.3838506, 0.1962042, -0.1608109, 
    -0.5885453, -0.594584, -0.5377312, -0.5714722, -0.4068561, -0.04902697, 
    0.2533813, 0.7174115, 0.9909143, 1.128903, 1.138327, 1.121415, 0.9976687, 
    0.3042774, 0.1524701, 0.1207647, -0.004983902,
  -0.1600947, -0.5319211, -0.7676141, -0.7227409, -0.9305048, -0.6105014, 
    -0.01470101, 0.07901633, 0.27358, 0.3427045, 0.1993945, -0.116442, 
    -0.09523487, 0.1587853, 0.01475859, -0.2498899, -0.1154172, 0.1795375, 
    -0.03421569, -0.3088087, -0.2319211, 0.03832629, -0.01881889, -0.2749549, 
    -0.2707557, -0.1384639, -0.05330782, 0.06109667, 0.05385351, -0.04896188, 
    -0.01321936, -0.08984685, -0.006611586, 0.3010869, 0.3993621, 0.4438443, 
    0.3863077, 0.3846645, 0.3098273, 0.1999149, 0.2792773, 0.2514939, 
    0.3727179, 0.4813769, 0.4679818, 0.6168261, 0.737627, 0.8793259, 
    1.009356, 1.132484, 1.310234, 1.480173, 1.613214, 1.710267, 1.692884, 
    1.550224, 1.27192, 0.9625769, 0.7200155, 0.5000448, 0.3161421, 0.2086878, 
    0.1536422, 0.2033324, 0.2590623, 0.3217574, 0.5324018, 0.2789025, 
    0.2078251, 0.3880007, 0.1880984, 0.5109012, 0.9694462, 0.7874966, 
    0.4132135, 0.3243294, -0.01668644, -0.3883176, -0.6825881, -0.8984737, 
    -0.9619827, -1.119405, -1.009427, -0.7480989, -0.4656284, 0.05336571, 
    0.6893685, 1.094072, 1.263669, 1.281768, 1.184241, 0.9564257, 0.2989223, 
    -0.1037304, -0.1697133, -0.1450882,
  -0.510469, -0.891963, -0.9296423, -0.7230344, -0.79141, -0.3553586, 
    0.008638799, 0.003951252, 0.2104454, 0.1436648, -0.05058974, 0.01155216, 
    0.1791466, 0.146741, -0.1375852, -0.07573621, 0.03144151, -0.06269914, 
    0.08723584, 0.1559695, 0.3343224, 0.5878706, 0.2495404, -0.2738971, 
    0.06186163, 0.5748985, -0.005488753, -0.2916216, 0.1578419, 0.167347, 
    0.2225063, 0.2592087, 0.3268191, 0.641696, 0.6179328, 0.6128058, 
    0.4713998, 0.2522264, 0.1807094, 0.201445, 0.3779421, 0.4510703, 
    0.5665978, 0.6154097, 0.7616175, 0.9786096, 1.032011, 1.17109, 1.155563, 
    1.183997, 1.37109, 1.48831, 1.547262, 1.579358, 1.600875, 1.426315, 
    1.090215, 0.796139, 0.5764773, 0.3722134, 0.1350548, 0.003658533, 
    -0.01416373, 0.1236455, 0.3436648, 0.3562299, 0.2611615, 0.2767868, 
    0.3828738, 0.1784793, -0.03489959, 0.4158003, 0.7022586, 0.30986, 
    0.07221299, -0.08745503, -0.5230019, -0.7473183, -0.9687863, -1.160534, 
    -1.20474, -1.311316, -1.235046, -1.106709, -0.7289588, -0.1321814, 
    0.4349897, 0.8940067, 1.003968, 0.9568813, 0.8337209, 0.5958462, 
    0.3239386, -0.1537304, -0.3752964, -0.3409863,
  -0.707621, -0.8784381, -0.870593, -0.8608106, -0.7351923, -0.576045, 
    -0.1763382, 0.07149744, 0.01287079, -0.1257362, 0.1171023, 0.1557254, 
    0.05502552, -0.1559771, -0.1796587, 0.1196415, -0.1386105, -0.3406938, 
    0.08437121, 0.1436974, 0.168242, 0.6000776, 0.5417607, -0.2798862, 
    -0.1112175, 0.1221476, -0.6644735, -0.01932341, 0.5761359, -0.03906631, 
    0.06173122, 0.2589643, 0.2814741, 0.5366986, 0.5342247, 0.5124962, 
    0.5502079, 0.4297162, 0.2754682, 0.1868941, 0.1792444, 0.2399378, 
    0.5020635, 0.7720828, 1.087269, 1.286813, 1.395277, 1.613554, 1.671546, 
    1.728365, 1.637366, 1.399931, 1.351331, 1.233411, 1.05776, 0.8519983, 
    0.5195764, 0.2727827, 0.04486927, -0.1699419, -0.3125038, -0.3287798, 
    -0.2206418, 0.04386014, 0.2871056, 0.149394, 0.1205206, 0.4632612, 
    0.4522914, 0.2129359, 0.135478, 0.3094851, 0.3254519, 0.09835234, 
    -0.05688855, -0.364587, -0.795821, -1.120544, -1.495202, -1.715238, 
    -1.691703, -1.582816, -1.352168, -1.080423, -0.7139031, -0.3037307, 
    0.1111455, 0.4225389, 0.4603804, 0.5080854, 0.3971154, 0.05732036, 
    -0.09588599, -0.200785, -0.2335325, -0.3518104,
  -0.9321001, -0.9092485, -0.7259796, -0.4227407, -0.3284211, -0.3324738, 
    -0.01958358, 0.1465297, -0.1811397, -0.2317259, 0.05974555, -0.01746795, 
    -0.1680702, -0.1273636, 0.06542587, 0.06238228, -0.118591, -0.02995175, 
    0.1746382, 0.1954226, 0.07823515, 0.2077434, 0.309746, 0.3989873, 
    0.04298162, -0.183727, -0.1625032, 0.3913537, 0.4637169, 0.01314726, 
    0.002291143, 0.2630821, 0.01348901, -0.0343788, -0.3104204, -0.4823443, 
    -0.1633013, -0.06779325, -0.332474, -0.2282097, 0.04062128, 0.1205368, 
    0.2380981, 0.4252238, 0.625257, 0.7744918, 0.9227991, 1.124866, 1.224703, 
    1.388684, 1.474019, 1.33888, 1.131067, 0.8677692, 0.6439579, 0.2942836, 
    -0.09212565, -0.1972041, -0.3680861, -0.5727084, -0.6487339, -0.6530306, 
    -0.5105994, -0.2426307, -0.1074908, -0.153389, -0.06888402, 0.06483996, 
    0.01822567, 0.03933573, 0.07602179, 0.1714482, 0.1877731, -0.009281158, 
    -0.2331907, -0.3745152, -0.6186562, -0.9484408, -1.209069, -1.272008, 
    -1.346032, -1.353193, -1.090172, -0.8379917, -0.6479197, -0.3821652, 
    -0.1503291, -0.08151412, -0.08805728, -0.09263051, -0.2105019, 
    -0.3223345, -0.3864295, -0.4591835, -0.6368853, -0.7367063,
  -1.179153, -1.201794, -0.7730179, -0.2795119, -0.1183954, -0.03768277, 
    0.03186472, -0.08143283, -0.2583371, -0.05262423, 0.0766401, -0.1314166, 
    -0.142061, 0.02078092, 0.1125288, 0.07203382, 0.256409, 0.2973107, 
    0.05474877, 0.3623823, 0.4140263, -0.05176127, -0.03148165, 0.01179635, 
    0.03549427, 0.2048302, 0.2360639, 0.003251433, -0.03200248, 0.001233339, 
    -0.03268576, -0.1106972, -0.2485227, -0.2128131, -0.2985058, -0.6045117, 
    -0.5913444, -0.4475946, -0.5890007, -0.4275427, -0.19906, -0.1473503, 
    -0.08795929, 0.07079697, 0.2238083, 0.2601519, 0.2695274, 0.3757777, 
    0.4628539, 0.4643354, 0.4292121, 0.3469033, 0.146204, -0.1376996, 
    -0.3801794, -0.7165241, -0.8572626, -0.7634478, -0.972497, -1.14237, 
    -1.014733, -0.8871942, -0.6179068, -0.2732134, -0.2782916, -0.3335162, 
    -0.1249551, -0.03763366, -0.02684307, -0.0443716, 0.05697894, 0.02375984, 
    0.02537107, -0.1362011, -0.2979038, -0.3898146, -0.5841506, -0.829267, 
    -0.8401079, -0.7437863, -0.7281775, -0.6768265, -0.5315952, -0.3699093, 
    -0.150557, 0.05785704, 0.005415916, -0.1332068, -0.199857, -0.342598, 
    -0.5208044, -0.6013057, -0.7578324, -0.9028845, -0.8078977, -0.9306515,
  -0.9418159, -0.8580923, -0.5164096, -0.2689328, -0.2765988, -0.1534055, 
    0.1155236, 0.05165625, 0.03632426, 0.2574506, 0.2619591, 0.2281214, 
    0.1126755, 0.2586713, 0.5228641, 0.6006798, 0.5120405, 0.3136029, 
    0.2013634, 0.2930789, 0.226396, -0.1682981, -0.2286171, -0.1752805, 
    -0.2604856, 0.03067648, 0.2167447, -0.4010289, -0.2128779, -0.03374362, 
    -0.4730015, -0.6218297, -0.5257845, -0.5474155, -0.276794, -0.394274, 
    -0.6109085, -0.5621128, -0.402071, -0.5077348, -0.5073929, -0.3225627, 
    -0.06016016, 0.1175747, 0.22402, 0.2238407, 0.1567345, 0.110445, 
    0.04117393, -0.1715212, -0.4408565, -0.6118364, -0.715971, -0.809721, 
    -0.9940147, -1.223572, -1.318981, -1.342224, -1.394876, -1.164196, 
    -0.8430209, -0.7755079, -0.6225295, -0.2638221, -0.1879107, -0.08074903, 
    -0.1139522, -0.4061885, -0.1996946, -0.02560568, -0.02653337, -0.1466997, 
    -0.07897425, -0.1508007, -0.1887727, -0.2511754, -0.4157748, -0.542695, 
    -0.4680204, -0.3918982, -0.2505894, -0.1071324, 0.03160429, 0.2739711, 
    0.4910774, 0.4825811, 0.3716593, 0.2751269, 0.09483719, -0.2675977, 
    -0.6488314, -1.029512, -1.352851, -1.345446, -1.042045, -0.9102247,
  -0.6781447, -0.4857296, -0.1469928, 0.1906862, 0.1118451, 0.07273412, 
    0.2406378, 0.1722298, 0.1992643, 0.2769008, 0.3336716, 0.4828255, 
    0.6358202, 0.7707156, 1.030774, 0.6849409, 0.2485313, 0.3031375, 
    0.5004031, 0.4651492, 0.2414676, 0.09823841, 0.02550077, -0.03849663, 
    -0.0824745, -0.001794145, -0.0725621, -0.34499, -0.2237988, -0.3071809, 
    -0.6679389, -0.5799675, -0.6186557, -0.5815787, -0.3299348, -0.07220411, 
    -0.1570511, -0.410274, -0.2729201, -0.130928, 0.06246328, 0.3114381, 
    0.4478474, 0.4441042, 0.3729129, 0.3130817, 0.3588667, 0.4050422, 
    0.2603641, -0.03574562, -0.2901893, -0.5264688, -0.7440634, -0.8453979, 
    -0.83184, -0.8919148, -1.092777, -1.293623, -1.308761, -1.124402, 
    -0.9547563, -0.8453975, -0.5926468, -0.136218, 0.08053005, 0.2997038, 
    0.1033978, -0.3873572, -0.3155804, -0.1980176, -0.1062536, 0.02555013, 
    0.1363084, 0.005074739, -0.1304234, -0.1368202, -0.1884966, -0.1779492, 
    -0.1559603, 0.02411771, 0.346611, 0.4537239, 0.4901977, 0.6895633, 
    0.7629027, 0.558557, 0.3794556, 0.1286907, -0.2664256, -0.5807981, 
    -0.7974806, -1.051126, -1.209964, -1.139831, -1.040937, -0.8707228,
  -0.2346225, -0.1167514, 0.04236269, 0.1345668, 0.103838, -0.0009796619, 
    0.1281703, 0.3200326, 0.5636196, 0.6041306, 0.550094, 0.628219, 
    0.7571416, 0.7184533, 0.531409, 0.2121219, 0.04158145, 0.08108342, 
    0.0634239, 0.007011056, 0.09202099, 0.1683719, 0.1147586, -0.06074597, 
    -0.04603195, -0.2411487, -0.344974, -0.4808307, -0.3177443, -0.4131382, 
    -0.5233264, -0.4503126, -0.4793327, -0.3627148, -0.04665041, 0.2376428, 
    0.2195604, 0.2231898, 0.2351203, 0.5983524, 0.9287076, 0.9807577, 
    0.8033166, 0.6210575, 0.4949999, 0.4409795, 0.5521126, 0.7243943, 
    0.6446414, 0.292623, -0.07002354, -0.3606968, -0.6279821, -0.8425493, 
    -0.9824252, -1.07917, -1.166507, -1.16086, -1.126273, -1.119617, 
    -1.054414, -0.7700883, -0.1973671, -0.09266335, 0.1893679, 0.1428022, 
    -0.1400752, -0.4390011, -0.2817254, -0.06803727, 0.1238735, 0.2456344, 
    0.3047652, 0.2270309, 0.1228155, 0.1053673, 0.1096641, 0.0370568, 
    0.09516251, 0.2791957, 0.4811332, 0.5259569, 0.7902958, 1.022051, 
    0.9852335, 0.7617805, 0.515296, 0.09713197, -0.4821811, -0.7860057, 
    -0.8568711, -0.8887889, -0.7561722, -0.4903026, -0.3678098, -0.3536,
  0.06726527, 0.4103966, 0.5320446, 0.2874641, 0.06630492, 0.1217906, 
    0.2887988, 0.4428353, 0.5470018, 0.5658982, 0.5382775, 0.4871707, 
    0.3990847, 0.2930952, 0.09690374, -0.1418495, -0.2845249, -0.2342155, 
    -0.2037797, -0.1798532, -0.05594444, 0.05650687, -0.01476598, 
    -0.01701164, -0.06333351, -0.183239, -0.2733271, -0.2596714, -0.407295, 
    -0.4977899, -0.5329297, -0.3665395, -0.08976579, 0.182972, 0.4003222, 
    0.4379365, 0.2900517, 0.3156052, 0.4558554, 0.6097941, 1.068779, 
    1.190279, 0.8656049, 0.832516, 0.9998823, 1.219869, 1.226201, 0.9672814, 
    0.5120893, -0.0123899, -0.3510942, -0.4609249, -0.5129271, -0.6092157, 
    -0.7947624, -1.039635, -1.192386, -1.124841, -0.8682816, -0.5759964, 
    -0.3414751, -0.09266305, -0.1111529, 0.0774539, 0.01018524, -0.06774449, 
    -0.2784705, -0.1543982, 0.1173308, 0.3099734, 0.4184046, 0.5735475, 
    0.8326788, 1.012823, 0.9937959, 0.9492478, 0.3680139, 0.18053, 0.3100388, 
    0.6787562, 1.227193, 1.347588, 1.641223, 1.625029, 1.267754, 0.882988, 
    0.5833299, 0.2428348, -0.03615236, -0.01120114, 0.07724237, 0.0157032, 
    -0.03698254, 0.0187304, -0.03354859, -0.09002614,
  0.6404755, 0.8396935, 0.7886196, 0.4526492, 0.4241663, 0.6653616, 
    0.8437628, 0.7396612, 0.5830366, 0.515849, 0.4951948, 0.3268353, 
    0.1715782, 0.1606733, 0.1087364, -0.05649799, -0.2019569, -0.2433953, 
    -0.216068, -0.2643263, -0.369616, -0.4629266, -0.4967971, -0.4430535, 
    -0.3844597, -0.3713089, -0.3122268, -0.356221, -0.2884802, -0.2483271, 
    -0.2066927, -0.18293, -0.07799816, 0.04721332, 0.2295539, 0.2725875, 
    0.3442669, 0.4310837, 0.4523566, 0.5760866, 0.8552215, 0.7714, 0.3281053, 
    0.3547325, 0.585885, 0.8601038, 0.8630502, 0.5586555, 0.1505823, 
    -0.1054398, -0.1300491, -0.07591534, -0.1067908, -0.224304, -0.3916705, 
    -0.6321978, -0.7656614, -0.6746783, -0.3831583, -0.04134464, -0.07720041, 
    0.04846656, 0.199101, 0.1704555, 0.1294398, 0.1268356, 0.1665814, 
    0.2978967, 0.4173139, 0.465019, 0.5903119, 0.9738573, 1.559876, 1.500468, 
    1.176624, 0.873157, 0.5163862, 0.7859502, 1.180026, 1.454212, 1.651412, 
    1.490345, 1.399264, 1.187627, 0.9309369, 0.7616501, 0.6958137, 0.5659469, 
    0.4789516, 0.5863736, 0.763359, 0.8032681, 0.7207813, 0.6620083, 
    0.5814908, 0.4878547,
  0.8182257, 0.7968389, 0.4596316, 0.3351687, 0.3541143, 0.5239062, 
    0.5892705, 0.6123823, 0.4800906, 0.4047, 0.3735639, 0.287366, 0.1523237, 
    0.05858997, -0.03429739, -0.1260292, -0.2344114, -0.3451372, -0.3403684, 
    -0.375964, -0.3827676, -0.3599321, -0.3614784, -0.3598671, -0.373067, 
    -0.3779659, -0.2848183, -0.1411494, -0.06546581, -0.09022141, -0.1434603, 
    -0.07899141, 0.003235817, 0.1003056, 0.09547162, 0.05014288, 0.04285085, 
    0.03503853, -0.05998087, -0.1232617, -0.1484897, -0.01932311, 
    -0.03812194, -0.08301139, -0.1598505, -0.1341341, -0.1370316, -0.1036496, 
    -0.1842327, -0.195756, -0.2551794, -0.3696001, -0.4654169, -0.6244175, 
    -0.6847038, -0.5669305, -0.4120965, -0.1042025, 0.05800462, 0.157874, 
    0.1714154, 0.1737104, 0.2215295, 0.2297653, 0.2106733, 0.3011844, 
    0.4074994, 0.4538862, 0.5158002, 0.6345503, 0.9421186, 1.268958, 
    1.063391, 0.5368777, 0.1103804, 0.1158978, 0.6652793, 1.193079, 1.277014, 
    0.9305627, 0.4157351, -0.1373248, -0.2349485, -0.1592973, 0.1614547, 
    0.8303999, 1.333753, 1.547652, 1.517607, 1.371155, 1.190865, 1.082076, 
    1.026835, 1.007418, 0.936129, 0.8557092,
  0.3029587, 0.3558885, 0.456686, 0.5277796, 0.6034795, 0.6648074, 0.7809369, 
    0.5290978, 0.396627, 0.2616174, 0.2238894, 0.1756473, 0.09913355, 
    -0.02423882, -0.136039, -0.1887896, -0.1821327, -0.2295122, -0.2679888, 
    -0.3146032, -0.3338742, -0.3259967, -0.2877316, -0.2712766, -0.2810585, 
    -0.2692746, -0.2185911, -0.2011428, -0.1931512, -0.08730817, -0.03180695, 
    0.02022731, 0.199394, 0.2466108, 0.1355431, -0.02751029, -0.1696815, 
    -0.1344928, -0.08017956, -0.03307676, -0.1009967, -0.0755409, 
    -0.08392304, -0.2745481, -0.4524449, -0.5178256, -0.4411654, -0.3592806, 
    -0.3827834, -0.6368198, -0.9417517, -1.470056, -0.9756219, -0.6385291, 
    -0.2777214, -0.08585954, 0.04276991, 0.08601511, 0.1195275, 0.1708133, 
    0.1896447, 0.242965, 0.3110802, 0.3449669, 0.3613406, 0.3979942, 
    0.4918907, 0.6027957, 0.705465, 0.7727501, 0.8104128, 0.798808, 
    0.6393842, 0.4708621, 0.2279747, 0.3331342, 0.5645633, 0.6409792, 
    0.3437136, -0.09547901, -0.4416542, -0.5601762, -0.3555858, -0.06950188, 
    0.117981, 0.2856739, 0.5745244, 1.281247, 1.69609, 1.821498, 1.678382, 
    1.184615, 1.124182, 0.8247684, 0.5544395, 0.3649865,
  0.1166792, 0.1462853, 0.1961225, 0.2939415, 0.4283816, 0.5382124, 0.528935, 
    0.4235476, 0.28914, 0.2235639, 0.2324343, 0.2557253, 0.3283979, 
    0.3580855, 0.1543745, 0.1240848, 0.0872196, -0.004642487, -0.1075233, 
    -0.1743528, -0.2235552, -0.226078, -0.2437699, -0.269242, -0.2283567, 
    -0.1746294, -0.1134474, -0.02340865, 0.07716107, 0.2140429, 0.3055954, 
    0.3929648, 0.4192507, 0.3264447, 0.2535443, 0.1870568, 0.1588504, 
    0.1872361, 0.3697067, 0.4680303, 0.4889777, 0.4174769, 0.3255007, 
    0.1549441, 0.03472928, 0.01365182, 0.008052856, -0.05421931, -0.2542193, 
    -0.4462928, -0.891052, -1.300671, -1.299417, -0.5371616, -0.1355829, 
    0.002356768, 0.06615853, 0.02561462, 0.09441352, 0.04208601, 0.09115827, 
    0.1986126, 0.2126915, 0.3124473, 0.3345664, 0.3817996, 0.4801232, 
    0.6435672, 0.7280886, 0.8049441, 0.6934858, 0.6791466, 0.6162235, 
    0.5887821, 0.5644493, 0.6443972, 0.5147587, 0.3137657, 0.158183, 
    -0.08533883, -0.08867568, -0.356693, 0.009908915, -0.172709, -0.3819373, 
    -0.6050652, -0.6079465, -0.4499875, -0.3207232, -0.2388548, -0.3906937, 
    -0.4952835, -0.3749875, -0.21405, -0.07283902, 0.05427682,
  -0.0167681, 0.177047, 0.3899213, 0.6129682, 0.7815557, 0.8545049, 
    0.8211387, 0.6944948, 0.5360799, 0.4399211, 0.456539, 0.5458781, 
    0.5863245, 0.4318813, 0.3374475, 0.2507285, 0.03222275, -0.06701225, 
    -0.1080604, -0.140287, -0.08428113, 0.009794394, 0.09708281, 0.1559206, 
    0.2201133, 0.2977993, 0.4273565, 0.5423956, 0.6570606, 0.801559, 
    0.7777635, 0.7996711, 0.774557, 0.7249639, 0.6574835, 0.5904751, 
    0.582158, 0.5617315, 0.5607874, 0.5590293, 0.4968874, 0.4347618, 
    0.3682253, 0.3038862, 0.2704389, 0.283118, 0.3100223, 0.3253543, 
    0.2906212, 0.2401167, 0.1753868, 0.133281, 0.1286099, 0.1644657, 
    0.2063279, 0.2382779, 0.2199017, 0.2019167, 0.2057904, 0.240556, 
    0.3002242, 0.4373176, 0.6137825, 0.4306605, 0.4849409, 0.5894005, 
    0.6285443, 0.6494265, 0.6137169, 0.6104943, 0.49373, 0.4182091, 
    0.3230919, 0.2857547, 0.1999799, 0.07141548, 0.002942145, -0.09653711, 
    -0.139522, -0.2956255, -0.3798865, -0.2419956, -0.03566432, -0.1180205, 
    -0.1229039, -0.07332736, -0.02588248, 0.07416582, 0.1680946, 0.07543588, 
    -0.170202, -0.2688679, -0.3675982, -0.5202512, -0.4528684, -0.2085162,
  -0.1052448, 0.345602, 0.8265915, 1.212757, 1.464466, 1.385657, 0.8800097, 
    0.414515, 0.2379196, 0.1062138, -0.002183914, -0.02134109, 0.008688211, 
    0.07397103, 0.1030074, 0.05097306, -0.004805207, -0.009150803, 
    0.01243109, 0.05370712, 0.1277956, 0.2408328, 0.3581831, 0.4908491, 
    0.574687, 0.6195111, 0.6777631, 0.6785769, 0.6940392, 0.6823041, 
    0.641256, 0.5584923, 0.504521, 0.4486453, 0.4102339, 0.3764285, 
    0.3289676, 0.3147098, 0.3123497, 0.3130659, 0.3313276, 0.3352664, 
    0.3355919, 0.3140424, 0.2901655, 0.2849897, 0.2986616, 0.3283817, 
    0.3510866, 0.3827273, 0.3841921, 0.3691857, 0.347213, 0.3257287, 
    0.3144655, 0.282939, 0.2495731, 0.2511355, 0.2916791, 0.3566856, 
    0.4063927, 0.4679487, 0.5570111, 0.6795046, 0.7689578, 0.593258, 
    0.5659468, 0.5507938, 0.5316368, 0.479993, 0.4373823, 0.3857872, 0.35234, 
    0.251933, 0.2467248, 0.1844689, 0.1414348, -0.08183956, 0.09345388, 
    0.1090784, 0.1731739, 0.1062469, -0.04894567, -0.06142926, 0.01378202, 
    0.1019821, 0.1464489, 0.2008591, 0.227356, 0.1907191, 0.06519818, 
    -0.1364943, -0.2429399, -0.3018593, -0.2640174, -0.2005572,
  -0.05268919, 0.06729758, 0.2530726, 0.3654263, 0.2306607, 0.2496221, 
    0.3026005, 0.3164837, 0.2496055, 0.1902468, 0.1332645, 0.101168, 
    0.09708279, 0.1205691, 0.1813763, 0.2577599, 0.3287234, 0.3850548, 
    0.4208946, 0.4546512, 0.4798465, 0.5060508, 0.549101, 0.5966271, 
    0.5919232, 0.508297, 0.4739057, 0.4186648, 0.365491, 0.3432254, 
    0.3575483, 0.3288862, 0.3074832, 0.3040164, 0.3008914, 0.2898888, 
    0.281702, 0.2701622, 0.2749962, 0.2907352, 0.3140587, 0.3291629, 
    0.3449995, 0.3383425, 0.327226, 0.3006147, 0.2597944, 0.2176394, 
    0.1724083, 0.1436811, 0.1366336, 0.1562462, 0.1876752, 0.2162885, 
    0.2503543, 0.2902467, 0.3553835, 0.4294884, 0.5010542, 0.5619428, 
    0.6127567, 0.6253217, 0.6077273, 0.5645958, 0.5241823, 0.4798463, 
    0.4629192, 0.4456667, 0.4088014, 0.3837852, 0.3780724, 0.2765262, 
    0.2423627, 0.1088341, 0.06518197, -0.03502953, -0.1312536, -0.2077022, 
    -0.3669631, -0.5054561, -0.5360227, -0.5864133, -0.5604693, -0.5214716, 
    -0.50002, -0.4508336, -0.3574581, -0.2107782, -0.06709337, 0.05193377, 
    0.09037757, 0.008785486, -0.008239508, -0.08970106, -0.1303749, -0.1132688,
  -0.2847206, -0.3321328, -0.3552772, -0.3640825, -0.3431841, -0.3193398, 
    -0.2886269, -0.2444537, -0.1844602, -0.1241087, -0.06784236, -0.01654029, 
    0.03002548, 0.06739521, 0.09848261, 0.1211876, 0.1416628, 0.1707156, 
    0.2063764, 0.2488568, 0.290312, 0.3260379, 0.3788048, 0.4200971, 
    0.464547, 0.4845991, 0.5124475, 0.5345502, 0.590019, 0.6227013, 
    0.6551557, 0.6779584, 0.6926231, 0.6924279, 0.682532, 0.6593875, 
    0.619202, 0.5749148, 0.5357872, 0.4897586, 0.4414839, 0.3919884, 
    0.3456343, 0.3066369, 0.2774376, 0.2595014, 0.2441694, 0.2312299, 
    0.2266727, 0.2165327, 0.2169884, 0.2155887, 0.21095, 0.2165652, 
    0.2339806, 0.2428999, 0.2476199, 0.2613894, 0.2699832, 0.2869591, 
    0.283769, 0.2837039, 0.2834923, 0.2828413, 0.2802534, 0.2725548, 
    0.2637006, 0.2566857, 0.2473432, 0.2313927, 0.2042116, 0.1681765, 
    0.1103966, 0.0431928, 0.04700142, -0.01717499, -0.05934624, -0.07975638, 
    -0.1097043, -0.0931353, -0.003926516, -0.04549527, 0.05154264, 
    0.06420553, 0.09532523, 0.1811976, 0.2227666, 0.2330368, 0.226917, 
    0.1763797, 0.104586, 0.02047139, -0.04655331, -0.1202349, -0.1860064, 
    -0.2408241,
  -0.4392291, -0.4318072, -0.4182492, -0.4000689, -0.3784381, -0.3510129, 
    -0.3229856, -0.2873899, -0.2521523, -0.2097043, -0.1658567, -0.1304073, 
    -0.09381896, -0.0538612, -0.01680058, 0.02069944, 0.05585569, 0.0879032, 
    0.1214318, 0.1546023, 0.1870242, 0.2202273, 0.2572716, 0.2935346, 
    0.3269982, 0.3617313, 0.3988081, 0.4268517, 0.4583133, 0.4882612, 
    0.5125288, 0.5334598, 0.5511193, 0.5693159, 0.5791954, 0.585299, 
    0.5935834, 0.5871869, 0.5805789, 0.5715131, 0.5664187, 0.5499799, 
    0.5330853, 0.5075808, 0.4851362, 0.4725385, 0.4537885, 0.4280398, 
    0.4002728, 0.3787397, 0.3574994, 0.33206, 0.3010216, 0.2724246, 
    0.2481245, 0.2260378, 0.200517, 0.1753217, 0.1515913, 0.1328738, 
    0.1135053, 0.1028445, 0.09786406, 0.0961225, 0.08349231, 0.06819284, 
    0.064547, 0.06202421, 0.06143827, 0.06350533, 0.06171497, 0.04713164, 
    0.03280872, 0.02286405, 0.005969524, -0.02021863, -0.0478879, -0.0721392, 
    -0.0912961, -0.1140988, -0.143591, -0.1704953, -0.2021034, -0.2319048, 
    -0.2589393, -0.284395, -0.3092323, -0.3284543, -0.3538287, -0.3752805, 
    -0.3926958, -0.4069048, -0.4187863, -0.4290728, -0.4416216, -0.4413776 ;
}
