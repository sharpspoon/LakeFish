netcdf CGMR_SRA1B_1_rsds-change_2070-2099 {
dimensions:
	time = 12 ;
	latitude = 48 ;
	longitude = 96 ;
	bounds = 2 ;
data:
 surface_downwelling_shortwave_flux_in_air_anomaly =
  -9.644806, -9.935394, -10.29141, -10.85913, -11.38229, -11.89532, 
    -12.34116, -12.82733, -13.43463, -14.00052, -14.37476, -14.6539, 
    -15.00208, -15.52216, -16.00156, -16.60391, -17.24557, -17.77994, 
    -18.1893, -18.59766, -19.14871, -19.48596, -19.81042, -19.97916, 
    -20.19141, -20.09195, -19.76434, -19.53983, -19.12604, -18.61093, 
    -18.11563, -17.8349, -17.59634, -17.26666, -16.91928, -16.52396, 
    -16.06042, -15.51981, -14.8414, -14.39868, -14.07007, -13.72345, 
    -13.63101, -13.48019, -13.47656, -13.82867, -14.30365, -14.9646, 
    -15.61328, -16.31589, -17.01016, -17.44009, -17.4711, -17.2854, 
    -16.61249, -15.72916, -14.67761, -13.74481, -12.76901, -11.86981, 
    -11.15729, -10.72943, -10.45883, -10.13724, -9.764862, -9.320587, 
    -9.048187, -8.959137, -8.573944, -8.266663, -8.179443, -8.176819, 
    -8.350769, -8.274475, -8.363281, -8.598175, -8.973175, -9.228638, 
    -9.429932, -9.584381, -9.689606, -9.635956, -9.722382, -9.969543, 
    -10.29556, -10.41483, -10.61746, -10.69507, -10.51587, -10.3815, 
    -10.12292, -9.746094, -9.299225, -9.331512, -9.405975, -9.458313,
  -22.90729, -22.71588, -21.79086, -19.95859, -18.04477, -16.97241, 
    -16.12344, -15.50961, -14.71146, -13.94217, -13.52216, -13.96353, 
    -14.90286, -16.29611, -18.0018, -19.75494, -21.62448, -23.46432, 
    -25.26303, -26.73386, -28.00937, -28.90808, -29.19272, -28.64142, 
    -27.33829, -25.43933, -23.17917, -21.28568, -18.90753, -17.27762, 
    -16.05783, -15.7229, -15.40155, -15.16171, -14.73749, -13.66223, 
    -12.79504, -12.38931, -12.14948, -11.33359, -10.22528, -9.515106, 
    -9.344788, -9.139832, -8.773956, -8.098694, -7.275024, -6.710144, 
    -6.692444, -7.333069, -7.981232, -8.610931, -9.650787, -11.85834, 
    -13.21457, -13.78699, -13.67682, -12.73282, -11.36432, -10.47162, 
    -10.28464, -9.952332, -8.594818, -7.264832, -6.0401, -5.448425, 
    -4.881256, -3.809631, -2.061707, -0.4315186, 1.654175, 3.5961, 4.496094, 
    6.048462, 7.326843, 7.300781, 6.149994, 4.388031, 2.62265, 1.706512, 
    1.06485, 0.6296997, 0.2049561, -0.5739441, -1.956238, -4.247131, 
    -6.880493, -8.550507, -10.91199, -13.50937, -15.90729, -17.60522, 
    -19.65704, -20.77838, -21.78671, -22.49948,
  -14.39685, -14.47266, -15.71329, -16.53568, -17.46222, -18.82422, 
    -19.49347, -18.44193, -17.58566, -17.48621, -17.63904, -16.98621, 
    -16.76718, -17.10129, -16.86691, -16.61145, -16.20389, -16.47733, 
    -17.81119, -18.69064, -20.92447, -23.0354, -24.98047, -26.10391, 
    -25.84244, -24.15912, -21.38699, -19.72266, -18.65079, -17.92889, 
    -18.23749, -18.8396, -19.85519, -20.65182, -21.13492, -22.03958, 
    -23.96198, -26.10938, -25.90573, -23.33228, -18.79971, -13.75443, 
    -9.210938, -5.841125, -2.960693, -2.158081, -1.872894, -1.3909, 
    -0.8442688, -0.8518372, -1.783569, -4.035675, -6.463013, -6.957275, 
    -5.301819, -3.245056, -0.9382629, 1.198181, 1.938782, 0.9505157, 
    -1.768738, -5.304169, -6.683594, -7.583328, -8.825516, -11.37006, 
    -13.56693, -13.87082, -13.09608, -10.12082, -5.205475, 0.6484375, 6.0271, 
    9.535431, 11.82135, 12.52344, 13.13959, 12.82498, 12.14322, 10.97812, 
    8.880981, 5.817993, 2.733856, -0.2466125, -3.371094, -5.558319, 
    -10.17499, -14.29871, -17.53802, -18.96643, -19.15469, -19.36978, 
    -19.56589, -18.68982, -17.70651, -15.74478,
  -10.66824, -8.791168, -5.79245, -2.336212, -1.834869, -3.868256, -6.217712, 
    -6.857056, -6.770569, -7.52005, -8.15625, -7.941681, -6.235931, 
    -5.243744, -5.987488, -7.366669, -7.454407, -8.521637, -9.7901, 
    -12.06143, -13.36743, -13.83722, -14.43854, -12.67032, -12.75156, 
    -14.0849, -15.17029, -14.95599, -14.8526, -15.07162, -14.96222, 
    -14.28516, -12.63437, -11.11224, -9.666931, -11.37137, -14.99008, 
    -19.84766, -22.87134, -23.66226, -21.52005, -15.44687, -7.929962, 
    -3.31015, -1.583588, -1.63385, -6.024231, -8.857574, -12.98517, 
    -9.633591, -8.845566, -12.70105, -15.21512, -12.08855, -6.076813, 
    -0.1635437, 7.950256, 10.92265, 8.381516, 3.828644, -1.135941, -5.294525, 
    -6.797409, -6.125519, -5.601563, -3.288544, 0.2049561, 2.249756, 
    6.058594, 7.126038, 8.277863, 8.838531, 6.384369, 5.036194, 6.137756, 
    6.654449, 5.762238, 4.240112, 5.003387, 4.453888, -0.9440002, -2.821106, 
    -7.431244, -12.78438, -16.91145, -20.60728, -23.25208, -26.31537, 
    -27.80026, -28.17474, -27.94296, -27.40677, -24.43958, -22.68515, 
    -20.22421, -15.30783,
  -2.1409, 1.280975, 2.476563, 3.180206, -1.395569, -6.5224, -8.985687, 
    -10.69818, -11.43777, -12.7659, -13.40964, -16.03125, -16.92267, 
    -13.21484, -10.84195, -7.863281, -5.438782, -7.539063, -9.532288, 
    -10.70886, -9.10965, -5.836456, -5.390106, -4.474762, -1.555725, 
    0.430481, -0.5619812, -2.5802, -4.231506, -6.525787, -7.784637, 
    -9.532288, -11.14948, -12.35519, -10.79321, -7.972107, -5.401031, 
    -7.2789, -9.836212, -11.58487, -15.42941, -16.19998, -15.9104, -13.57605, 
    -10.60522, -9.715363, -14.65128, -13.71225, -8.948181, -0.2005157, 
    5.523956, 9.17395, 7.550522, 1.329681, -3.073441, -6.723434, -12.00261, 
    -14.45963, -17.05676, -17.57266, -16.76122, -16.28618, -15.50807, 
    -14.9922, -14.92293, -14.05467, -10.82343, -4.748688, -1.76355, 
    -0.07003784, 2.652603, -7.358337, -12.65051, -15.33855, -10.0961, 
    -2.923172, -1.539581, -1.206772, -1.085938, -0.6742096, -1.802872, 
    0.1015625, -0.7848816, -2.311707, -3.381256, -6.289856, -9.793488, 
    -12.26772, -17.62994, -25.13748, -32.02267, -26.29636, -26.8508, 
    -21.85025, -15.42578, -8.876831,
  -18.94324, -9.366669, -3.5383, -1.934906, -4.431244, -5.851318, -10.66849, 
    -15.08826, -16.49454, -16.0672, -17.22552, -19.70261, -21.22424, 
    -16.95651, -12.58646, -5.795319, -1.039856, 1.058075, 1.122131, 
    -0.8661499, -2.163544, -3.155731, -2.007294, -3.595062, -6.020844, 
    -4.711975, -4.491425, -4.366394, -4.202362, -5.993744, -10.88229, 
    -13.50861, -12.18335, -8.748169, -2.699738, 2.090363, 2.553375, 
    -0.03671265, -0.5596619, -1.815887, -1.476288, -0.04141235, -1.015625, 
    -6.689575, -14.15887, -8.900513, -8.315628, -9.317444, -8.525269, 
    -4.541138, -0.138031, 0.4885406, -1.730728, -6.077087, -4.092438, 
    1.798965, 3.683319, 1.746613, -7.539581, -14.42604, -16.07344, -12.54558, 
    -8.418762, -11.02214, -15.71666, -16.91277, -11.89427, -6.375519, 
    -5.251556, -8.494278, -16.54767, -15.54532, -14.29843, -14.55728, 
    -16.86745, -17.61511, -10.15521, -3.065109, -2.019012, -2.013535, 
    -12.73724, -10.7065, -15.78334, -25.89009, -31.65285, -34.37733, 
    -32.15105, -28.64038, -23.23282, -21.1927, -21.12473, -24.46899, 
    -25.32944, -26.48541, -28.96146, -27.01822,
  -59.65884, -53.24245, -51.01251, -51.19087, -50.27631, -46.40729, 
    -47.98465, -51.12657, -54.51511, -54.09558, -55.19975, -52.21667, 
    -45.73697, -41.64896, -37.95181, -28.17398, -16.79504, -12.77084, 
    -15.63931, -17.47212, -15.95285, -15.16016, -13.93414, -16.08279, 
    -17.85419, -15.68567, -12.91876, -12.64063, -15.92969, -20.42654, 
    -21.7211, -24.14166, -27.21484, -20.4729, -10.62033, -4.792725, 
    -17.56613, -21.86275, -13.91354, -10.05, -9.497406, -6.419006, -1.729675, 
    -0.0223999, -2.305984, 0.5338593, -1.601044, -1.320572, 2.754425, 
    4.002853, 2.277344, -0.7497406, -4.850525, -9.605209, -11.27473, 
    -8.745834, -5.240112, -12.30312, -17.6526, -14.00652, -5.717957, 
    -3.835938, -7.961716, -12.48932, -13.11719, -6.179169, 1.463547, 
    -1.587753, -7.014069, -8.268753, -7.654175, -6.343231, -3.942184, 
    -5.069534, -7.216934, -9.21199, -6.879944, -3.490372, -3.407028, 
    -22.04504, -38.49271, -36.17995, -24.94115, -18.00287, -20.31615, 
    -29.9362, -38.46225, -41.51118, -44.08125, -49.26122, -48.80077, 
    -48.84608, -52.36693, -57.16171, -63.37267, -63.23332,
  -12.67162, -12.42813, -12.14948, -8.469009, -8.621353, -14.66589, 
    -15.16588, -9.983856, -6.630981, -7.047668, -12.28645, -14.37865, 
    -13.40807, -9.807556, -6.897125, -2.556503, 6.68541, 6.541931, 3.768753, 
    3.522919, 5.245834, 3.48645, 0.686203, -0.1591187, -2.1875, -2.479172, 
    -3.27655, -3.923431, -7.382278, -8.568756, -10.76772, -12.68489, 
    -14.56979, -16.27449, -12.46458, -4.403641, -0.9617157, -0.06797791, 
    -1.334122, -1.489334, 0.6838531, 3.484116, 5.141937, 4.476303, 0.828125, 
    -5.067444, -9.109894, -10.40182, -9.627075, -14.74609, -17.06694, 
    -14.2263, -10.28229, -5.070313, -1.337234, -1.120575, -4.597397, 
    -12.20599, -20.47839, -15.46199, -11.10495, -12.94688, -21.40366, 
    -20.05209, -9.008331, -3.619003, -1.512512, -2.575256, -2.709641, 
    -0.0148468, 3.134903, -0.08514404, -0.2268219, 3.123444, -0.1580811, 
    -4.638275, -6.247406, -7.240891, -8.114059, -5.637756, -2.076294, 
    -2.380981, -4.41301, -9.880203, -11.17787, -14.14818, -14.90105, 
    -16.72058, -20.94818, -18.35469, -12.89322, -10.35834, -11.56979, 
    -17.82448, -18.13385, -14.75546,
  -9.6026, -7.289581, -7.316925, -7.21199, -5.413025, -11.95313, -9.863281, 
    -8.206512, -5.698441, -8.473709, -8.12265, -5.388809, -0.8585815, 
    -1.024475, -2.296097, -2.831512, -3.451553, -3.007553, -3.265091, 
    -6.27005, -3.421616, -4.982819, -7.544525, -6.121872, -3.950012, 
    -9.670578, -14.28699, -13.9586, -11.8737, -12.10052, -14.18385, 
    -15.29974, -14.8802, -13.01224, -16.36171, -16.11874, -13.99037, 
    -9.371613, -9.765366, -4.158325, -0.7098999, 0.8716125, -2.219269, 
    -6.579422, -3.205475, -3.053391, -4.540359, -8.966934, -8.272919, 
    -10.23021, -13.00365, -11.38152, -6.246872, -9.208862, -13.00807, 
    -8.437241, -2.891922, -7.56041, -13.33098, -12.55521, -8.408081, 
    -10.60832, -14.11015, -10.39688, -9.887238, -6.04245, -9.058868, 
    -10.58855, -10.2552, -7.449997, -5.267197, -7.033585, -3.901291, 
    0.1856842, 1.823959, -2.143234, -9.636719, -8.870834, -3.895309, -3.3638, 
    -7.121872, -5.184891, -1.463806, -0.3697968, -5.637497, -11.12109, 
    -9.179428, -9.532547, -15.05208, -15.31354, -6.016663, -5.409637, 
    -10.18646, -6.597382, -4.914063, -6.353638,
  -4.624222, 3.848175, -3.61824, -12.12657, -8.00885, -4.401566, -1.000778, 
    -3.754181, -7.634109, -7.228653, -3.220306, -2.566406, -4.976822, 
    -8.324478, -1.334381, 3.110931, 4.025513, 1.727341, 3.13855, 3.143753, 
    6.535934, 5.576294, -2.063797, -1.441147, -2.780731, -8.831512, -11.8573, 
    -9.366409, -9.207031, -12.46381, -8.33255, -9.247925, -8.652603, 
    -11.41353, -8.386444, -2.446091, -2.973694, -9.341919, -6.061981, 
    -0.6622314, -0.3179626, -1.844788, 0.3158875, 0.3674469, -1.246094, 
    -1.397919, -1.238022, -5.689575, -6.723434, -7.553894, -9.260941, 
    -7.146881, -3.953903, -4.252075, -7.137756, -7.571091, -7.483841, 
    -9.738541, -7.970825, -3.349228, -10.52031, -10.46379, -6.209641, 
    -1.566147, 0.5395966, -2.257553, -4.183853, -0.653656, -5.486969, 
    -9.832291, -11.41901, -6.098694, 0.1078033, -0.9898376, -4.509384, 
    -4.508072, -11.5, -13.30626, -11.52187, -8.585159, -7.300781, -11.25861, 
    -7.529175, -5.341919, -6.017441, -11.99348, -10.67682, -15.61458, 
    -22.32005, -14.62837, -7.332291, -11.7901, -10.57631, -2.279434, 
    -3.711456, -9.450256,
  -0.4460907, -5.937759, -6.388794, -3.12735, 4.964844, 2.071365, 0.973175, 
    5.612503, -0.7294312, -2.551559, 5.322128, 7.775772, 3.140106, 2.534119, 
    3.070053, 5.072403, 9.250519, 8.208603, 5.756256, 8.791656, 9.109894, 
    5.9263, 5.047134, 1.4039, 0.9000092, -3.069016, -0.1822968, -0.3213501, 
    -2.121353, -3.795837, -0.1013031, 0.759903, -5.675003, -6.778641, 
    -0.683075, 1.351044, -4.915375, -5.759628, 1.253906, 2.792709, -2.316132, 
    -3.326569, -0.7963562, 4.982544, 4.657028, 1.031769, 4.321884, 3.774475, 
    -0.4507751, 4.921356, 1.505997, -2.056778, 2.537231, 0.9098969, 
    -6.835159, -6.832031, -14.09921, -12.67995, -7.248962, -8.167709, 
    -8.979691, -4.831253, -0.7885437, -2.951569, -4.180481, -4.191666, 
    -5.695572, -5.736206, 1.194519, 0.768219, -1.302078, 0.0690155, 
    -3.445053, -4.9552, -5.611206, -5.280472, 0.8190155, 0.9658813, -2.38205, 
    5.194275, 2.786713, -4.483841, -2.944778, 0.97995, -0.6622314, 0.7338409, 
    2.702347, -2.713272, -5.136978, 0.4051971, -2.288803, -8.160934, 
    -5.879944, -3.725769, -1.350784, -1.000778,
  -0.2890625, -1.978653, -0.08984375, 4.776031, 2.960419, -1.445831, 
    2.999725, 8.924484, 11.67526, 6.659119, 4.0289, 1.980728, 6.291931, 
    7.180725, -0.9755249, 2.421616, 9.954697, 9.894272, 5.626816, 6.145584, 
    5.176834, 4.208069, 6.154938, 6.49791, 0.1619873, 3.552353, 8.26329, 
    5.515625, 2.916931, 1.507034, 3.753647, 5.764069, 2.247925, 2.965897, 
    4.627075, 3.738037, 5.348694, 4.831253, 6.226563, -0.5604248, -1.098969, 
    3.036194, 1.8703, 4.122131, 6.727875, 13.10963, 13.79375, 12.33151, 
    4.696625, 12.08517, 14.48465, 9.072906, 8.811203, 4.636475, 1.934372, 
    0.2151184, 4.070831, 4.435944, -0.1359558, -2.191925, 3.4039, 6.612488, 
    1.509094, -2.530472, -0.4916687, 2.189056, -0.1171875, -0.8388062, 5.681, 
    9.779434, 0.05807495, -0.5489655, 3.500244, 5.166138, 3.787491, 
    -1.009109, -4.0401, 13.94141, 12.80678, 9.927612, 7.563812, 2.808594, 
    1.200806, 2.970856, 5.065094, 3.692688, -0.7861938, -1.122925, 1.019287, 
    2.531525, -4.20105, 0.8622437, 9.397919, 7.540894, 2.894272, 1.6138,
  4.144012, 3.836456, 9.769806, 6.661713, 8.671875, 17.625, 10.90259, 
    8.646851, 11.50391, 13.45544, 9.952606, 5.388, 5.424713, 4.03125, 
    5.231262, 10.66122, 7.139069, 2.634888, 5.048706, 11.92212, 9.692688, 
    7.638794, 5.973419, 5.656494, 4.140625, 9.06485, 11.87659, 10.63565, 
    12.27292, 11.12396, 13.99869, 12.93387, 10.9841, 9.926575, 11.62762, 
    12.03986, 7.476044, 0.4604187, 6.096619, 11.29037, 7.957275, 9.440369, 
    7.988556, 6.154419, 7.084381, 13.91275, 25.32396, 17.46277, 17.43359, 
    15.77267, 16.36771, 12.26068, 9.904175, 6.580719, 12.3367, 10.32187, 
    9.402344, 6.203125, 7.370575, 7.375793, 5.1828, 6.101807, 3.773956, 
    7.52005, 7.338806, 8.286987, 6.765381, 2.902863, 4.71405, 4.492737, 
    5.980469, 2.337494, 0.75, 0.4080811, 3.135406, 3.577362, 8.988556, 
    22.69374, 27.0672, 14.49609, 1.150787, 2.273193, 11.04401, 5.090118, 
    -0.9841003, 1.654419, 4.860168, 4.345306, 3.372406, 0.8392944, -1.262238, 
    -2.040649, 0.2453308, 1.310699, 0.2109375, 0.5078125,
  2.757263, 4.615875, 5.722656, 6.453918, 5.281006, 4.681488, 7.023956, 
    8.534119, 9.724731, 5.729156, 7.761444, 8.413818, 9.344788, 8.945313, 
    12.62344, 11.73047, 9.168762, 6.774994, 10.44376, 9.680725, 5.21875, 
    3.618744, 2.226044, 4.44455, 4.645844, 6.144531, 12.81354, 14.15234, 
    19.25601, 14.76953, 13.52136, 7.9534, 7.528107, 12.66953, 10.43384, 
    8.123962, 5.775513, 3.882538, 25.89218, 37.69583, 23.06693, 14.08698, 
    9.264832, 11.11615, 10.60831, 10.12213, 22.38959, 34.59271, 22.15625, 
    16.38907, 19.21719, 15.45209, 7.519287, 13.9487, 14.28308, 9.410156, 
    4.142181, 2.885162, 10.9711, 12.98489, 8.675537, 7.305206, 5.525787, 
    4.146088, 5.421356, 4.726044, 9.362244, 5.847656, 0.7874756, 3.102081, 
    1.2034, -3.582306, 0.9901123, 2.639313, -0.8997192, 0.9893188, 11.90781, 
    20.00522, 24.47137, 13.54193, 1.616425, 3.083099, 5.394012, -0.754425, 
    3.420837, 1.995575, -5.786194, -3.762512, -3.603119, -2.646332, 1.5672, 
    0.5471497, -1.155212, 3.932556, 3.512238, 2.425537,
  -3.378113, -1.380737, -1.984894, -7.094543, -4.010651, 2.132813, 1.821869, 
    -1.982544, -3.083344, 2.527863, 8.7117, 4.661469, -2.646362, 0.9518127, 
    -7.910156, -2.173676, -2.690613, -2.808075, -1.308594, -0.7307129, 
    1.22995, 7.666138, 3.061432, 4.321869, 1.946075, 3.226318, 5.413269, 
    1.020325, 6.645294, 3.497406, 4.149475, 5.693481, 1.891388, 1.441925, 
    -0.9750061, -1.137482, 7.134125, 12.42578, 15.46069, 18.57214, 9.715607, 
    -0.3640747, 2.072662, 1.626312, 2.064575, 5.89505, 7.464569, 13.13126, 
    10.46512, 9.311981, 11.13983, 7.800781, 9.805206, 8.877594, 4.862518, 
    6.747131, 2.742432, 2.360687, 4.039825, 2.408081, 7.955994, 7.872375, 
    7.794769, -1.144531, 1.836731, -0.2622375, 1.914581, -1.061462, 
    -4.747925, 1.278107, -0.6023254, -2.264832, -0.06668091, -5.729431, 
    -6.75, -0.6841125, 2.438782, 5.427338, 10.06744, -0.1046753, -9.125519, 
    -3.644531, -7.439331, -10.17499, -6.0755, -7.172668, -5.996887, 3.077362, 
    4.717712, 4.272919, 0.8638, -0.2630005, 3.163544, 3.240112, -7.915619, 
    -4.166138,
  -5.792694, -2.411987, -4.294525, 0.3919373, -0.1104126, -0.6138, -4.292175, 
    -12.23749, -18.75235, -13.00443, -2.400787, -6.058319, -10.49585, 
    -6.37265, -2.321594, -2.518738, 2.952362, -2.566132, 0.03125, -2.848694, 
    0.6484375, 0.4067688, -4.360657, -5.342712, -7.505463, -6.333588, 
    -7.166656, -6.430481, 0.01693726, 2.196869, 5.0224, 1.746338, -3.807556, 
    -7.029419, -0.09844971, 2.219543, 3.149994, 3.08725, 2.767456, 3.003906, 
    -2.501556, -7.17865, -10.02084, -7.507263, -9.517456, -6.118469, 
    -8.714325, -5.511719, 1.688568, 4.222931, 1.681488, -1.669006, 0.7791748, 
    0.06222534, -1.135132, -1.353119, -3.727081, -2.068237, 2.764038, 
    4.900513, 2.202087, -0.0552063, 0.6276245, 0.7145996, 1.023438, 
    -3.692963, 0.5177002, 2.289307, 4.489319, -2.11145, -1.395844, -3.005737, 
    -5.019012, -6.414307, -1.053131, -4.75235, -4.453125, -0.8557434, 
    5.387756, -12.82291, -21.87866, -5.250244, -14.39346, -9.215363, -5.9599, 
    -2.479156, 5.628662, 5.720581, 9.3638, 9.666382, 5.322388, -3.766937, 
    -6.041931, -7.505737, -0.336731, -4.4888,
  -4.003662, -6.760681, -4.016144, -7.689331, -4.7388, -8.371613, -12.91199, 
    -19.56613, -16.59663, -6.351318, -14.30103, -7.571075, -11.08905, 
    -5.458588, 2.967987, -0.6760254, -3.73645, -1.390106, -4.295319, 
    -4.96875, -7.599976, -6.695557, -11.44763, -14.2677, -13.18878, 
    -8.645844, -6.722382, 4.204956, 6.7211, -0.5614624, -6.485931, -12.11511, 
    -8.705444, -5.894806, -3.115112, 4.53595, 3.404419, -1.388824, -2.950775, 
    -7.408875, -8.308594, -14.20911, -15.72345, -12.67944, -17.23724, 
    -12.96042, -10.12448, -6.199463, -4.837494, -6.26355, -8.307556, 
    -8.337769, -8.904175, -9.280212, -6.312225, -0.06588745, 1.264343, 
    0.6867371, -2.767975, 1.900513, 0.7067871, 1.551056, 1.290375, 
    -0.3622437, 0.3557434, 0.1893311, -3.654694, -7.173187, -11.04269, 
    -8.112244, -14.16302, -6.057281, -5.497925, -2.354675, -4.360443, 
    -5.587494, -3.075531, -0.6950378, 14.81589, 0.5117188, -8.328888, 
    2.079681, -10.59895, -2.120819, -6.581238, -3.634888, 1.715881, 2.172638, 
    -1.828125, -3.71405, -6.493225, -8.899994, -4.940857, -4.888031, 
    -1.777069, -4.478638,
  -3.046875, -0.09973145, -5.517212, -5.273956, -10.33203, -13.19556, 
    -18.1651, -20.84271, -10.13983, -3.761719, -3.470306, -3.883881, 
    -7.201294, -8.094788, -0.3781433, -1.910919, -1.86615, -1.805725, 
    -9.003387, -6.496887, -9.738525, -6.464569, -9.485413, -5.769806, 
    -9.400269, -0.2098999, 3.728638, 7.172394, 12.19141, 3.073975, -9.705994, 
    -10.18829, -7.663269, -2.855194, 0.6799622, 5.170074, 4.83905, -2.850494, 
    -10.37628, -13.47501, -12.24869, -11.37109, -8.601563, -14.13019, 
    -12.11404, -9.513306, -4.277344, 0.2846375, -4.313568, -7.598694, 
    -12.5065, -13.25912, -7.338806, -9.289307, -3.568237, 0.0385437, 
    -1.635437, -4.262756, -4.840881, -3.158569, -0.317688, -3.183075, 
    -0.0869751, -2.284912, -5.414612, -10.59116, -17.88959, -18.5466, 
    -12.73856, -5.969269, -6.680481, -0.5432434, -0.7325439, -1.627594, 
    1.552063, 6.045563, 2.291931, 1.006256, 27.04739, 8.046097, -8.020569, 
    19.96223, -1.842987, -4.065109, 0.5385437, 11.76068, 8.538544, 2.901306, 
    -6.079956, -13.59766, -16.03723, -13.26849, -7.138, 0.4637756, -2.980194, 
    1.65155,
  -1.33725, -1.792175, -8.977325, -4.788025, -15.78177, -19.70105, -25.42606, 
    -16.17032, -4.122131, 6.032043, -0.5986938, -10.73856, -17.85182, 
    6.878387, 2.232574, 8.144287, 6.60495, -1.281494, -2.814056, -5.740356, 
    -7.618744, -9.497406, -8.024994, -4.102356, -3.059113, 0.02420044, 
    4.4888, 11.25833, 11.45236, -1.684631, -14.11301, -9.16275, -1.584656, 
    0.2528687, 2.30835, -1.411194, -1.058594, -5.232544, -12.79166, 
    -13.36771, -13.83594, -9.410431, -9.61615, -14.25363, -11.41382, 
    -11.86041, -10.99194, -13.66666, -16.53229, -14.806, -11.26382, 
    -12.31198, -12.26016, -5.985413, -7.358582, -4.63855, -6.603912, 
    -10.24191, -7.291138, -7.918243, -9.840881, -10.62759, -13.29141, 
    -21.53409, -21.03073, -19.65445, -18.55209, -11.56485, -10.15442, 
    -1.461731, -0.3757629, 4.103882, 0.3963623, 7.4646, 8.756775, -4.096375, 
    1.755737, 5.759644, 43.27342, 5.963547, -9.345337, 9.848953, -4.739075, 
    5.686707, 25.13387, 23.85104, 5.425018, -7.004181, -5.109375, -18.00912, 
    -12.07602, -7.827057, -3.182037, -3.813263, -2.867462, -2.265106,
  8.15625, 4.386993, 6.299988, 1.415344, -17.1422, -17.68463, -11.61484, 
    2.409119, 4.979675, 6.736969, 10.14714, -5.748444, -4.751572, 13.32396, 
    0.0723877, 10.75208, 9.63205, 5.315643, 3.06485, -2.286713, -4.449738, 
    -4.716675, -4.739349, -2.492706, -2.341156, 0.1549377, 1.37735, 2.002869, 
    1.075531, -2.083588, -11.90729, -12.60574, -3.161987, 0.9547119, 
    1.714844, -3.078369, -4.886719, -5.170074, -10.38333, -11.34634, 
    -15.83725, -13.84845, -9.269806, -17.10312, -12.94244, -13.00674, 
    -26.50391, -29.11926, -20.85861, -16.72812, -12.01849, -8.299225, 
    -8.570313, -2.378662, -1.078888, -3.559875, 0.4406433, -5.460938, 
    -4.310944, -8.564575, -11.99347, -12.67502, -18.96823, -19.21249, 
    -20.3284, -14.45496, -12.43958, -5.644516, -4.350021, 0.9429626, 
    2.420059, 2.095856, 3.037231, 6.483582, -0.291687, -2.332031, -0.109375, 
    32.10158, 39.16589, 2.552078, -1.814301, 8.161728, 3.545563, 16.56302, 
    22.17239, 16.94583, -10.31277, -9.146637, -10.25259, -8.00885, -5.58725, 
    -4.247925, 1.146362, 4.045837, 3.181, 8.878387,
  9.990906, 4.297119, 0.2033997, -3.73671, -8.461731, -10.78488, -2.739319, 
    9.125, 3.846878, 7.930984, 15.51901, 6.085419, -0.7385559, -0.3882751, 
    1.629669, 1.264313, 1.514832, 7.471619, 2.586456, -0.6989746, -2.179688, 
    2.365875, -3.077606, 1.290649, 0.7697754, 0.882019, -3.688538, -4.246887, 
    -6.109894, -7.126312, -9.031006, -7.233337, -4.378906, -2.019531, 
    -6.443481, -5.501053, -5.184113, -15.82605, -23.18152, -19.0896, 
    -15.69531, -16.28671, -15.95442, -16.8, -21.79037, -26.39374, -39.40547, 
    -40.19244, -28.33098, -22.6823, -15.80417, -10.32683, -5.52684, 
    -2.503387, 4.794281, 2.101563, 0.5924377, -0.7161255, -0.6653748, 
    -8.526306, -9.244019, -13.59271, -16.25494, -10.17032, -14.35443, 
    -6.684128, -1.911194, 5.215363, 4.055725, 6.717438, 10.28201, 7.205231, 
    10.31589, 1.275269, -0.6138, -10.22552, -16.77943, -3.730728, 12.80156, 
    1.767441, 5.151825, 7.930984, 14.33307, 19.12395, 14.02005, 2.683075, 
    -11.15234, -4.755463, -3.422913, -3.514069, -0.1252441, 4.191406, 
    5.245819, 5.416412, 10.33801, 12.23856,
  8.914337, 5.286194, -0.8828125, -13.306, -5.635941, -5.254944, -4.072906, 
    -8.899231, -5.717972, 1.004425, -0.455719, -2.083328, 0.4489594, 
    0.630722, 2.70546, -10.07603, -0.7190094, 7.645309, 5.24115, 7.302338, 
    1.836975, 3.43045, 2.632813, -0.6038818, -1.457031, -6.029175, -9.967712, 
    -9.320587, -7.468231, -7.053375, -12.18542, -6.243469, -3.823456, 
    -5.408081, -0.7945251, -6.834625, -13.72473, -8.356506, -6.369781, 
    -19.97604, -24.54922, -25.33022, -24.81589, -27.39218, -42.94427, 
    -47.40884, -48.31224, -49.11874, -37.63957, -35.19818, -23.3349, 
    -10.56485, -2.336197, -2.669006, 2.961456, 4.5224, 1.612213, -0.7669067, 
    -2.026306, -1.38385, -6.521118, -6.938019, -9.707825, -7.789063, 
    -4.085693, -2.360687, -0.1421814, 3.00705, 8.536713, 11.6586, 18.07867, 
    13.17398, 6.957031, -2.028137, -5.240631, -13.01511, -5.926559, 16.40053, 
    6.571106, 2.911972, 13.3862, 14.24374, 19.03697, 17.91145, 11.52527, 
    -8.194016, -10.67293, -6.789856, -9.4552, -9.4729, -3.459625, -1.161987, 
    5.624725, 7.368225, 11.33282, 13.70053,
  -3.036743, -5.813293, -8.802094, -8.183838, -3.221878, -4.153397, 
    -1.237503, -5.169266, -23.44089, -33.82916, -21.83907, -7.415359, 
    -1.653915, 6.333603, 7.990356, 3.4953, 3.065872, 9.806503, 8.034119, 
    0.5091248, -2.022659, 0.4533844, -2.286987, -3.228149, 1.036469, 
    -1.529938, -4.463531, -6.753143, -7.136978, -10.46719, -13.1711, 
    -8.931763, -2.687759, -4.967972, 2.624741, 4.063019, -6.994522, 1.988022, 
    7.762238, -7.894791, -24.87161, -24.67291, -18.49506, -20.80391, 
    -32.40936, -33.46407, -40.91667, -44.39766, -34.58333, -29.08047, 
    -21.92371, -18.15781, -14.79819, -19.69714, -10.99141, -6.810425, 
    -7.461197, -12.53152, -9.989075, -10.95079, -5.891937, -11.68826, 
    -8.674225, -8.583069, -6.036194, -7.64035, -3.9711, -7.91275, -5.138306, 
    -9.298431, -10.0979, -9.250763, -8.48465, -11.89948, -14.02135, 
    -6.987488, -0.8656311, 8.098175, 8.122665, 1.88829, 11.57657, 9.633331, 
    12.61224, 20.41302, 10.85051, -8.495834, -1.65625, -8.940369, -8.717682, 
    -6.4617, -3.183319, -2.450012, 1.592712, 3.132019, 1.867981, -1.905457,
  -2.052338, -2.823425, -2.641663, 1.557297, 3.481247, 6.234375, 1.2052, 
    -2.312759, -26.95546, -41.26537, -23.98386, -6.898438, -2.459366, 
    3.737762, 3.773438, 6.55574, 0.2255249, -3.334641, -6.196609, -4.603378, 
    -4.133072, -2.796875, -5.371094, 0.5164032, -0.1117096, -4.329956, 
    1.666397, 2.701569, 2.973953, 9.086456, 3.140106, -11.12109, -8.245316, 
    -8.800781, 4.402069, 6.671875, -8.274994, -10.54218, -11.27499, 
    -20.39375, -18.01588, -11.07864, -15.24817, -11.74609, -9.770584, 
    -11.49583, -16.62917, -11.7672, -4.277603, 8.681519, 7.499466, 6.776825, 
    3.392197, -3.802597, -7.722672, -6.2724, -11.05469, -12.48566, -11.83517, 
    -12.60025, -13.22629, -12.49686, -12.87006, -12.30939, -6.410431, 
    -8.71405, -3.671356, -3.479675, -6.56459, -3.109375, -5.938797, 
    -7.304688, -10.05313, -19.21667, 5.266418, 1.482033, -15.36511, 
    -10.16432, -4.942978, 0.3747253, 4.342453, 8.309128, 18.34557, 16.56953, 
    7.750519, -2.919769, -0.2843628, -2.359131, -4.647125, -2.016144, 
    0.002593994, -3.692444, -0.9377747, 1.191132, 4.021088, -1.740356,
  -1.662781, -1.02655, 9.283081, 19.30911, 4.275787, -2.271103, -8.617706, 
    -15.24635, -28.11302, -24.20285, -16.05417, -11.44635, -9.844269, 
    -5.403397, -6.668503, -1.216141, -1.947144, 0.615097, 0.5911407, 
    3.011978, 1.976044, 0.7119904, -1.396362, -3.370056, -5.179153, 
    -7.433853, 9.070313, 3.379166, 2.652344, 8.656509, 0.5622406, -9.733597, 
    -4.469269, -7.133591, 0.6101685, 1.416412, -8.395584, -6.214066, 
    -2.799225, 1.920303, 0.7809906, -1.771347, -1.826035, -4.91095, 
    -6.588287, -5.061203, -0.4682312, 5.389847, 5.068222, 7.057816, 9.555466, 
    13.4203, 14.41354, 12.55026, 9.096878, 5.683594, -1.051544, -4.449738, 
    -5.71405, -7.2435, -7.887238, -7.804138, -6.9375, -7.203644, -5.669281, 
    -4.077362, -1.215637, -0.2229004, -0.3559875, 0.8416748, 2.640884, 
    -5.405212, -7.250778, -19.33542, -16.79193, -8.984894, -24.09427, 
    -15.29089, -11.70755, -6.221085, 7.697418, 15.22736, 22.63333, 10.55626, 
    2.519257, 10.59766, 10.54349, 8.014069, 5.049744, 1.614868, 2.403656, 
    0.6065063, 2.0737, 0.05728149, -0.8486938, -0.9328003,
  -2.837524, -2.396088, 3.860168, 3.600769, -3.5112, -4.560425, -3.916656, 
    -6.581787, -9.446625, -7.916916, -29.68152, -17.48882, -8.563553, 
    0.2885284, 1.655212, -2.36171, -6.373947, -2.74324, 1.537231, 6.316406, 
    3.895569, 4.236984, 4.620056, 0.4505157, -4.877853, -9.677856, 2.754944, 
    5.032028, 6.652603, 9.217438, 0.02838135, -1.425003, -1.989059, 1.154694, 
    3.817703, -0.0619812, -3.182037, -0.9039001, -0.2203217, 1.784378, 
    0.7302094, 0.234375, 2.615631, 2.836716, -0.4880219, 2.433075, 1.949997, 
    1.835159, 1.258331, 1.492188, 4.9375, 3.769257, 3.521881, 8.210678, 
    15.09245, 14.95103, 15.95963, 17.14192, 11.12032, 14.33516, 13.88515, 
    11.77786, 9.740097, 9.241928, 7.745316, 6.214325, 6.825516, 1.440109, 
    3.971344, 1.309372, 4.162506, 5.250259, -4.874207, -18.44009, -22.3521, 
    -23.01198, -7.440109, -2.355988, -5.442963, 22.75339, 12.72084, 23.35678, 
    6.479431, -2.878647, -1.318237, -3.735413, -0.4734497, -0.5593719, 
    0.4825439, 4.778641, 3.244293, -0.1098938, -1.528656, -1.001282, 
    3.077087, -0.3213654,
  -3.549469, -3.628143, -2.513519, -2.473694, -3.492462, -4.922913, 
    -5.269806, -5.341675, -6.099731, -8.833069, -26.1987, -14.2177, 
    -8.860138, -5.711472, 5.996887, 0.6872406, 0.2580719, -1.815369, 
    -0.02812195, 1.162491, -2.3414, 1.886978, 8.843231, 2.870575, 0.4963531, 
    -3.248703, -2.582794, 0.4195404, 1.554947, 0.4130249, 2.839844, 
    -1.825256, -3.606506, 0.8197937, 1.636978, -4.097916, -4.779419, 
    -2.389069, 0.7914124, 2.826813, 2.053375, 2.844788, 5.021088, 9.819534, 
    7.731522, 6.111465, 4.912506, 5.526306, 5.026566, 6.027084, 9.032822, 
    7.430984, 4.992966, 5.902603, 11.36536, 12.72865, 11.28647, 16.55495, 
    18.40547, 23.21849, 23.35782, 22.62968, 23.54922, 18.83151, 17.80443, 
    14.84714, 14.48776, 10.0638, 9.016144, 4.887238, 6.969528, -4.494797, 
    -9.207794, -8.123199, 3.186981, 8.019272, 20.33932, 9.999741, 6.777344, 
    12.12135, 3.688019, 0.5731812, 0.1109467, 0.2932281, -3.972916, 
    -1.692444, -1.425781, 5.713287, 3.737228, 4.646606, 1.988007, 1.267456, 
    1.178375, 2.595291, 1.350525, -1.80545,
  -0.5872345, -0.5760345, -1.537766, -2.016663, -1.922913, -3.155731, 
    -3.555725, -3.9328, -6.191666, -7.749496, -9.524994, -8.037766, 
    -7.058075, -5.440109, 3.024734, 4.248947, 7.57579, 4.061981, 1.264069, 
    -2.012238, -7.856766, 4.142975, -3.563019, 0.3885498, 1.676559, 
    -1.503387, -3.020569, -5.258591, 6.092194, 3.631256, -0.5690002, 
    -4.413284, -2.873962, 0.6903687, -1.640625, -0.6156311, 2.069534, 
    -0.495575, 2.09584, 5.255997, 3.832031, -0.1518097, 2.313278, 3.599731, 
    5.282822, 6.358856, 8.193497, 5.205994, 3.556778, 2.602859, 8.894272, 
    8.374222, 7.601303, 9.181763, 9.131775, 10.75443, 8.102859, 12.66719, 
    16.25313, 14.13229, 16.19218, 19.84947, 18.68489, 16.26848, 14.53204, 
    18.39168, 20.58072, 18.39557, 13.36665, 2.911453, 0.8445282, -6.11615, 
    -4.210938, 12.87839, 6.798187, -1.86824, -5.6362, 0.8916779, 1.556763, 
    -2.998703, -4.053909, 1.726822, 3.382294, 1.139832, 0.2804718, 2.178131, 
    0.9364624, 5.79454, 6.32579, 2.201828, 3.372391, 3.737244, 4.248962, 
    5.855209, 3.277603, 1.730469,
  1.536194, 1.196091, 1.618225, 0.7624969, 0.4346466, -0.3411407, -2.201553, 
    -2.852356, -3.209366, -4.107803, -3.717178, -6.259384, -5.547913, 
    -7.423172, -4.825516, -2.568222, 7.221863, 3.546616, 3.259644, -3.596619, 
    -8.053131, -9.501297, -7.987503, -3.614334, -0.6757813, -1.911713, 
    -4.879425, -5.731506, 1.21875, -2.584106, 1.003387, -0.5164032, 
    -2.804947, -7.621872, -6.087769, -1.540894, -2.327347, -2.871094, 
    0.1213684, -2.933075, 1.219269, 0.6140594, -0.4197998, 4.409637, 
    0.7281189, 4.887512, 3.190369, -1.660416, 1.6073, -1.821365, -0.7984314, 
    5.279434, 2.934891, 9.425003, 7.490097, 7.471619, 6.228394, 7.090103, 
    8.770569, 9.586975, 9.353912, 12.4763, 14.08359, 13.96381, 13.72084, 
    16.756, 19.58932, 18.9034, 13.89661, 6.389313, 2.614075, 19.46797, 
    12.20235, 6.947403, -2.556503, -1.097137, -2.933075, -1.695313, 1.649994, 
    -2.747391, -5.339584, -1.624222, -4.581772, -3.710938, -1.376816, 
    1.026825, 6.115891, 6.127594, 5.773438, 3.509369, 0.5421753, 3.352081, 
    4.236191, 3.033081, 3.454681, 1.020828,
  3.152084, 0.6075592, -0.4255219, 0.5640564, 1.974991, 1.634109, -0.2364502, 
    -1.838531, -2.447662, -2.560944, 1.075516, -6.271347, -8.945053, 
    -5.474213, -3.649994, -5.186981, -2.879684, 3.212234, -0.516922, 
    -4.296875, -7.888031, -12.41927, -8.558319, -6.322144, -4.752869, 
    -0.2171936, -1.18959, -9.142456, -7.424988, -2.303909, -0.5726624, 
    0.3734436, 1.001556, -4.237503, -4.961716, -2.108856, -6.906509, 
    -5.894272, -1.243744, -3.44635, 3.436447, -3.296356, -5.48465, 0.5203094, 
    -1.288803, 1.704163, 3.007294, 3.324478, 3.715881, -0.6687469, -2.077347, 
    7.275528, 6.896606, 4.351303, 5.250259, 6.046616, 4.236984, 2.260941, 
    3.730728, 2.286194, 6.778381, 7.713806, 5.961197, 7.018494, 6.203644, 
    7.862503, 12.99974, 17.97578, 14.36433, 14.47162, 16.43125, 17.98333, 
    6.108597, -0.9614563, 0.514328, -0.5557251, -2.487762, -7.136719, 
    -0.1179657, 0.6890717, -4.978653, -0.910675, -2.720322, -3.451813, 
    -4.098175, -0.9690094, -0.02005005, 4.528122, 2.286972, 4.081512, 
    0.9640656, -0.5471344, -0.8354187, -1.143234, 1.033859, 2.769791,
  -0.45755, -0.6570282, 1.741928, 1.858337, 2.580475, 2.170563, 3.036713, 
    -0.5112, -0.71875, -1.730209, -2.699219, -1.708847, -8.105728, -9.773178, 
    -5.862244, -1.294281, -0.04896545, 7.309113, 4.725784, 1.151031, 
    -2.383331, -5.220306, -4.640625, -6.552597, -7.151306, -5.242981, 
    -1.524216, -13.8737, -9.166145, -0.4432297, 0.5286484, 5.634895, 
    3.670052, 2.263023, 2.496094, 2.501297, 0.2236938, 1.103119, 2.351044, 
    -1.327347, 0.01145935, -0.4104156, -0.408844, -2.215118, -3.20105, 
    0.1171875, -0.640625, 2.046875, 4.1315, -0.5476532, -0.4132843, 4.400787, 
    6.933594, 7.977859, 0.151825, 4.217194, 6.558334, 2.078384, 1.225006, 
    -1.536987, -0.546875, 6.91301, 5.020309, 2.931763, 4.471085, 4.078125, 
    4.700256, 7.446365, 12.88489, 19.37136, 10.00053, 4.017448, 2.988541, 
    -1.206512, -1.456772, -2.723694, -3.440109, -3.148972, 2.359375, 
    -2.470047, -5.661987, -5.148697, -2.997391, -1.244019, -4.015366, 
    -4.394531, 0.2752533, 2.144791, -0.032547, 0.170578, -0.900528, 
    -2.561981, -0.9885406, -1.558853, -2.385162, -1.915894,
  -2.675247, -1.802856, 1.995316, 6.524475, 6.271088, 5.507294, 5.445572, 
    2.107819, -1.007294, -1.465622, -1.472397, -3.361725, -4.20755, 
    -4.335403, -4.872147, -3.419006, 4.194275, 11.49843, 9.760162, 8.718491, 
    6.588806, 3.86145, -0.1906281, -2.929688, -6.332291, -6.888802, 1.496887, 
    -14.02995, -15.50338, 1.074478, -1.625259, -0.8033829, 2.070839, 
    7.461197, 6.168495, 5.223953, 4.961456, 6.094269, 5.907547, 6.950523, 
    6.239853, 4.677078, 4.553391, 3.994522, 2.427078, 2.931503, 1.645828, 
    2.511719, 6.203644, -0.4703064, 3.110931, 0.6984406, 2.103653, 2.53125, 
    -2.996613, 1.443756, 6.566933, 1.625267, -1.199738, 2.937492, 1.410934, 
    1.329422, 1.963028, 0.9666595, 2.652344, 4.359634, 2.062759, 3.435425, 
    6.373962, 7.630219, 6.561203, 3.011459, 1.3013, 0.9593811, 0.4315109, 
    1.927864, 1.940102, -1.856766, -0.8768311, 0.1687622, -1.538803, 
    -4.632034, -8.70105, 0.1125031, 0.674469, -1.728897, 1.143753, 2.290367, 
    5.1586, 5.273438, 2.952332, -0.3184967, 0.1583252, -0.0877533, 
    -0.7416687, 0.3013,
  3.787766, 4.440887, 4.951309, 5.384384, 7.234642, 5.628387, 12.94401, 
    9.49427, 3.551567, 2.245834, 0.4893341, -1.796356, 0.4789124, 0.84375, 
    -4.567184, -6.932297, -4.429169, 0.329422, 6.174744, 6.831772, 4.15416, 
    -2.924225, -3.481506, -3.574738, -1.900513, -0.0765686, -1.812241, 
    -6.486191, -8.630989, 3.95417, -0.1356812, -10.89974, -8.902077, 
    2.412498, 4.126556, 2.674744, 3.077866, 3.498695, 0.4807281, -1.162498, 
    0.08854675, 1.277344, 1.762764, 2.382034, 2.447136, 3.78125, 2.25573, 
    1.267189, 1.330467, 1.392708, 4.947655, 2.744011, 1.471092, -0.5239563, 
    -3.236977, 0.296875, 2.433594, 2.849998, 1.684372, 1.285156, 2.205467, 
    2.626305, 2.230728, 1.602615, -1.104691, 1.466934, 3.393478, 1.812241, 
    4.520309, 0.7203217, 0.4273453, -3.278381, 1.24662, -1.414581, -3.242706, 
    -4.781769, -1.100006, -0.434639, -1.115623, -2.092194, 0.02083588, 
    -0.0851593, 1.388542, 0.9127655, 0.3440094, -0.6531296, 1.823959, 
    3.326561, 4.435417, 1.753128, 1.631767, 3.828384, 4.562241, 0.0838623, 
    2.173172, 3.354431,
  7.694267, 12.91511, 13.73515, 9.703384, 6.412758, 9.495834, 8.724739, 
    5.159378, 8.563286, 4.107811, 4.271095, 3.214584, -1.378647, -0.5286407, 
    -1.062759, -5.490883, -7.857025, -1.846092, 2.587761, 1.553642, 
    -2.730988, -4.143997, -3.37291, -4.171616, -6.032547, -5.723434, 
    -3.800781, -2.718491, -1.180992, 0.779686, -3.199997, -6.491669, 
    -4.876823, -2.439583, -3.353127, 0.5835953, -1.04557, -1.419266, 4.34375, 
    0.640625, -0.06848907, 1.769005, -2.333328, -2.245827, -2.826561, 
    -0.8346329, -1.539581, -2.50235, -1.185936, -3.585159, -2.251305, 2.5, 
    2.478386, -0.5716095, -0.7528687, -2.767189, -3.829422, 1.438797, 
    -1.089584, -3.928383, -0.7687454, 1.13073, -1.368484, -2.032295, 
    -2.911194, -1.567711, 0.9927063, -0.4854202, -1.000519, -0.8822937, 
    -1.627609, -4.585938, -3.026566, -3.572914, -4.319794, -1.756508, 
    2.773964, 2.742706, 1.027344, -0.6299515, 0.3000031, 0.2651062, 
    -0.1119843, 3.426819, 1.079689, 0.441925, 0.7572937, 3.881248, 1.794266, 
    -3.789841, -0.8776016, -1.506767, 2.637505, 2.750519, -0.1567688, 3.001564,
  5.013802, 6.403641, 10.89505, 7.997398, 5.273964, 3.58828, 0.5075455, 
    0.1752548, 4.12188, 3.285938, 2.202347, -3.861198, -5.995316, -3.182289, 
    -3.377869, -3.870834, -3.715103, -5.162498, -3.0513, 1.098694, -1.416405, 
    -5.027084, -5.682549, -2.5112, -3.629692, -5.24115, -5.078644, -2.831245, 
    -2.787239, -2.937759, -2.73333, -1.487762, -2.050781, -5.371872, 
    -5.075516, 0.7390594, 1.804947, -4.390625, -1.1875, -2.670311, -3.78854, 
    -0.5046883, -1.960159, -1.719536, -4.139328, -3.238022, -3.024223, 
    -3.785683, -2.521614, -2.429955, -0.9997406, -0.1260376, -3.587242, 
    -1.864059, 0.2479095, -0.5223999, -0.03541565, 1.004425, 1.369278, 
    0.6658859, 1.003387, 0.7695313, 1.060158, 0.4986954, -4.967186, 
    -4.522133, -3.501564, -3.56823, -5.151825, -4.374474, -2.751305, 
    -5.71067, -5.457291, -3.26432, -2.185158, -2.657288, -3.577866, 
    -1.063278, 3.524223, 1.988281, -1.164063, 1.697395, 0.9283829, 0.8658829, 
    0.5757828, -3.317192, -2.437241, -1.091148, 0.2322922, -0.8671875, 
    -3.455727, -3.191147, 0.6315079, -0.5630264, -1.248962, -1.035942,
  -1.018749, 0.7213593, 0.4614563, -1.942448, -2.381767, -2.102345, 
    -5.280209, -2.52943, -2.294533, -0.6010437, -0.6677094, -2.528126, 
    -2.151566, -1.651299, -4.636459, -6.590363, -7.283859, -12.20339, 
    -7.666145, -5.909378, -4.19088, -4.591667, -4.767708, -4.836983, 
    -4.306252, -4.085938, -5.009895, -4.513542, -4.2388, -2.482811, 
    -1.786194, -2.746613, -2.146873, -1.993752, -3.800514, -3.122658, 
    -2.825783, -3.164322, -1.891144, -3.58073, -3.965626, -2.002865, 
    -2.173695, 0.06015396, -1.629166, -2.688282, -1.619007, -0.5544281, 
    -3.403645, -4.933075, -3.105469, -2.366146, -2.700001, -0.6044273, 
    -0.717968, 0.9320297, 1.744011, 1.51302, 1.763283, 1.429688, -1.141666, 
    1.39505, 2.275257, 3.160938, -0.5010452, -1.777081, -3.065624, -3.774994, 
    -1.861717, -2.323433, -5.739326, -6.200264, -9.270309, -8.14323, 
    -5.730206, -5.172916, -4.067451, -2.480469, 0.5846405, 1.493229, 
    -0.1947899, 1.091408, 0.05989456, -2.956512, -2.754948, -2.938801, 
    0.8846359, -0.6880188, -1.093487, -1.009377, -2.340885, -1.394791, 
    -0.105732, -3.870834, -6.103127, -5.850262,
  -5.266148, -5.603649, -6.88932, -7.971355, -6.635677, -4.485939, -2.45573, 
    0.01250076, -4.530991, -4.602345, -4.037243, -5.613281, -5.046875, 
    -2.693489, -4.993752, -5.098698, -4.634113, -5.866928, -4.842186, 
    -5.450779, -4.276043, -4.378384, -3.178383, -3.348183, -4.569271, 
    -4.572914, -5.353127, -3.098183, -3.081764, -4.543488, -3.942444, 
    -4.871353, -3.160156, -3.155983, -4.555988, -4.738808, -1.206245, 
    -1.797653, -1.90078, -5.025257, -3.197395, -1.236458, -2.03698, 
    -0.2315102, -0.3151016, -2.657291, -2.632553, -2.428123, -1.910938, 
    -0.1104164, -1.114323, -2.687759, -2.616928, -0.814064, -1.953648, 
    -3.868229, -0.7765617, 0.2661438, -0.3158836, -0.6283836, -1.020832, 
    1.936459, 5.481251, 2.10677, -1.061718, -0.8041649, -2.247658, -2.363541, 
    -1.458076, -0.9994812, -2.248699, -2.522915, -2.243229, -3.629425, 
    -2.927605, -3.708073, -5.952084, -4.322395, -1.821095, -1.344013, 
    0.5916672, 0.5096359, -0.8541679, -1.096355, -1.002342, -0.9919281, 
    -0.2252579, -1.489063, -1.53125, -1.56953, -2.954945, -3.398956, 
    -3.022919, -2.663544, -3.366146, -4.910416,
  -1.589844, -4.067448, -4.269011, -4.563541, -2.098959, -3.218229, 
    -3.773438, -2.629686, -2.395311, -1.335676, -2.182552, -5.166407, 
    -4.63047, -4.349739, -3.632549, -4.775782, -3.540886, -1.93568, 
    -0.283596, 0.07734299, -1.370312, -2.948177, -2.302868, -2.892708, 
    -2.471874, -3.066669, -4.647655, -5.465626, -4.61797, -3.850521, 
    -4.041409, -3.194271, -3.472656, -3.817188, -3.678127, -1.630207, 
    -1.933853, -2.728909, -7.20052, -4.501041, -0.7835922, -0.2447929, 
    -1.77969, -1.513544, -0.8799477, -0.5750008, -1.90052, -1.947138, 
    -1.422394, -1.052864, -1.679428, -2.203384, -0.7192726, -0.1291656, 
    -0.01458359, -0.2432289, 0.2294273, -0.7263031, -0.9721336, 0.3054695, 
    1.210938, 1.755728, 0.5348969, -0.08463478, -0.6098957, -2.017708, 
    -0.7257843, -0.1630211, 0.07265472, -1.215103, -1.788803, -1.266148, 
    -1.397919, -2.758335, -4.047655, -4.15625, -4.793749, -5.05703, 
    -4.284634, -3.487759, -0.6132813, 0.1549473, 0.2406235, 1.701561, 
    -1.282553, -0.4466152, 0.2117195, -1.594791, -1.802086, -1.511459, 
    -2.771355, -3.032551, -1.758595, -1.465626, -1.070313, -1.335678,
  -0.1507816, -2.211458, -3.187241, -4.101824, -3.754686, -3.207813, 
    -3.255468, -3.902344, -1.920313, -1.348438, -1.882032, -1.521875, 
    -2.896355, -3.048437, -3.580729, -1.95599, -0.4065094, -0.4979172, 
    -0.9697914, -0.566927, 0.3976555, -0.1135426, -1.513021, -3.004688, 
    -3.354427, -2.503386, -2.717188, -3.712502, -3.642448, -3.282291, 
    -3.024218, -2.954947, -2.769793, -2.746355, -3.011457, -2.775002, 
    -2.870573, -4.740625, -8.213022, -5.76302, -3.073177, 0.3533859, 
    0.9742203, -1.557814, -1.880728, -1.395834, -0.3119793, 1.010418, 
    1.146095, 0.9841137, 0.3341141, -0.2861977, -0.5023441, -1.21875, 
    -2.626564, -2.030991, -0.7338524, -1.103645, -0.5309906, 0.8768234, 
    1.331772, -0.001823425, -0.1906252, 0.2914047, 0.4299488, -0.8200512, 
    -1.368229, -0.9036465, -0.2236977, -0.4249992, -0.3781242, -1.357292, 
    -3.053907, -4.46875, -5.940365, -9.253906, -6.391666, -5.439583, 
    -3.401041, -3.249477, -3.475, -4.610418, -0.9804688, 0.2721348, 
    -1.217447, -0.9320316, 0.2320309, -0.05520821, -0.9825516, -0.2890625, 
    -0.5817699, -0.8687515, -1.71875, -1.664845, -0.8109379, 0.006250381,
  -0.8684893, -1.127343, -1.428386, -1.063802, -1.420312, -2.036979, 
    -1.262761, -0.9020834, -0.5346355, -1.635677, -2.229426, -1.778386, 
    -1.196615, -1.407292, -1.859115, -1.398958, -0.8947916, -0.5755205, 
    -0.4096355, -0.375, -0.9445314, -1.204167, -1.027864, -0.8471355, 
    -1.046875, -1.938021, -1.805729, -1.396093, -1.338542, -1.871354, 
    -2.490625, -1.970833, -1.736198, -2.215364, -2.360416, -1.889845, 
    -1.88698, -3.813803, -6.263541, -5.939061, -5.171875, -3.81927, 
    -2.186458, -0.9153652, -0.7302084, 0.2057295, 0.4557285, 0.1716146, 
    -0.02682304, -0.4539061, -0.2895832, -0.6703129, -1.121094, -1.270312, 
    -1.345052, -0.9830723, -1.197657, -1.388281, -1.295833, -1.012239, 
    -0.959115, -1.185938, -1.342969, -0.7919264, -0.6955729, -0.6950521, 
    -1.042188, -1.090365, -1.520573, -1.954688, -3.084115, -3.439063, 
    -5.691928, -6.149218, -6.307031, -6.361198, -4.501303, -2.961458, 
    -1.951563, -2.345572, -4.554949, -3.385677, -1.836198, -1.121354, 
    -1.692448, -1.211719, -0.8075523, -0.01484394, 0.09895897, -0.3153648, 
    -0.6013021, -1.18177, -1.109635, -0.917448, -1.337239, -1.015885,
  0.03541708, 0.2791667, -0.3539062, -0.8658855, -0.8934896, -0.9229169, 
    -0.9213543, -1.015885, -0.8356771, -0.7229171, -0.676302, -0.7023439, 
    -0.9010415, -0.6377606, -0.4710937, -0.6062503, -0.7122397, -0.4825521, 
    -0.1742187, 0.1736979, -0.005208015, -0.5976563, -0.5898438, -0.3867188, 
    -0.2661457, -0.4854169, -0.6591148, -0.6989584, -0.5322914, -1.090104, 
    -1.271615, -1.009635, -0.8057294, -1.057552, -1.332552, -1.096614, 
    -0.4325514, -0.7674484, -1.314583, -1.596615, -1.030468, -0.6221356, 
    -1.015365, -1.008073, -0.7057295, -1.127604, -2.365886, -2.938542, 
    -2.672656, -2.979167, -3.294791, -3.294011, -2.323177, -2.077083, 
    -2.242709, -2.207031, -1.948958, -1.665364, -1.633333, -1.81875, 
    -1.508594, -1.477604, -1.146354, -0.8809896, -0.8114581, -1.040104, 
    -1.094792, -1.196094, -1.309115, -1.865104, -2.336459, -2.938802, 
    -2.738281, -2.969792, -3.159896, -2.959636, -2.426302, -2.272396, 
    -2.320313, -2.159115, -2.298698, -2.200781, -1.900521, -1.623178, 
    -1.255208, -0.8388019, -0.4049482, -0.03515625, -0.4445314, -0.4458332, 
    -0.3416662, -0.2875004, 0.2236977, 0.05234385, -0.2403646, -0.0406251,
  0.103125, 0.2304688, 0.2101561, -0.001822829, -0.0789063, -0.1104167, 
    -0.375, -0.421875, -0.321875, -0.1033853, 0.01588547, -0.1234375, 
    -0.2541667, -0.2046875, -0.01510417, 0.09921873, 0.1466146, -0.1565104, 
    -0.2210938, -0.1697916, -0.1432292, -0.07291663, -0.0526042, -0.0583334, 
    -0.0234375, -0.1463542, -0.2507812, -0.0859375, -0.1083331, -0.2770834, 
    -0.2932291, -0.3151041, -0.2445314, -0.2080729, -0.2947915, -0.3268228, 
    -0.3651042, -0.5309894, -0.5671875, -0.6166668, -0.5046874, -0.4351562, 
    -0.4088542, -0.4065105, -0.3023438, -0.1515627, -0.1096356, -0.2752604, 
    -0.3104167, -0.3606772, -0.5557293, -0.8390625, -0.5929687, -0.4791667, 
    -0.4257813, -0.5286458, -0.4523439, -0.4796875, -0.4614582, -0.475, 
    -0.4570313, -0.5690105, -0.5421876, -0.4783854, -0.4203124, -0.4486978, 
    -0.5929688, -0.6721354, -0.8041666, -0.6815104, -0.7356772, -0.8005207, 
    -0.8497396, -0.9502604, -1.014844, -0.8820312, -0.6908855, -0.6929686, 
    -0.6927083, -0.6729167, -0.8059897, -0.6265626, -0.454427, -0.484375, 
    -0.3757813, -0.3677083, -0.2434895, -0.1067709, 0.0539062, 0.03880215, 
    0.0369792, -0.008593798, 0.07343757, 0.02083337, -0.1218749, -0.009635329,
  -0.0005208403, -0.00442709, 0.009895831, 0.02552083, 0.03411458, 
    0.03463542, 0.00833334, -0.001562506, -0.01432292, -0.02786458, 
    -0.03463542, -0.04583333, -0.06432292, -0.06119792, -0.05078125, 
    -0.02447917, -0.0005208254, 0.00390625, -0.0109375, -0.02968751, 
    -0.03203125, -0.04479165, -0.01796876, 0.001041666, -0.02135417, 
    -0.04010417, -0.03723958, -0.02890626, -0.03229167, -0.02109376, 
    -0.0252604, -0.04453126, -0.04322916, -0.04088542, -0.03697917, 
    -0.0440104, -0.04921874, -0.07213542, -0.06796876, -0.06015624, 
    -0.03854166, -0.03932291, -0.05546877, -0.04427083, -0.03593749, 
    -0.02395834, -0.01744792, -0.01093748, -0.009895831, -0.02968749, 
    -0.04010415, -0.06979167, -0.09739584, -0.08151039, -0.07682294, 
    -0.09348957, -0.09661458, -0.09114581, -0.08723956, -0.07135415, 
    -0.0809896, -0.1195312, -0.09192708, -0.09765625, -0.08828124, 
    -0.06796873, -0.05755207, -0.08203125, -0.1286458, -0.1567708, 
    -0.1286458, -0.0984375, -0.1054688, -0.1598958, -0.146875, -0.1669271, 
    -0.1460938, -0.1414063, -0.1393229, -0.1481771, -0.07942706, -0.05364582, 
    -0.03958333, -0.04062501, -0.05963543, -0.06510416, -0.06093749, 
    -0.03671876, -0.03932291, -0.04296875, -0.05260417, -0.07187501, 
    -0.06822917, -0.01927082, 0.02135417, 0.01744792,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.8721313, -1.361191, -2.031509, -2.78125, -3.566666, -4.37709, -5.153641, 
    -5.73204, -6.048187, -6.302094, -6.567978, -6.748962, -6.908066, 
    -7.122925, -7.279175, -7.308594, -7.447662, -7.508865, -7.707809, 
    -7.977859, -8.234894, -8.513016, -8.786194, -8.987228, -9.166412, 
    -9.415115, -9.63829, -9.957565, -10.09975, -10.25938, -10.32265, 
    -10.37265, -10.59479, -10.76901, -11.13959, -11.60078, -12.19688, 
    -12.60184, -12.84166, -13.34584, -13.89818, -14.45338, -15.24713, 
    -16.13751, -16.96249, -17.52448, -18.02552, -18.33176, -18.88177, 
    -19.47421, -20.01432, -20.43672, -20.76588, -21.18333, -21.38203, 
    -21.47292, -21.30624, -21.14766, -21.01823, -20.69661, -20.12344, 
    -19.41093, -18.51953, -17.71354, -16.63698, -15.33255, -13.87682, 
    -12.4836, -11.26563, -10.0052, -8.676041, -7.474228, -6.117447, 
    -5.103119, -4.280472, -3.286194, -2.015884, -0.8713531, 0.1770782, 
    1.445831, 2.377853, 3.128906, 3.642441, 4.098694, 4.327072, 4.29921, 
    4.090363, 3.78334, 3.463287, 3.009125, 2.416397, 1.931244, 1.623962, 
    1.146347, 0.5065155, -0.1755066,
  -7.295319, -8.288803, -9.511719, -10.58566, -11.63228, -12.67969, 
    -13.26614, -13.40573, -13.66588, -14.41119, -14.61121, -14.46277, 
    -14.60782, -14.75677, -15.42682, -16.36771, -17.29088, -18.10728, 
    -18.72292, -18.85834, -19.08099, -19.28073, -19.26927, -18.75391, 
    -17.84714, -16.74844, -15.28854, -13.34064, -11.45364, -9.960938, 
    -9.135422, -8.958069, -9.160156, -9.862244, -11.07892, -12.26251, 
    -13.24765, -14.30495, -15.39766, -16.30313, -16.74323, -16.89244, 
    -17.14713, -17.26302, -17.39973, -17.36926, -17.99505, -18.56145, 
    -19.50313, -20.88594, -22.08723, -22.38776, -21.84531, -20.75182, 
    -19.75495, -18.80078, -17.19245, -15.64635, -14.39973, -13.48568, 
    -12.49088, -11.03099, -10.0414, -10.04245, -10.33308, -9.846611, 
    -9.238014, -8.758591, -7.955467, -7.492973, -6.649475, -5.777863, 
    -4.459381, -2.807297, -1.407288, -1.220306, -0.6445313, -0.2705688, 
    0.3421936, 1.619522, 2.831512, 3.976028, 5.297394, 5.880219, 6.057281, 
    5.963287, 5.478119, 4.251038, 2.985931, 1.883087, 0.1046906, -1.4599, 
    -2.615891, -3.524216, -4.5737, -5.876556,
  -10.09036, -11.54532, -12.74454, -15.00703, -17.75781, -19.81302, 
    -21.21797, -21.7065, -21.26172, -20.16641, -19.39948, -18.64114, 
    -17.59193, -16.34843, -15.36354, -14.83151, -14.0724, -13.76537, 
    -13.40157, -13.43568, -13.35391, -13.12161, -12.97682, -12.88959, 
    -13.0573, -13.31328, -13.55234, -13.78073, -13.60989, -12.85599, 
    -12.39114, -12.48645, -12.66745, -12.52942, -13.07629, -13.22943, -14.05, 
    -14.42891, -14.34869, -14.1599, -13.55911, -12.75938, -12.38594, 
    -12.12004, -11.89792, -11.70808, -11.1888, -11.2164, -11.34792, 
    -11.25417, -12.77552, -14.12786, -14.40573, -13.53542, -10.12318, 
    -7.428383, -5.156769, -3.8862, -2.825005, -2.082031, -2.106781, 
    -2.345322, -2.574226, -3.006248, -3.642448, -5.851563, -6.802597, 
    -5.576828, -4.797653, -4.424469, -5.516418, -6.516922, -6.613815, 
    -5.377609, -4.596344, -4.251038, -3.583069, -2.304688, -1.635941, 
    -1.059113, -0.4213562, -0.08308411, -0.6015625, -0.6906281, -1.216675, 
    -2.379944, -3.417709, -4.863022, -5.568497, -6.419281, -7.220322, 
    -6.615891, -6.224213, -6.444534, -7.302597, -8.291656,
  -11.52682, -11.73282, -13.16484, -14.73567, -16.21536, -16.23854, 
    -14.84973, -14.37526, -14.14009, -13.37213, -12.79089, -11.96225, 
    -10.35104, -9.491135, -8.681763, -7.107285, -6.596878, -5.810944, 
    -4.992188, -4.094788, -3.478638, -2.985413, -3.190109, -4.169266, 
    -5.912491, -8.277603, -11.02786, -13.03619, -14.24532, -15.57474, 
    -16.52525, -15.55937, -13.74973, -11.78749, -10.04036, -8.191925, 
    -6.963547, -8.138535, -11.76457, -13.82448, -15.00363, -15.39975, 
    -15.21562, -16.60312, -17.15677, -17.74297, -17.86693, -15.64973, 
    -16.1539, -13.72186, -12.25548, -12.25287, -12.38333, -10.7289, 
    -7.577858, -5.68541, -4.383331, 0.2898407, 0.4197922, 2.0914, 3.4198, 
    3.048965, 2.055466, 0.7419281, -0.2338562, -1.069534, -2.583328, 
    -3.861465, -3.603653, -2.300262, -1.844269, -2.369019, -1.869537, 
    -2.993759, -2.619537, -0.6869812, 0.3966217, 0.89505, 2.29895, 2.532806, 
    0.3945313, -0.4690094, -3.434128, -6.437759, -8.119797, -7.759903, 
    -6.023438, -6.569016, -6.423691, -7.5065, -9.122131, -9.739319, 
    -11.31718, -12.16432, -12.70105, -11.9875,
  -5.628387, -7.114594, -9.947403, -11.825, -12.45522, -13.0638, -13.86615, 
    -13.95807, -12.63046, -12.5573, -12.98828, -14.28673, -15.56927, 
    -14.82344, -10.575, -4.916412, -1.961716, 0.3721466, 1.810669, 1.231522, 
    1.331253, 1.387238, 0.3507843, -0.7424469, -1.463791, -1.554688, 
    -2.945572, -4.764587, -4.198959, -5.528641, -7.874481, -8.17865, 
    -6.485672, -5.178131, -5.482819, -5.507553, -4.769272, -3.263535, 
    -3.105728, -5.04921, -6.564056, -7.149216, -7.02475, -6.991394, 
    -5.628128, -4.347916, -5.798187, -1.842972, 2.835159, 2.748947, 0.9888, 
    0.170578, -1.6409, -4.037498, -5.148705, -6.441673, -9.33255, -12.12163, 
    -13.45651, -14.94376, -13.8013, -12.1422, -10.88463, -9.888535, 
    -9.213547, -8.838028, -7.184113, -4.868225, -3.723434, -2.782288, 
    -1.916397, -7.156769, -7.830994, -7.369537, -6.166931, -3.901566, 
    -0.7820282, -0.2406311, 0.3885498, 0.2640533, -0.6075592, 2.130203, 
    0.3408813, -3.344528, -6.588013, -9.445831, -11.04947, -11.94688, 
    -12.57552, -12.52188, -14.59088, -5.015884, -4.867706, -4.778641, 
    -6.36145, -6.761459,
  -5.074738, -5.2276, -4.027863, -3.288803, -2.733078, -2.426559, -3.204956, 
    -3.979172, -7.166412, -6.496094, -6.157562, -8.726822, -14.08099, 
    -16.06328, -11.63307, -6.563278, -3.304428, -2.444534, -3.951828, 
    -4.114059, -1.680206, -0.2929688, 0.8895874, 0.3463593, -0.0377655, 
    -0.9242249, -3.701035, -4.603653, -7.560669, -12.63385, -16.05678, 
    -17.56537, -15.83333, -11.44193, -6.792191, -1.805481, 3.508591, 
    5.330719, 5.386459, 4.164841, 2.085419, 0.170578, -0.9492188, -1.552872, 
    -2.876038, 1.75235, 0.5361938, -2.261192, -3.566406, -5.024483, 
    -4.696091, -5.973434, -7.157555, -6.346619, -6.021347, -6.426559, 
    -8.194534, -11.04063, -15.49166, -15.19167, -14.29244, -13.68542, 
    -14.27423, -16.7336, -15.49089, -14.22083, -9.539063, -3.922134, 
    -2.320831, -3.971619, -4.915359, -6.016663, -3.355209, -3.610153, 
    -2.077866, 0.5343781, -0.2002716, 1.138016, 2.853394, -1.696091, 
    -10.87265, -11.86719, -16.2724, -23.08881, -29.16692, -32.20442, 
    -31.37709, -29.63881, -26.36745, -24.91406, -23.17917, -21.24454, 
    -20.5349, -22.56979, -17.32292, -12.1086,
  -31.20938, -33.26407, -33.30756, -26.3073, -19.24037, -13.29767, -11.81017, 
    -12.7112, -12.73178, -12.15364, -17.3013, -26.27499, -28.70834, 
    -30.42082, -25.44844, -19.15468, -13.82031, -14.22031, -14.80963, 
    -13.46718, -13.51198, -13.67004, -10.42552, -9.870575, -7.235428, 
    -4.154434, -9.253387, -13.58932, -12.51224, -15.42162, -19.15364, 
    -23.60521, -22.35287, -21.36328, -16.02318, -14.50233, -26.98932, 
    -6.889847, -1.047409, -1.038025, -3.295837, -5.595581, -6.030731, 
    -6.411713, -2.791138, -1.316147, -2.429153, -3.253647, -0.2617188, 
    1.5578, 2.556778, -2.763535, -9.920059, -12.34116, -11.67578, -10.77109, 
    -10.12213, -11.39738, -13.79897, -12.47682, -5.08905, -2.317184, 
    -2.142715, -6.698181, -10.95573, -8.649994, -6.223953, -6.741409, 
    -4.758591, -2.132813, -0.4395752, 3.132813, 2.750259, -1.757553, 
    -4.229172, -3.973953, -3.609634, -3.870316, -3.186447, -7.523697, 
    -21.41302, -20.325, -16.55339, -13.87553, -8.635422, -9.860153, 
    -14.48698, -18.91614, -19.65755, -20.16512, -25.92004, -30.67188, 
    -31.6039, -26.86848, -24.10391, -27.64531,
  -6.023438, -0.3552094, 0.4476624, -2.809891, -6.73645, -3.178116, 
    0.8377533, 2.553909, -0.3807373, -2.836456, -4.120056, -4.204697, 
    -5.396866, -7.614838, -4.954422, -5.328384, -4.663803, -6.886978, 
    -9.782806, -8.129684, -7.813538, -9.403381, -10.78645, -13.28801, 
    -4.711716, -0.02812195, -0.4268188, -1.538284, -3.499481, -5.454422, 
    -10.62917, -10.95522, -9.18306, -8.051559, -6.456772, -5.320572, 
    -7.289841, -7.204697, -8.771866, -5.682541, -5.191147, -2.307037, 
    -2.118744, -4.304688, -0.8203125, 0.883606, -0.8981781, -3.910156, 
    -6.889587, -6.579422, -8.149475, -9.501038, -8.817703, -7.1138, 
    -8.292969, -11.71849, -11.2039, -9.802597, -11.84584, -15.4823, 
    -12.59714, -9.087753, -7.391144, -5.047134, -1.759109, -5.236984, 
    -7.760681, -10.67032, -10.17969, -5.789581, -1.205215, 1.286972, 
    2.538788, 1.531509, -0.3078003, -2.222656, -2.833862, -8.679169, 
    -8.975769, -3.713287, -1.943481, -6.288528, -11.68646, -12.58516, 
    -8.889053, -8.176041, -11.51431, -12.09714, -13.19896, -8.481247, 
    -5.054947, -3.997131, -4.31041, -5.199478, -5.374481, -8.657547,
  -8.473953, -4.510941, -4.123428, -10.02214, -12.05547, -7.020309, 
    -1.597397, -0.9442749, -1.644012, -2.971878, -5.910156, -7.795319, 
    -5.066666, -5.653381, -6.763535, -6.4487, -4.059631, -4.269272, 
    -5.715363, -6.196091, -3.263794, -6.867966, -11.62839, -9.004944, 
    -3.409103, -1.011978, -2.445572, -5.7789, -7.034637, -5.437759, 
    -4.794006, -2.295578, -0.6070251, -1.351303, 1.059372, 4.450775, 
    4.173965, 1.529419, -2.369278, -4.671616, -4.140625, -1.9599, -2.758072, 
    -5.121613, -4.21875, -0.1765594, -1.712234, -2.939056, -3.570053, 
    -5.031509, -7.858337, -6.016663, -6.071884, -7.53801, -10.10469, 
    -7.890884, -7.3237, -8.585938, -6.975769, -6.816925, -7.857819, 
    -7.415894, -7.297409, -6.585159, -2.169785, -0.2052155, -2.858078, 
    -3.52005, -1.877609, -0.7773438, -2.853653, -3.015884, -2.58725, 
    -4.443237, -5.013535, -4.034103, -6.391678, -5.650513, -4.585159, 
    -0.8859406, -2.028656, -4.636459, -5.976822, -7.671875, -4.080719, 
    -6.765884, -12.01979, -12.45676, -8.666656, -8.834366, -11.65964, 
    -10.96979, -11.19348, -8.884628, -8.985153, -9.927094,
  -10.21327, -8.256256, -6.678391, -7.713806, -4.699478, -2.910934, 
    -1.144531, -1.441925, -0.6385345, 2.516144, 0.5622406, -3.258331, 
    -3.067963, 2.569534, 6.571625, 6.68074, 7.670319, 7.297653, -1.342712, 
    -2.565094, 4.505219, 4.866928, -2.852341, -4.558334, -3.614059, 
    -0.9401093, 2.945053, 3.130997, -1.584641, -8.172653, -9.138535, 
    -3.476303, -0.6010437, -3.199997, -7.110413, -4.729431, -2.582291, 
    -5.073959, -0.6364594, -0.08932495, -2.95079, -4.05365, -4.593491, 
    -2.999222, -0.8809967, -3.61145, -2.834366, -3.046097, -5.551041, 
    -3.249222, -4.126572, -2.569794, -2.655457, -4.019272, -6.043228, 
    -2.608337, 2.551559, 3.160416, -0.9864502, -7.291153, -10.30209, 
    -3.68074, -1.653122, -2.249222, 0.5020905, 0.6114502, -5.171082, 
    -9.44635, -6.358582, -3.771088, -3.374481, 3.201569, 1.286713, -3.648178, 
    -1.854691, -3.200775, -3.112228, -2.058594, -3.114838, -4.666153, 
    -2.997665, -5.203903, -6.617706, -4.890625, -4.119019, -5.5289, 
    -5.860413, -4.929688, -1.383072, -7.026566, -5.632813, 0.5260315, 
    -0.9385376, -5.420837, -8.132019, -7.820313,
  1.68959, 0.0705719, -0.1526031, 0.7723999, 1.821869, -0.2687531, -1.413788, 
    0.9552155, 1.8302, 2.995834, 7.568756, 7.26355, 5.764847, 6.783585, 
    5.733597, 4.876816, 4.744522, 0.3312378, -1.873688, 4.714066, 4.856506, 
    2.744537, 3.052856, 3.496094, 6.544525, 3.363541, 3.238022, 6.778397, 
    0.6585999, -2.437759, -3.252075, 0.5164185, 2.359894, -1.797134, 
    -2.784897, -6.021606, -4.030212, -1.471085, 0.6184998, 6.670059, 
    7.163284, 4.379684, 4.313538, 5.184891, 2.02475, 1.133347, 5.353134, 
    13.20651, 13.74713, 3.789841, 4.354691, 4.033844, 4.627075, 1.708847, 
    -2.722656, -6.184113, -5.063797, 0.2065125, -1.20546, -1.320572, 
    -3.753128, -1.924744, 1.25209, 4.746872, 4.463547, 0.5929718, -2.37265, 
    0.9104156, 3.4776, 1.074478, -3.315887, -4.303131, -5.698441, -5.31041, 
    -2.179169, 2.058853, 0.7729187, 7.188812, -1.414581, -2.163528, 2.449478, 
    1.123703, -2.020569, -4.199738, -0.2127533, 0.1429749, -2.766663, 
    -1.200775, -0.1580811, -1.093491, -1.921616, 2.089325, 1.713806, 
    -5.924484, -2.405716, 0.6921844,
  1.933334, 5.996353, 6.265366, 5.327866, 7.079422, 5.728653, 7.25209, 
    3.901566, 2.626556, 4.628387, 4.518234, 9.355728, 8.665894, 2.65625, 
    3.996353, 3.291672, 0.7002716, -2.001038, -0.1460876, 3.638535, 3.420319, 
    3.659882, 4.599991, 1.703125, 3.664322, 2.739578, 2.385162, 5.974747, 
    4.440613, -0.6442719, 3.685944, 2.268494, -0.7789154, 4.681244, 2.203125, 
    -1.636719, 2.365631, 4.320053, 4.0961, 0.8101654, 0.5088501, 6.303909, 
    7.870056, 6.933853, 5.581253, 11.256, 9.376816, 11.17838, 4.709885, 
    1.814316, 4.498962, 4.301559, 2.371613, 2.614319, 0.7156219, 2.671875, 
    -4.119278, -2.4823, -0.1273346, 7.193481, 5.603119, 0.5244904, 0.6354065, 
    0.4424591, 0.5643158, -2.036972, -0.6596375, 0.1489563, 1.238281, 
    -1.803635, -3.8013, 0.7320251, -2.320313, 2.182037, 8.110947, 6.740616, 
    13.56874, 28.0974, 20.56667, 5.596619, -2.3414, 0.1481781, 0.5554657, 
    0.4781342, 2.326035, 3.140366, 1.263809, -0.005477905, 4.9776, 3.409897, 
    0.9888153, 1.137772, 2.104935, 1.326569, 1.679688, 2.647385,
  -0.733078, 0.0776062, 1.280472, 5.180725, 6.964325, 8.892715, 4.067184, 
    4.2677, 10.44376, 11.89192, 3.339844, 5.460678, 6.723434, 2.37735, 
    -0.9312439, 4.315369, 5.309631, 4.879166, 9.046356, 12.32813, 14.0737, 
    11.12631, 9.980469, 9.682297, 10.92056, 10.2216, 11.07813, 7.941925, 
    7.534897, 7.802612, 10.9651, 7.738281, 4.911713, 6.446869, 4.29245, 
    7.266937, 3.026031, 3.836731, 5.385406, 4.818481, 2.897675, -1.675018, 
    2.631256, 7.219803, 8.036453, 13.80989, 19.25676, 9.832809, 11.22525, 
    14.08516, 8.933075, 8.834106, 6.151306, 3.930725, 2.636459, 1.236725, 
    7.203384, 9.672668, 8.110931, 8.784378, 9.254166, 8.790359, 6.403122, 
    5.070053, -0.3406219, 1.566666, 6.452332, 5.35495, 1.942963, 7.173706, 
    2.170319, 2.600525, 5.95079, 6.518494, 7.870316, 5.158325, 28.73647, 
    53.37344, 28.59558, 5.998169, -2.938263, -2.320313, 0.1231689, -5.671875, 
    -5.188293, 2.310669, -1.911469, -5.423431, -4.417969, 0.1078186, 
    1.210678, 5.135406, 1.617447, 1.888535, 3.018219, -1.570831,
  8.331497, 10.24478, 6.757813, 2.157837, -0.5734253, 0.05209351, 1.138306, 
    3.373688, 2.339569, -0.8919373, 0.39505, 3.679169, 1.86615, 1.495056, 
    3.891144, 3.697906, 1.8797, 1.006531, 3.31015, 3.704437, 4.658066, 
    5.502853, 6.027588, 7.728363, 4.644775, 5.389587, 6.708832, 4.283081, 
    2.2388, 2.819519, 2.652588, 5.327087, 6.11145, 4.138275, 4.443756, 
    3.807281, 1.222412, 6.329163, 20.84689, 18.81119, 7.498932, 0.3932495, 
    3.474213, 7.197906, 0.7401123, 3.783081, 10.76797, 15.09349, 6.228638, 
    2.863281, 1.059662, 0.3828125, -0.1510315, 3.075256, 3.060669, 8.713821, 
    10.62761, 8.330994, 6.650009, 7.720047, 2.175522, 11.79895, 12.0224, 
    6.335678, 4.1539, 8.076828, 7.469025, 12.80208, 11.27345, 6.167725, 
    -0.4315186, 5.72345, 3.773438, 3.397156, 2.53775, 0.5596313, 16.28723, 
    23.95233, 6.814606, -2.516937, -8.9776, -8.174469, -6.1474, -6.300507, 
    -1.251312, -2.024475, -1.784637, -0.6182251, 0.6768188, 0.7505188, 
    -2.081512, -4.318222, -2.703903, 2.752075, 4.603912, 6.008072,
  -2.230743, -5.293488, -7.579407, -7.726807, -6.777344, -1.867981, 
    -6.952362, 0.1763, 1.781494, -3.382813, -1.413544, -2.094269, -6.063293, 
    1.749481, -0.9692688, -7.782013, -9.041687, -5.181244, -0.1348877, 
    -3.435425, -1.60675, 3.414337, -0.6398315, -1.550507, -8.383057, 
    -5.591156, -2.848175, -4.428619, -7.252869, -6.847382, -6.201294, 
    -7.605988, -6.130981, -1.225494, -4.287231, -2.660675, 6.588013, 7.95285, 
    8.845032, 3.652344, -5.7612, -10.85886, -3.871613, -3.208618, -2.182037, 
    -5.756775, -4.50885, -6.529938, -6.440338, -7.581787, -9.652344, 
    -8.206512, -2.492432, -0.6731567, 7.998169, 16.33359, 11.50964, 9.2966, 
    0.5262756, 0.4450378, 3.904419, 7.351837, 4.394531, 4.164063, 5.395844, 
    3.60495, 3.406006, 3.404938, 1.216431, -0.7109375, -1.865356, -5.381775, 
    -4.229156, -4.257813, 1.690094, 4.41745, 1.837738, 2.801819, -0.7049255, 
    -9.947418, -3.524994, -1.081238, -4.439575, -0.9447937, -3.499207, 
    -5.119781, -4.7612, -1.801819, 0.4104004, -1.80545, -2.9375, -1.496338, 
    -4.437256, -2.233856, -0.836731, -1.521881,
  -11.84921, -10.09842, -8.310944, 0.725769, 0.9197998, 0.2255249, -2.283356, 
    2.859894, 5.809097, -2.198456, -2.434631, -4.747406, -6.894806, 1.984894, 
    -4.083588, -8.504181, -8.413544, -6.836212, -1.62735, -8.505463, 
    -5.738037, -8.887756, -11.13959, -10.46588, -5.547913, -8.839325, 
    -12.54138, -8.739319, -8.131256, -3.186981, -5.309875, -6.573181, 
    -4.538788, -4.113281, 0.07525635, 1.096619, 3.481262, 1.45105, -9.2229, 
    -13.67993, -13.54321, -16.27289, -11.37628, -8.690094, -5.675018, 
    -10.5914, -14.59921, -6.965607, -8.025269, -4.025238, -2.802887, 
    -1.128662, 4.598694, 4.905457, 9.570313, 3.825287, -1.420837, 0.377594, 
    -0.40625, 5.191132, 7.195831, 6.104675, 5.639313, 2.896881, 0.1554565, 
    4.134644, 8.107574, 3.519257, -2.664825, -4.912231, -9.537506, -13.29376, 
    -7.013824, -6.513031, -4.791382, -8.813538, -2.334381, -0.9289246, 
    0.7203064, -13.52527, -9.208313, -5.834106, -9.439575, 1.419525, 
    -4.327606, -5.327362, -5.781525, -14.19193, -11.53021, -13.48932, 
    -4.374481, -5.692444, -5.445038, -4.613007, -6.432556, -5.462494,
  -1.997131, -4.596619, 1.370575, -6.001587, -4.247375, -8.098938, -8.383057, 
    10.18803, 11.56979, -5.874207, -10.92343, -7.705719, -8.621368, 
    0.8867188, 2.565369, 3.297119, 0.8994751, -7.096863, -1.493469, 
    -6.117188, -4.767731, -7.463013, -11.64948, -13.69193, -7.074768, 
    -5.997925, -3.118225, 0.2166748, 0.2723999, -5.81665, -9.447906, 
    -11.62787, -5.280212, -4.754944, -7.534882, 0.567688, -2.092194, 
    -7.354156, -12.80026, -17.38333, -18.84195, -16.77759, -5.830444, 
    -8.976288, -3.229431, -6.486176, -11.68152, -6.262756, -0.7619629, 
    -0.102356, -6.23645, -3.660431, 1.376556, -1.234375, -0.2388, 1.715118, 
    2.536438, 3.776062, 7.711975, 6.975006, 4.488037, 4.101837, 2.835693, 
    -1.07605, -0.04870605, -1.49115, -0.9502563, -6.936707, -11.91382, 
    -9.237213, -11.85782, -7.438293, -3.70755, -5.246338, -7.651031, 
    -8.333618, -2.264069, -2.313019, 6.672913, -4.638031, -10.6716, 6.884109, 
    1.46199, 13.89662, 2.412262, -8.4375, -12.22604, -17.44272, -10.85367, 
    -9.661713, -9.895844, -13.80026, -10.7341, -12.25989, -11.60913, -9.701813,
  -4.710419, -5.807037, -7.340881, -6.1026, -10.94922, -10.48776, -1.731232, 
    6.985413, 10.02032, 4.852325, -1.4552, -7.192963, -7.863281, 1.371887, 
    6.674225, 6.775513, 2.429169, -1.428894, 0.9091187, 1.767456, 1.354401, 
    -2.494781, -3.624725, -4.95105, -1.916138, -1.847656, -3.467468, 
    -2.267975, -2.828369, -5.545563, -8.818237, -6.061188, -1.592194, 
    -4.949219, -7.224213, -3.561737, -4.375519, -11.4534, -12.17682, 
    -16.70782, -21.16617, -13.67395, -8.801575, -11.84818, -7.914856, 
    -7.552094, -11.98151, -1.513031, 1.828888, -4.640381, -6.781525, 
    -11.19922, -6.097656, 0.3013306, -0.6598816, 0.01382446, 2.001312, 
    5.095032, 3.320831, 4.119537, -0.8406067, -1.7146, -1.30365, -3.390625, 
    -4.688293, -12.3862, -14.58307, -13.53412, -13.53647, -11.09766, 
    -6.769287, -1.066925, -4.092194, -6.907837, -7.970306, -1.864868, 
    -2.338287, -3.010651, 24.81848, -5.466156, -11.25494, 17.70677, 15.03699, 
    9.652603, -0.05807495, -7.043488, -9.889069, -6.996094, -3.590637, 
    -4.870575, -6.019531, -9.367188, -9.706512, -5.504425, -8.467438, 
    -0.9836121,
  -8.027863, -6.771362, -10.43152, -3.4198, 0.1228943, 5.365112, 9.7836, 
    16.63544, 15.78436, 14.06198, -7.827087, -17.65259, -24.91927, 0.1856689, 
    4.8797, 0.6455994, -6.502594, -6.561218, -0.9494934, 5.661713, -1.242981, 
    -0.9895935, -1.815887, -5.5672, -5.937775, -4.071625, -3.817963, 
    -1.372681, 0.7120056, -1.219788, -4.344543, -6.169037, -2.076569, 
    -2.265625, -8.183075, -8.459381, -10.42734, -12.96329, -13.30106, 
    -12.07135, -13.31796, -8.550781, -13.14896, -12.39609, -9.409119, 
    -13.43958, -9.805725, -6.612244, -7.720032, -4.419281, -6.135162, 
    -13.89999, -14.61719, -14.34268, -6.757813, -2.333588, -2.540619, 
    -0.366394, 0.1580811, -5.3461, -2.415894, -4.101837, -9.070038, 
    -6.447632, -15.65808, -16.37814, -12.88281, -10.75938, -8.043747, 
    -6.931778, -4.775543, -3.06955, -4.223175, -1.391144, 7.740356, 
    -3.511459, -2.940094, -2.006256, 27.14453, -7.270584, -4.564331, 
    7.855469, 8.201813, 8.274734, 2.6427, -0.978653, -4.9104, -0.2539063, 
    -0.0385437, -1.143738, -6.071106, -11.10339, -9.505219, -10.66458, 
    -1.878143, -1.108337,
  6.047638, -2.734894, -2.108612, 4.131256, 5.655472, 3.477875, 7.1315, 
    11.61276, 5.017715, 3.586197, -6.5159, -12.39612, -18.82005, -7.432541, 
    4.116943, 3.732025, -4.914581, -11.02112, -3.124207, 11.35886, 8.451569, 
    4.917175, 1.692444, 0.3234253, 0.272644, 0.7374878, 0.1564941, 2.4422, 
    -4.297119, -7.188019, -1.562775, -4.005219, -1.447418, -2.430725, 
    -11.21747, -16.05054, -15.61639, -20.99402, -22.19766, -16.22006, 
    -20.21042, -13.9966, -20.13438, -18.26927, -12.9211, -13.98282, 
    -14.49298, -13.52605, -7.354431, 2.396088, 1.764053, -10.89844, 
    -15.09193, -15.02527, -8.178925, -3.876801, -0.6911316, -2.434113, 
    -6.190369, -12.74377, -9.131775, -14.36795, -12.08542, -14.29974, 
    -16.25494, -14.05469, -15.96642, -7.781769, -4.265884, -2.449997, 
    -3.070831, -0.9664001, -2.605988, 1.954407, 1.000519, -5.936707, 
    -3.126831, 18.97057, 13.14272, -1.171097, -3.581757, 5.586716, 5.634109, 
    13.69089, -1.354172, 1.261978, -6.690887, 0.9801941, 2.7435, 2.900787, 
    -1.575775, -3.203644, -0.5638123, -2.873688, -3.255737, 2.317169,
  4.705475, 3.694519, 5.331512, 2.986206, 11.494, -0.2234344, 3.713028, 
    2.791656, -1.943222, -8.509125, -7.066406, -14.57135, -6.863281, 
    -0.6091156, 9.978119, 2.857834, -6.003922, -8.75885, -4.642456, 3.433594, 
    3.510956, 2.689087, 3.788269, 6.427612, 0.6442566, -4.169556, -5.248962, 
    0.848175, 0.1283875, -4.517456, -1.308319, -0.0604248, -0.3007813, 
    -6.742981, -16.45181, -23.7047, -11.0276, -23.64531, -28.92371, 
    -19.69218, -19.75131, -19.89973, -30.30367, -26.63463, -29.15208, 
    -21.54974, -28.4888, -33.93697, -20.71484, -9.1586, 1.231766, -13.50235, 
    -15.62032, -10.25728, -6.568237, -8.385651, -1.513794, -3.1875, 
    -6.951843, -8.606018, -3.940369, -11.83463, -13.42264, -11.90652, 
    -13.03256, -12.12057, -4.366928, 2.459122, 1.620056, 5.784637, 9.253632, 
    9.082031, 11.05026, 8.585938, -7.516663, -11.73697, 7.465881, 2.868492, 
    3.805481, 0.8216248, -1.648697, 5.851563, 8.412491, 11.29401, 10.90392, 
    -5.936203, -4.125519, -2.183838, -4.4422, -0.3932495, -2.805481, 
    2.680206, 6.23465, 6.591675, 5.888, 8.054962,
  7.00885, 4.874756, 2.261719, -0.3130188, 1, -8.802078, -6.010681, 1.764053, 
    3.796356, -7.980728, -14.5177, -17.02942, -11.44583, -8.054947, 
    -10.31952, -15.27655, -7.361465, -10.37422, -3.547668, 4.759369, 
    3.437256, -0.6695251, 0.2190247, 3.862, 5.5513, 3.190613, 0.5900879, 
    0.02032471, -1.332825, -0.3395996, -0.03878784, 3.458313, -2.60025, 
    -0.8973999, -1.759613, 0.651825, -3.1008, -18.57108, -9.068237, 
    -4.557816, -17.57057, -27.36458, -42.03697, -35.79897, -31.58514, 
    -29.97943, -32.0276, -33.67188, -27.06744, -15.22006, -8.248703, 
    -19.15964, -17.37761, -9.110153, -7.253387, -7.673691, -7.954956, 
    -8.405457, -4.264862, -2.54245, -1.363007, -2.716125, -2.832275, 
    -1.870575, -5.343475, -4.938538, 0.7664185, 1.677063, 6.852356, 9.377075, 
    13.25806, 9.868744, 9.345306, 0.9638062, -15.25989, -3.227341, 3.271873, 
    3.488281, -4.599243, 0.9093781, 5.431763, -6.395309, 8.561203, 17.57343, 
    19.63776, -5.952332, 5.507553, -3.669006, -4.251038, -1.485168, 
    -1.197144, -2.049469, 2.171356, 4.238281, 4.362762, 5.47525,
  -3.417694, -2.611725, -4.639313, -0.3934937, 4.628403, 4.110413, 6.259109, 
    6.241669, -7.887238, -26.00156, -36.97162, -23.34166, -18.03229, 
    -13.58592, -9.256775, -7.532806, -6.960159, -2.262497, 0.3986969, 
    1.349472, 4.461441, 3.027893, -0.9669189, 4.213287, 3.229706, 4.900269, 
    -2.588287, -3.599487, -1.912231, -5.083069, -6.877075, -9.71405, 
    -3.346619, -0.5447845, 10.22108, 5.746872, -19.69272, -6.494263, 
    6.286194, 3.726563, -16.47812, -17.8914, -20.58698, -19.10547, -21.78647, 
    -22.00989, -4.436981, -9.607025, -9.97345, -6.559113, -4.818756, 
    -4.162766, -0.6190186, -0.9466095, -4.310928, -8.904953, -8.273956, 
    -7.129425, -6.4263, -6.752609, -5.432816, -6.272156, -2.145325, 
    -4.136169, -3.442444, -7.4328, -4.942169, -6.313538, -3.091125, 
    -6.654144, 3.6539, -0.40625, -6.8685, -7.831238, -12.2901, -7.133591, 
    -5.478897, -1.549728, 10.84375, 6.566925, 11.67032, -1.619797, 2.975784, 
    13.1427, 3.367981, -3.816406, 10.36172, 4.019012, -0.1669006, -2.376038, 
    0.6047058, 1.121857, -0.5671997, -2.173431, -1.230713, -1.9039,
  0.3127441, 0.6968689, -0.8666687, 5.039322, 10.69922, 12.30339, 14.43437, 
    13.11693, 2.257813, -32.48073, -23.55652, -9.698456, -11.84506, 
    -6.603638, -5.605988, -1.84375, -3.52475, -3.598175, 0.7210999, 6.727081, 
    4.084106, 1.192719, -1.681519, -0.4023438, -0.971344, -1.36615, -6.5849, 
    2.261459, 0.3458405, -9.6026, -5.373703, -8.503647, -6.27343, -1.480728, 
    11.86667, 5.209106, -18.24557, -20.86772, -23.631, -18.90808, -11.019, 
    -10.18542, -3.760406, -3.272919, 7.419266, 7.035675, 13.55078, 14.49922, 
    12.39635, 15.11433, 15.58881, 13.39165, 13.74895, 13.30028, 6.339081, 
    1.132813, 1.325012, 2.054932, 0.2257996, -2.605988, -4.762756, -7.634369, 
    -8.720306, -9.835663, -8.66095, -5.380707, -8.572113, -4.716675, 
    -0.7799377, -5.179169, 1.88205, -5.365891, -9.542709, -11.41016, 
    -4.775787, 6.396881, -11.49557, -3.604691, -2.829941, -6.736969, 
    0.7755127, 3.130707, 8.281006, 16.7039, 10.67839, 0.7296753, 3.352875, 
    2.927338, 6.488281, 1.870056, 1.720856, 0.4380188, 0.5648499, 0.5315247, 
    0.9153748, -2.335938,
  -1.090363, -3.013, 0.3247375, 21.12421, 20.8802, 17.60027, 10.74452, 
    11.96225, 0.5945282, -17.44141, -13.52814, -6.273193, -5.052063, 
    -1.372406, -5.260925, -2.438019, -6.595825, -7.972137, -0.393219, 
    1.636475, 3.850769, -0.3494873, -0.8260498, 0.526825, -0.7533875, 
    -3.258331, -0.6888123, 9.56459, -7.898712, -7.096085, -1.740372, 
    -9.72084, -14.95755, -2.485428, 6.886978, 7.815887, -1.766922, -8.557297, 
    -3.184891, -2.604172, -3.962769, -2.11145, 1.72995, -0.1440125, 2.889587, 
    8.052856, 7.259644, 5.597107, 8.392456, 12.02316, 11.14896, 8.783081, 
    12.84219, 8.818481, 7.436737, 5.092712, 3.047638, -0.471344, 3.390106, 
    2.420319, 1.307526, -0.5872192, -1.728394, -4.153656, -5.058594, 
    -5.347382, -5.154694, -5.262238, -1.17865, -2.679413, -4.24765, 
    -3.989075, -15.94896, -13.55963, -8.822662, 5.233597, -14.31406, 
    -10.29245, -9.942169, -10.51041, 0.7950745, 7.8703, 16.50417, 7.504684, 
    6.6297, 8.227356, 8.4534, 5.210419, 3.035431, -0.3403625, 0.6028748, 
    -0.7773438, -2.279968, -3.111725, -2.39505, -4.170563,
  0.8768311, -1.385132, 8.400269, 9.737488, 5.719788, 10.08228, 8.455719, 
    0.9460754, -1.882813, -3.684357, -11.04323, -5.169525, -3.255737, 
    6.948425, -0.9158936, -1.907288, -0.8588562, -1.5867, -1.747925, 
    -0.4080811, -5.013031, -1.59375, 2.057007, 1.607025, 1.060944, -2.552856, 
    4.65625, -1.427094, -12.06302, -3.249756, -4.997925, -11.51172, 
    -14.39322, 0.5442657, 2.568497, 1.177353, 2.750519, 2.08699, 4.443222, 
    1.32135, 0.7221375, 4.025787, 2.228363, 3.197906, 0.7567749, 1.829956, 
    0.7088623, -0.3479004, -1.308594, -1.47345, -1.821609, -0.8653717, 
    -0.3005219, 2.501312, 5.091675, 9.372391, 12.01744, 15.65286, 8.609116, 
    11.84975, 9.214066, 10.83853, 5.329163, 6.016418, 4.744003, 1.974747, 
    1.60495, -0.04165649, 3.784912, 0.4721375, -1.550262, 4.099243, 
    -3.780975, -17.10052, -21.13126, -13.97369, -15.74219, -4.494507, 
    -7.44165, 11.37189, 11.13203, 6.722137, 3.152084, -2.431519, 0.1385498, 
    1.2836, 1.325256, -0.1927032, 1.383575, 2.304413, 0.7437439, -2.340363, 
    -3.814331, -0.3528748, 4.838287, 1.115082,
  -1.843506, -2.202087, 0.06381226, 1.083344, 0.2125244, 0.4794312, 0.153656, 
    -1.413818, -2.501312, -2.287231, -3.619797, -3.843475, -3.342468, 
    -0.651825, 9.199738, 5.139328, 9.410156, 2.460938, -0.07241821, 
    -4.373199, -4.903625, -4.949997, 0.1448059, 2.789063, -2.587524, 
    -2.605469, -4.325256, -5.774475, -2.798187, -3.322418, -6.366943, 
    -7.767715, -9.094788, -5.488022, -8.186447, -5.733856, 1.99765, 
    -1.161194, -1.306, 1.207031, 0.7984467, 1.474762, 1.286728, 3.517975, 
    2.883347, 4.845306, 6.137222, 5.864853, 5.286987, 6.232559, 5.027344, 
    7.640106, 1.905472, 3.255478, 5.891663, 6.093231, 9.75235, 12.50131, 
    11.46822, 12.04506, 9.904953, 13.82787, 12.94557, 12.77162, 12.73334, 
    7.988281, 9.791916, 6.087769, 4.654968, 7.201569, 2.620819, -6.39325, 
    -11.25937, -7.887238, -4.882813, 0.9026031, 12.38438, 5.67421, 4.796082, 
    5.225006, -4.931519, -4.027603, -7.711716, -4.337234, 0.382019, 
    -0.045578, 0.9630127, 5.625778, 3.190094, 1.617706, -1.808075, -3.235687, 
    -3.483337, -0.5617371, 0.8153687, -2.012482,
  0.3825378, 0.5856934, 0.1244812, 0.5778503, -0.5632629, -0.5734253, 
    -1.070038, -0.6195374, -2.880219, -4.003906, -2.692719, -3.839081, 
    -3.005219, 0.03384399, 10.01563, 3.70755, 14.01537, 9.565643, -2.510162, 
    -9.10025, -5.889587, 4.13829, -8.247681, -5.748169, -2.776031, -2.875, 
    -4.713531, 5.110947, 10.78125, -0.8541718, -3.139847, -5.041153, 
    -4.173187, -7.670044, -4.463013, -0.9015656, -0.6828156, -1.644791, 
    2.628387, -1.001556, -0.4098816, -1.50676, -1.478638, -0.478653, 
    0.735672, 4.21405, 1.787506, 5.534637, 1.34375, 6.51329, 8.404953, 
    10.29271, 11.26094, 9.078125, 9.648438, 8.570831, 11.75052, 11.70103, 
    9.866928, 11.22136, 12.30937, 9.009628, 9.642975, 12.41484, 14.37109, 
    13.4073, 9.956772, 10.85339, 6.762497, 2.741394, -0.775238, -7.74115, 
    -6.596603, 11.47058, 4.230988, -4.670303, -5.44165, -6.53801, -2.753906, 
    -6.980988, -6.346878, -0.0945282, 2.429169, 1.446106, -2.411194, 5.06926, 
    3.899216, 3.410416, 3.6073, 2.523956, 1.319794, -0.06719971, 0.9283752, 
    2.409637, 1.534882, 0.6497192,
  2.739594, 2.536194, 2.025543, 2.501556, 0.6528625, 0.7320251, 0.06848145, 
    0.5583496, -0.1669312, -3.319, -3.846375, -3.097656, -2.590607, 
    -2.228668, -0.4390564, 2.718735, 2.009109, -0.3721313, -0.2484436, 
    -4.997925, -10.76511, -1.755997, -5.254425, -6.858826, -9.35675, 
    -1.997131, -2.263275, 3.333847, 8.396088, -8.2276, -3.604431, -7.497406, 
    -2.351288, -13.21198, -8.589066, -4.416397, -0.589325, 0.2841187, 
    -1.791931, -1.576294, 1.264587, -1.488022, -3.922134, -5.880219, 
    -1.532043, 5.371353, 5.953903, 4.08046, 3.797653, 4.017441, 4.97995, 
    8.353119, 5.028122, 9.396088, 5.266144, 5.998444, 4.638031, 7.342194, 
    6.289841, 7.346863, 9.149734, 9.023178, 14.84167, 14.98412, 21.28725, 
    15.69141, 12.67162, 10.23151, 5.380737, 12.70207, 8.754684, 15.67578, 
    14.8, 5.141159, -6.700256, -4.290359, -5.905212, -9.289856, -5.400009, 
    -0.9406281, -3.854172, -5.260941, -0.8322906, 1.828644, 3.107025, 
    5.383072, 5.087234, 7.216141, 6.118744, 1.731262, 0.225769, 1.833588, 
    0.5770874, 2.016144, 4.330963, 2.603638,
  3.736481, 3.341675, 0.8023376, 1.235657, 3.717438, 3.439056, 2.184906, 
    -0.6374817, 0.4510193, -0.9437561, 3.004944, -0.3830872, -3.310699, 
    -3.925262, -0.5783997, 1.481247, 3.509903, -1.77005, -2.888275, 
    -3.385406, -8.097137, -10.58723, -8.207275, -7.311981, -6.127838, 
    -5.100525, -12.63177, -16.41797, -10.54271, -0.7450562, 2.323166, 
    -5.074478, -2.516144, -2.137756, -5.018219, -5.837494, -8.224487, 
    -2.113281, 1.474991, 1.591934, 1.14949, -0.3874969, 0.2773438, -1.048965, 
    -1.763275, 1.439575, 3.659119, 2.008331, 8.357544, 4.465363, 4.296097, 
    10.54973, 3.55574, 3.303909, 1.680206, 4.620316, 5.169525, 3.987503, 
    3.166931, 0.3692627, 2.533585, 3.598434, 9.125259, 10.41615, 12.48151, 
    9.640106, 10.25833, 9.116928, 9.946869, 21.47266, 17.675, 14.28125, 
    6.603653, 2.314316, 2.429428, -1.130981, -3.655212, -7, -8.671875, 
    -10.63387, -7.900009, -11.41953, -2.93074, -4.123962, -1.12709, 1.736969, 
    2.870834, 9.115372, 7.316406, 3.339066, -2.931503, -1.093994, 2.065094, 
    -0.7059937, 1.421875, 2.479431,
  1.596359, 2.645828, 3.999741, 3.228119, 0.6567688, 2.573181, 4.385941, 
    3.360672, 0.8083344, 0.7731781, 0.8359375, -0.4101563, -1.778915, 
    0.6708374, 2.047653, 0.9255219, 6.082825, 1.8862, -0.625, -1.329941, 
    -3.124466, -5.582031, -4.483337, -4.694016, -6.2724, -6.530731, 
    -5.731506, -16.11902, -25.07396, -7.674484, 0.5562515, 4.226303, 
    0.8070374, 3.039581, 9.212494, 6.687241, 5.521881, -0.9294281, -1.783325, 
    -4.294266, -4.288284, -1.259109, -2.431503, 0.3119812, -0.5703125, 
    4.443497, 2.309891, 4.24115, 1.206512, -0.7395782, 5.283081, 6.543228, 
    6.348175, 3.780212, 0.6023407, 4.127869, 3.86824, -1.370316, 0.7958374, 
    -3.274216, 1.304947, -0.3033905, 6.759628, 6.980469, 10.07031, 6.59584, 
    5.947403, 9.550781, 12.3138, 22.58514, 13.03673, -0.1799469, 0.5502625, 
    1.226303, 0.6398468, 0.1419373, -5.101563, -4.750259, -4.223434, 
    -4.941147, -8.373444, -3.36824, -2.479172, -6.450256, -0.610672, 
    -1.402344, -0.7427063, 1.137238, 3.447922, 6.92421, -0.3197937, 
    -0.3734283, 0.3312531, -0.6276093, -0.2046967, 0.7742157,
  -0.3096313, 0.377594, 3.015091, 2.31485, 2.650253, 4.774216, 5.3974, 
    5.061966, 1.91954, 4.67865, 6.104691, 1.749222, 1.925262, 4.9599, 
    9.574478, 9.918747, 16.27109, 14.16328, 7.401825, 6.32605, 2.128128, 
    0.190094, -2.516678, -1.878387, -4.340363, -21.74532, -7.084885, 
    -16.7323, -25.13724, -14.03568, -0.6945343, -3.865623, 3.253387, 
    2.550522, 10.75339, 5.493484, 9.555466, 10.2263, 10.38853, 6.864853, 
    0.1822815, -0.9289093, -4.424728, -0.441925, 3.694794, 6.963287, 
    3.795837, 5.598969, 3.877609, 4.795578, 4.586975, 2.387772, 5.233063, 
    5.63855, 4.028381, 4.676559, 0.6091156, 0.2010345, -1.585159, 0.1140594, 
    -2.119781, 0.7179718, 4.424225, 7.449478, 3.534378, 4.039063, 8.699219, 
    12.42682, 14.24896, 10.99532, 11.67606, 7.264313, 4.197922, 3.97995, 
    2.326309, -1.205994, -1.48204, -4.241135, -3.602615, -5.377853, 
    -4.319534, -5.807037, -6.706512, -2.385681, -0.2502594, -0.4315033, 
    -3.119278, 1.55365, 4.215363, 3.25209, 4.113541, 2.853134, 3.492447, 
    1.740875, 1.032028, -0.08306885,
  5.152863, 4.695313, 4.308334, 3.203644, 3.319275, 2.703384, 7.997131, 
    9.004684, 5.205719, 13.57526, 13.90677, 9.787231, 5.496872, 9.282806, 
    12.08073, 9.671616, 7.698441, 12.92421, 22.03777, 12.20547, 7.35704, 
    -3.930725, -2.471619, -3.222916, -1.869522, -3.110413, -3.761459, 
    -8.266144, -17.11615, -11.50469, -7.436188, -12.58281, -12.91251, 
    -1.044266, 0.9802094, 5.020309, 1.184113, 5.807297, 8.647911, 3.349998, 
    5.409119, 3.967194, 3.137497, 6.679428, 6.294266, 1.133591, -1.936447, 
    -0.9455719, -1.983337, 0.2023468, 1.406769, 2.169022, 5.726044, 4.907562, 
    -0.06459045, -1.535156, -2.787491, -2.245056, -2.143494, 0.09532166, 
    0.5690155, 2.544266, 8.303131, 7.09166, 4.295563, 5.204163, 9.75885, 
    11.57864, 12.04869, 9.416138, 6.825256, 3.92865, 1.201035, 3.872391, 
    4.224487, -2.915894, 0.7239532, -0.5195313, 0.3010406, 0.8367157, 
    1.130203, 0.6273499, 1.058594, -1.7612, -0.9059906, -1.492981, -1.416153, 
    -0.0942688, 3.045044, 0.8872375, 4.305222, 2.883331, 6.020569, 6.251297, 
    13.90443, 13.99687,
  16.94766, 17.82812, 17.82083, 13.25052, 4.438797, 1.83255, 7.12291, 
    9.169525, 13.14949, 14.18282, 18.53515, 13.9711, 13.43933, 5.844009, 
    4.104691, 1.302597, 0.2427063, 0.1500092, 1.777603, 0.0406189, -4.032043, 
    -2.447144, -2.873184, -4.064835, -8.334106, -4.450272, -4.367966, 
    -1.193481, -8.22084, -2.278122, -1.723694, -5.515106, -8.04895, 
    -6.668488, -11.31667, -5.932556, -4.49427, -8.913803, -1.755722, 
    -1.409378, -2.155731, 1.422653, 0.3161469, -0.8440094, -0.454689, 
    0.1572952, -4.66172, -3.097397, -1.157288, -1.636719, -4.530464, 
    -5.735672, -0.5125046, -0.752861, -4.167961, -3.545822, -3.065613, 
    2.071609, -1.265099, -0.1890564, 2.03334, 0.3453064, 1.707809, 6.665634, 
    9.488281, 5.488541, 3.5401, -2.6922, -0.8859253, 1.239319, 1.459641, 
    -0.7692566, -2.001831, -3.406509, -0.3838577, 1.119003, -0.02786255, 
    -0.02812195, -0.7932358, 1.402603, 4.886719, 2.675781, 0.01483917, 
    -3.560944, -0.7825546, -0.9637985, -5.124733, -2.289841, -3.47213, 
    -4.957809, -0.8862, -1.048172, 2.5625, 5.609116, 10.52292, 15.38203,
  8.064064, 6.730988, 7.577087, 8.408333, 3.261971, 7.665359, 4.524475, 
    3.465363, 5.218231, 4.135674, 4.879692, -3.809898, -4.604172, 0.6679688, 
    -0.05807495, -5.148697, -7.344528, -6.542969, -7.064331, -2.719803, 
    -4.5513, -8.474991, -6.666153, -3.809891, -4.707031, -4.297653, 
    -6.181244, -2.485168, -2.199478, -3.656525, -1.987503, -1.958069, 
    -2.771103, -4.603912, -7.68985, -2.348434, -1.623955, -11.23307, 
    -5.646355, -4.621613, -6.34687, -4.089325, -1.195839, -5.852867, 
    -5.625786, -3.465103, -3.910934, -6.148438, -2.650002, -2.479431, 
    -3.032028, -2.351303, -1.887497, -6.289848, -7.387756, -5.058594, 
    -4.066406, -3.669533, -0.984375, -1.144272, 0.467186, 2.177605, 7.481773, 
    6.686455, 3.854683, -5.56015, -7.977089, -9.496094, -7.692459, -5.473953, 
    -7.616409, -9.818748, -9.403648, -11.37579, -9.285156, -12.24635, 
    -7.518234, -0.3156281, 0.5752563, 2.274742, -0.3799515, 1.122658, 
    5.023956, 3.898956, 2.11615, -0.2781296, -6.125, -4.945831, -4.739326, 
    -2.435936, -3.328392, -6.289063, -2.837242, 0.5927048, 7.084641, 10.04297,
  -3.147133, 1.072395, 1.189842, -1.045578, -0.3065109, -0.9416733, 
    -10.31719, -6.37162, -4.057289, -7.021088, -5.445572, -5.143753, 
    -6.657288, -2.13047, -7.136978, -12.59714, -14.47812, -15.99583, 
    -10.88126, -7.006775, -6.74453, -7.739586, -4.785675, -5.765884, -3.8349, 
    -3.413284, -5.251556, -3.827072, -2.067459, -2.22084, -0.7098999, 
    -1.845062, -2.50209, -2.686462, -5.505219, -3.874481, -1.326302, 
    -3.828903, -6.603386, -6.385422, -7.52813, -3.986458, -1.888802, 
    -1.652344, 1.880203, -0.3140564, -3.24765, -3.365623, -2.653122, 
    -2.490883, -3.404686, -4.813545, -3.089058, -1.396095, -4.648178, 
    -4.500259, -4.610161, -5.772392, -0.9473953, -0.5690155, -2.712753, 
    0.07395935, 3.89505, 6.044014, -3.891151, -6.082031, -3.213806, 
    -5.463799, -7.591148, -7.208336, -10.38776, -12.31693, -11.12135, 
    -13.33151, -13.525, -10.75651, -9.657036, -10.09792, -8.091141, 
    -2.923691, -2.303642, 1.713539, 5.333076, 1.438805, -0.3445358, 
    0.3372421, -0.5385361, -0.9950562, -4.54583, -5.540108, -3.903648, 
    -1.819794, -1.210938, -0.5859375, 3.558334, 2.32943,
  -4.082291, -4.3013, -9.055729, -7.670052, -5.680466, -6.526566, -7.157028, 
    -4.001556, -6.72422, -12.82994, -9.674477, -10.70703, -9.57917, 
    -7.458076, -9.200783, -11.05598, -6.72213, -5.414589, -6.360939, 
    -6.179169, -8.379425, -7.697914, -5.489319, -6.747917, -7.455208, 
    -6.394791, -6.006767, -3.238022, -2.821617, -4.302345, -6.264328, 
    -6.980728, -5.249481, -4.852348, -7.460938, -3.737503, -1.322395, 
    -2.641411, -1.462761, -3.925522, -0.4791641, -0.5208282, -4.242966, 
    -4.368752, 0.9562531, -1.439323, -5.507027, -2.652863, -0.735939, 
    -0.1236954, 1.61068, -1.500259, -2.886459, -0.7005157, -2.541405, 
    -3.194016, -2.480209, -2.304169, 0.6328125, 1.907547, 1.603912, 4.537758, 
    5.025002, 0.5026054, -3.023174, 2.052864, -0.390625, -2.936974, 
    -6.730728, -6.659897, -7.658859, -7.402603, -8.348701, -18.51224, 
    -9.580986, -7.488541, -7.030205, -7.466927, -5.859375, -6.579689, 
    -3.221092, -0.2286453, 1.02787, 1.284378, 2.112762, 3.471878, 2.484642, 
    1.782028, 0.1114578, -1.771355, -0.623436, 0.3947906, -2.967186, -1.6987, 
    -0.7479172, -3.317707,
  -6.09375, -7.007813, -9.982555, -10.23776, -9.853645, -10.13203, -8.231251, 
    -7.041924, -9.644012, -8.058075, -6.560677, -10.84714, -11.32161, 
    -7.333328, -5.885933, -9.148697, -9.322914, -4.854431, -5.611984, 
    -4.467972, -5.154686, -8.410416, -7.704163, -7.776817, -6.67318, 
    -5.870316, -5.872917, -7.559113, -9.871613, -7.148178, -6.596619, 
    -5.867188, -6.602348, -5.416931, -5.445831, -5.568489, -4.235939, 
    -0.1151047, -7.612762, -20.03958, -12.82031, -6.697132, -3.813805, 
    -2.628387, -0.7992249, -2.108337, -1.2388, 1.27969, -0.4205704, 
    -3.589325, -1.589844, 0.1348953, 0.09296417, 0.08724213, -0.2984352, 
    0.1591148, 0.4557266, 1.140099, 0.4481812, -0.6283836, 1.105209, 
    1.789845, -0.03620148, -3.060677, -2.636459, -1.824219, -4.647919, 
    -2.079689, -1.379951, -4.482033, -3.688545, -4.192451, -4.59037, 
    -4.605995, -6.121613, -5.240623, -9.688805, -10.59166, -6.724739, 
    -2.5849, -2.644005, -2.511719, -4.8638, 0.2283821, -0.6580696, 1.357811, 
    3.134636, 4.605988, 2.461197, 0.3216133, -2.234116, -2.539322, 
    -0.9528656, -2.625263, -4.548962, -5.711979,
  -3.097656, -3.755989, -5.740623, -7.753124, -7.298958, -7.273956, 
    -5.121094, -6.987499, -8.626564, -7.108593, -3.397137, -3.98724, 
    -5.144012, -6.594269, -8.999218, -11.15911, -8.024738, -6.601818, 
    -8.879425, -8.652081, -3.455727, -3.455727, -5.523956, -6.314323, 
    -6.686977, -6.106247, -5.483856, -5.311718, -6.309635, -8.403126, 
    -7.309895, -7.025002, -7.701042, -6.024994, -4.862495, -5.023178, 
    -3.939583, -4.273438, -11.65885, -21.75625, -18.21875, -9.69323, -3, 
    -1.448959, 0.5583344, -0.7317696, -2.642971, -1.473698, -1.327343, 
    0.1421852, -0.2322922, -0.5296898, -1.502083, -1.947918, -1.438545, 
    -3.047138, -2.223175, 1.342709, 1.43177, 1.609898, -0.8729172, -4.851563, 
    -3.878124, -2.648438, -1.964844, -3.791927, -1.728645, -0.6513023, 
    0.8304672, -0.6041679, -0.5911446, -1.25, -2.972397, -6.920055, 
    -7.011196, -10.89896, -10.48672, -8.364326, -6.052082, -6.816143, 
    -7.059372, -13.0612, -9.988022, -3.221352, -0.9406242, 0.6091156, 
    0.8557281, 0.5294266, 1.496616, 1.194012, -0.9869804, -0.967186, 
    -0.1028633, -1.788021, -2.351303, -2.780991,
  -2.755211, -3.574741, -5.519531, -5.865103, -4.201824, -2.031513, 
    -2.695049, -2.266666, -3.060677, -3.799477, -3.189842, -2.963543, 
    -3.871616, -4.254688, -6.773701, -4.667969, -3.444271, -5.090103, 
    -6.02005, -6.502605, -6.982292, -5.91198, -5.706249, -3.527866, -2.51823, 
    -5.50729, -6.108334, -3.519272, -2.260159, -5.087502, -6.983334, 
    -5.767967, -5.134377, -4.248699, -5.373177, -3.867447, -4.234894, 
    -5.608852, -10.17786, -13.53464, -13.09661, -8.489323, -5.030727, 
    -2.191666, -3.347397, -0.7250004, -1.691406, -2.732811, -4.140362, 
    -3.114323, -1.405731, -1.691666, -3.167446, -1.527866, -2.560158, 
    -2.638542, -3.431774, -3.165886, -1.976299, -2.837761, -5.437761, 
    -4.969271, -4.06823, -2.076305, -3.036198, -1.620312, -0.5677109, 
    -0.1778641, -2.072136, -1.34375, -1.182552, -1.809895, -3.424999, 
    -4.376823, -5.856251, -7.344528, -7.771618, -6.008072, -4.121876, 
    -5.655991, -9.53828, -11.93255, -7.565365, -1.752865, 0.6500015, 
    1.372917, 0.188282, -0.3997383, -0.5013008, -1.31953, -1.159634, 
    -2.707031, -2.622654, -2.669529, -2.53828, -2.16823,
  -1.957291, -2.625523, -1.704428, -1.371355, -0.994791, -2.854948, 
    -0.3760433, -0.1036453, 0.4619789, -0.08437538, -1.297398, -2.638802, 
    -2.246614, -2.07526, -2.604687, -2.505468, -2.961458, -4.641928, 
    -2.430988, -0.124218, -1.811718, -4.562759, -4.774479, -2.357031, 
    -2.339062, -4.056252, -4.696354, -2.906511, -1.411457, -2.693748, 
    -4.20755, -4.008852, -4.04401, -3.73177, -4.208332, -5.088541, -4.350262, 
    -4.513542, -5.778385, -6.60677, -6.515886, -5.879948, -4.432032, 
    -3.550259, -2.210155, -2.948698, -7.046616, -11.78125, -11.64818, 
    -11.58073, -11.76614, -9.608335, -5.252346, -3.181772, -3.126562, 
    -3.839064, -3.276302, -4.335676, -5.735678, -6.235416, -5.237501, 
    -3.504427, -0.5856762, 0.1273441, 0.767189, 0.3111992, -0.9372387, 
    -2.134113, -2.669271, -1.920572, -1.327866, -2.805729, -4.191147, 
    -5.308075, -5.387497, -5.964062, -5.999737, -6.138542, -5.403908, 
    -5.285156, -5.293491, -4.25703, -1.776825, -0.8789063, -1.139322, 
    -0.2265625, 0.9122391, 0.7729168, -0.1567707, -1.497656, -1.747656, 
    -0.1927071, 1.453125, 1.016407, -0.5406246, -1.29479,
  0.36901, 0.5205727, 0.04296875, -1.193749, -1.244532, -0.8252602, 
    -1.860937, -1.248959, -1.183332, -0.4364586, -0.1484375, -0.4710932, 
    -1.447395, -1.401563, -1.210938, -1.554428, -2.63724, -3.461719, 
    -3.347397, -3.370313, -3.100782, -2.937239, -1.876561, -1.147917, 
    -1.455729, -2.413021, -2.75651, -1.857031, -1.548178, -2.676563, 
    -3.126562, -2.872395, -2.237499, -1.889063, -3.006771, -3.89974, 
    -4.193228, -3.979427, -4.356251, -4.758072, -4.691406, -4.014845, 
    -3.792707, -3.094271, -2.926043, -2.647657, -2.664324, -2.938021, 
    -2.36849, -2.030729, -1.870573, -2.350521, -2.268749, -2.396093, 
    -2.079687, -2.031771, -2.698698, -3.239323, -3.63229, -3.008074, 
    -1.957552, -1.625521, -1.801041, -1.7125, -1.243229, -1.039324, 
    -1.590364, -1.994793, -2.170053, -1.739325, -1.411198, -1.355728, 
    -2.467709, -3.654947, -3.609896, -3.478386, -3.195833, -2.983072, 
    -2.370834, -2.284636, -2.1625, -1.357552, -0.645052, -0.5815105, 
    -0.3070316, 0.09114647, 0.4401045, 0.8544273, 1.326302, 0.4221354, 
    -0.5778646, -0.3830729, -0.2059898, -1.064583, -1.674999, -0.714323,
  0.8911462, 1.008594, 0.7992187, 0.7166672, 0.6463537, 0.8497396, 0.6216149, 
    0.08307266, -0.3572917, -0.4981775, -0.625782, -1.759896, -1.834114, 
    -1.82448, -1.815104, -1.752604, -1.654427, -1.611198, -1.702084, 
    -1.579688, -1.453906, -1.729688, -1.704948, -1.752344, -2.119532, 
    -2.341927, -2.120573, -1.877604, -1.760417, -1.932291, -2.171354, 
    -2.366927, -1.950781, -1.648698, -1.433073, -1.596093, -2.315886, 
    -2.761979, -3.099219, -2.907552, -3.208334, -3.547916, -3.637501, 
    -3.423178, -3.132813, -2.720053, -2.697396, -2.672396, -2.925261, 
    -3.309375, -3.427865, -3.189063, -3.141147, -2.676042, -2.390365, 
    -2.294532, -2.507552, -2.39349, -1.912761, -1.221354, -1.003646, 
    -1.020573, -1.321094, -1.842187, -1.332031, -0.6648436, -0.6973953, 
    -0.759635, -1.414063, -2.05, -1.96849, -1.936458, -2.107291, -2.465103, 
    -2.275521, -2.684114, -2.403125, -2.338802, -2.313021, -1.679688, 
    -0.5859375, -0.2213535, 0.02057362, -0.3312502, -1.051042, -0.953125, 
    -0.2385416, 0.5028639, 0.4721355, 0.5486984, -0.0348959, -1.821355, 
    -2.388021, -1.503646, -0.2328129, 0.2114582,
  -0.0703125, -0.03932309, 0.06875014, 0.263021, 0.4020832, 0.5221355, 
    0.3632813, 0.1377606, -0.1945312, -0.5239584, -0.9221354, -1.03099, 
    -1.136458, -1.061198, -1.005469, -0.8966148, -1.007031, -1.113021, 
    -1.202083, -0.8976562, -0.8630211, -0.9476562, -1.175781, -1.192188, 
    -1.165104, -1.172136, -1.074739, -1.046354, -0.9861979, -1.075521, 
    -1.146875, -1.148698, -1.280469, -1.328646, -1.379948, -1.43776, 
    -1.408333, -1.464323, -1.4125, -1.315625, -1.383333, -1.607292, 
    -1.811458, -1.990104, -2.057552, -1.932292, -1.605469, -1.418229, 
    -1.255729, -1.234375, -1.262761, -1.260156, -1.295052, -1.180729, 
    -0.9270835, -0.8658857, -0.8945313, -0.8153644, -0.7901044, -0.7835937, 
    -0.7809896, -0.734375, -0.9825521, -1.088802, -1.067188, -0.8736982, 
    -0.7981772, -0.9276042, -1.054167, -1.290625, -1.170834, -1.168489, 
    -1.252604, -1.205469, -1.146875, -1.013802, -0.8479166, -0.7841144, 
    -0.7713542, -0.5111976, -0.1705732, 0.04374981, 0.1171875, -0.03984404, 
    -0.3294272, -0.6382813, -0.6156249, -0.511198, -0.4195313, -0.4734378, 
    -0.4440103, -0.3283854, -0.578125, -0.7955728, -0.7757812, -0.3200521,
  -0.03281248, -0.01640624, 0.03177083, 0.01041663, 0.001302063, -0.09062499, 
    -0.2432292, -0.3312501, -0.3515626, -0.3143229, -0.3304687, -0.2255208, 
    -0.1312499, -0.1510416, -0.1877605, -0.2919271, -0.4098959, -0.4447916, 
    -0.4333333, -0.4630208, -0.4791667, -0.4007813, -0.2622396, -0.2773437, 
    -0.2726563, -0.2776042, -0.2802083, -0.2309896, -0.2044271, -0.2052084, 
    -0.2044271, -0.2533854, -0.2945312, -0.3447917, -0.3653646, -0.3973958, 
    -0.4299479, -0.4822917, -0.4921875, -0.3885417, -0.3239584, -0.3710938, 
    -0.3911459, -0.4125, -0.3885416, -0.3653646, -0.3802083, -0.3552084, 
    -0.3132813, -0.3419271, -0.3752604, -0.3927083, -0.3934896, -0.4242188, 
    -0.4356771, -0.3848958, -0.334375, -0.2638022, -0.179948, -0.2085937, 
    -0.2450521, -0.2338542, -0.2398437, -0.2393229, -0.2174479, -0.1354166, 
    -0.145573, -0.1924479, -0.2403647, -0.273698, -0.3075521, -0.3166667, 
    -0.309375, -0.3229167, -0.3322917, -0.3406249, -0.2385417, -0.1346354, 
    -0.05989587, -0.05703115, -0.07994795, -0.07630217, -0.0533855, 
    -0.05442715, -0.0958333, -0.1460937, -0.1505209, -0.1666667, -0.1583333, 
    -0.1359375, -0.09713542, -0.0226562, -0.02083337, -0.02734375, 
    -0.06874996, -0.06848961,
  -0.02109375, -0.02083334, -0.01796875, -0.01640625, -0.009375002, 
    -0.002343748, 0.004427083, 0.008072913, 0.004947916, 0.002083331, 0, 
    -0.009635419, -0.01901042, -0.02838542, -0.03463542, -0.03828125, 
    -0.03932292, -0.03567708, -0.02578125, -0.01640625, -0.009635411, 
    -0.007291667, -0.005729169, -0.00807292, -0.01406249, -0.01484375, 
    -0.01979167, -0.025, -0.028125, -0.025, -0.025, -0.01927083, -0.01822916, 
    -0.01458333, -0.01770833, -0.02317708, -0.02473959, -0.02838542, 
    -0.02421875, -0.021875, -0.021875, -0.02109375, -0.01692709, -0.015625, 
    -0.02005209, -0.01927083, -0.01744791, -0.01848958, -0.02057292, 
    -0.01822916, -0.01223958, -0.0125, -0.01510417, -0.01692709, -0.02109375, 
    -0.01510416, -0.01875, -0.01848958, -0.01770833, -0.02161458, 
    -0.02161458, -0.02786459, -0.02942708, -0.02838542, -0.03385416, 
    -0.03098958, -0.02083334, -0.01614583, -0.01223958, -0.00755208, 
    -0.01171875, -0.008854166, -0.008333333, -0.01276042, -0.0171875, 
    -0.01901042, -0.02135416, -0.01979167, -0.02265625, -0.01953125, 
    -0.01901042, -0.02057292, -0.01614583, -0.01041667, -0.007031254, 
    -0.004947916, -0.004166663, -0.007031247, -0.007291667, -0.002864584, 
    -0.005729169, 0.0002604201, -0.002604172, -0.01302084, -0.01640625, 
    -0.02135416,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -1.861547, -1.736025, -1.659201, -1.638109, -1.648264, -1.727171, 
    -1.815453, -1.887068, -1.969097, -2.027952, -2.152693, -2.266493, 
    -2.327951, -2.382118, -2.466234, -2.566494, -2.679255, -2.766754, 
    -2.86936, -2.973785, -3.125347, -3.276911, -3.424305, -3.546181, 
    -3.678734, -3.813629, -3.909203, -4.028994, -4.053734, -4.066233, 
    -4.098524, -4.112329, -4.095661, -4.074306, -4.044098, -4.046701, 
    -4.033421, -4.068838, -4.131598, -4.120401, -4.07066, -4.002434, 
    -3.953213, -3.895922, -3.865454, -3.857901, -3.852431, -3.816234, 
    -3.757119, -3.680557, -3.629516, -3.548786, -3.406076, -3.226389, 
    -2.982638, -2.707379, -2.441234, -2.190451, -1.986805, -1.803733, 
    -1.642015, -1.531338, -1.440972, -1.323784, -1.232378, -1.15712, 
    -1.05113, -1.000349, -0.9782124, -0.9815979, -1.036024, -1.031076, 
    -1.067797, -1.130556, -1.140972, -1.222744, -1.363108, -1.519619, 
    -1.643576, -1.80842, -2.056858, -2.224045, -2.411024, -2.563889, 
    -2.685764, -2.790972, -2.762327, -2.752171, -2.711546, -2.667536, 
    -2.603994, -2.508421, -2.42066, -2.317795, -2.206078, -2.034721,
  -2.436283, -2.123001, -1.736019, -1.424824, -1.367794, -1.446438, 
    -1.640186, -1.838104, -2.049824, -2.260239, -2.462585, -2.638889, 
    -2.674297, -2.612835, -2.458931, -2.253723, -2.101898, -1.96492, 
    -1.892265, -1.976379, -2.156586, -2.417267, -2.742786, -2.99044, 
    -3.167786, -3.276382, -3.4631, -3.616745, -3.819088, -3.910236, 
    -3.905029, -4.043571, -4.289928, -4.654251, -4.922218, -5.125866, 
    -5.383678, -5.50477, -5.621958, -5.570913, -5.660236, -5.624041, 
    -5.487064, -5.468056, -5.261806, -4.953733, -4.785244, -4.741755, 
    -4.617796, -4.447224, -4.258421, -3.780035, -3.50712, -3.109722, 
    -2.742796, -2.424566, -2.105558, -1.888632, -1.824047, -1.676651, 
    -1.359983, -1.118578, -1.148525, -1.175348, -1.168318, -1.417017, 
    -1.600349, -1.574566, -1.406336, -1.36936, -1.490713, -2.024565, 
    -2.406855, -2.662066, -2.787846, -2.982901, -2.997744, -2.921963, 
    -2.775864, -2.637585, -2.594093, -2.559458, -2.487583, -2.524042, 
    -2.703207, -3.033415, -3.233414, -3.435759, -3.687061, -3.885498, 
    -3.858936, -3.618311, -3.389666, -3.121696, -2.834721, -2.643051,
  -2.455555, -2.520138, -2.763885, -2.961544, -3.176388, -3.356068, 
    -3.276642, -2.98941, -2.848526, -2.566235, -2.073006, -1.756599, 
    -1.747486, -2.036549, -2.469883, -2.902695, -3.074829, -3.076653, 
    -2.982903, -2.819359, -2.58004, -2.306599, -2.224567, -2.229778, 
    -2.644882, -3.213371, -3.816235, -4.237846, -4.711285, -4.8316, 
    -4.598267, -3.96936, -3.650093, -3.927952, -4.110504, -4.367798, 
    -4.440453, -4.473267, -4.68108, -5.378983, -6.18185, -6.851646, 
    -6.862846, -6.49305, -6.349819, -7.022736, -7.467529, -7.511801, 
    -6.87925, -6.326645, -5.690187, -5.138626, -4.332375, -3.12925, 
    -2.029253, -1.766752, -1.737585, -1.97118, -2.311024, -2.208414, 
    -1.674301, -1.237844, -1.355032, -1.547216, -1.919611, -2.234455, 
    -2.741226, -3.308416, -3.639404, -4.320915, -4.463886, -4.796432, 
    -5.237316, -5.786026, -5.388889, -5.272484, -4.836025, -4.356075, 
    -4.388889, -4.491486, -4.864403, -5.057114, -4.884716, -4.314926, 
    -3.782635, -3.050079, -2.278984, -1.342007, -0.3912277, -0.1201324, 
    -0.08185196, -0.6506004, -1.503204, -2.148262, -2.312325, -2.538368,
  0.1066895, 0.03636932, -0.8456726, -1.603462, -2.10321, -2.418312, 
    -2.20295, -1.723259, -1.668579, -2.399834, -3.249313, -3.478737, 
    -3.136543, -3.225868, -3.781593, -4.508942, -4.874313, -5.214149, 
    -5.73317, -6.688629, -7.054001, -6.808685, -5.666496, -4.622231, 
    -3.681862, -3.084465, -2.676125, -2.416229, -2.545662, -2.475883, 
    -2.90374, -3.524063, -3.655045, -3.552437, -3.230827, -2.980827, 
    -3.172501, -4.043854, -4.505051, -4.495941, -4.682396, -4.970398, 
    -5.116486, -4.799309, -4.566502, -5.168839, -6.645409, -8.405556, 
    -9.217793, -8.200348, -6.500599, -5.593567, -4.712578, -3.363628, 
    -2.1842, -1.629253, -1.818836, -0.7138824, -0.2315941, -0.4409714, 
    -0.8610191, -1.895912, -2.702164, -3.485241, -5.479771, -6.976646, 
    -6.957638, -6.831081, -7.114674, -7.158413, -6.866489, -6.63628, 
    -6.159981, -5.434975, -4.828728, -5.156071, -5.084461, -4.605549, 
    -4.397221, -4.73941, -5.466492, -6.215973, -6.711025, -6.833683, 
    -5.579517, -4.293839, -3.390453, -1.885769, -0.5909729, 0.7793388, 
    1.037937, 0.6644936, 0.7480888, 0.8184013, 0.1538086, -0.02170563,
  0.5543289, 0.8077164, -0.05973053, -0.1732788, 0.2189102, 1.805367, 
    2.236099, 2.985588, 3.221008, 1.468132, -0.9389038, -2.63343, -3.773796, 
    -3.745934, -2.955826, -2.060501, -1.896965, -1.913109, -2.654785, 
    -3.373543, -4.565994, -4.649841, -4.112083, -4.048279, -3.089684, 
    -2.300087, -2.103737, -2.816238, -3.621445, -3.76519, -3.96936, 
    -5.512589, -5.857384, -5.147224, -4.571182, -5.011803, -4.996445, 
    -3.817017, -3.035767, -3.2342, -2.931602, -2.759201, -1.888107, 
    -1.105827, -0.6308289, -0.1214294, -0.585762, -2.314423, -1.581341, 
    -0.1865463, -0.3886299, -0.9662361, -1.396706, -2.177952, -2.46492, 
    -2.344101, -2.171444, -4.184986, -4.746185, -4.900871, -4.228733, 
    -3.659206, -3.25061, -3.983162, -5.399307, -7.861031, -10.0006, 
    -10.93445, -10.09566, -8.951126, -6.408676, -8.062843, -8.504517, 
    -9.046703, -8.492016, -7.601913, -5.755558, -5.838112, -4.248268, 
    -3.6605, -4.046181, -4.105827, -3.887856, -4.040722, -4.383423, 
    -5.528736, -6.008163, -4.511555, -2.494621, -1.312065, -1.586548, 
    1.694443, 1.064751, 1.605377, 1.050957, 0.2780304,
  -6.557915, -5.975365, -2.359474, -2.05349, -1.016762, 0.1217804, 0.4577179, 
    0.3741226, 1.155632, 0.8035507, 0.2566757, -0.9339447, -2.940712, 
    -5.47847, -8.08577, -7.534988, -5.099571, -4.163368, -4.130043, 
    -4.717018, -5.216492, -5.595139, -5.073265, -4.797745, -3.05426, 
    -0.91259, -1.077179, -2.242538, -2.115189, -2.500084, -2.950874, 
    -3.644623, -3.847221, -3.813629, -2.794357, -1.982124, -2.797485, 
    -4.211815, -5.598785, -5.726913, -6.400085, -4.789932, -3.591751, 
    -0.9443741, -0.707901, 1.114487, 1.863457, 1.401215, -1.886547, 
    -4.286808, -4.210506, -3.187069, -1.945404, -1.663631, -0.9391518, 
    -0.8204002, 0.03142548, 0.2488594, -0.5964432, -0.6378517, -0.4188385, 
    -2.718578, -4.802692, -5.235756, -5.89748, -6.820652, -5.965206, 
    -4.953743, -5.026653, -4.970921, -6.164932, -8.794621, -8.766491, 
    -7.628731, -5.659462, -3.835236, -3.432899, -3.418587, -2.913372, 
    -3.943577, -5.685242, -6.220917, -7.258171, -8.886551, -10.75322, 
    -12.3165, -14.79567, -14.00504, -11.96807, -10.60635, -8.908951, 
    -7.718842, -8.136292, -7.815727, -7.200363, -6.738129,
  -13.71599, -14.65089, -13.21624, -10.98994, -10.4053, -9.858177, -9.087608, 
    -7.427704, -6.977188, -6.410774, -5.51963, -6.347244, -7.353752, 
    -10.9975, -12.24463, -13.2553, -11.87562, -11.78577, -11.66911, 
    -10.38786, -11.34984, -12.97927, -10.17248, -9.758415, -7.784462, 
    -7.022224, -5.611809, -3.584206, -3.511803, -2.785507, -3.332649, 
    -3.982391, -3.552956, -4.57795, -5.875092, -7.64801, -14.76807, 
    -10.75192, -10.48396, -8.589691, -9.568069, -8.393074, -6.092018, 
    -3.834717, -1.967789, 0.5290909, 1.849915, 1.145485, -0.9274292, 
    -1.398781, -0.8128433, -0.7993011, -1.35685, -2.119354, -3.634987, 
    -1.85894, -0.2758636, 0.5827179, 0.2626686, 0.5220413, 0.7431335, 
    1.34626, -2.676643, -5.341492, -6.288109, -5.057121, -4.443062, 
    -5.125099, -8.20974, -8.50061, -5.261543, -4.111549, -4.878731, 
    -5.339417, -2.742271, -0.8386307, -1.518326, -3.138885, -1.625343, 
    -2.908684, -9.183434, -9.011551, -9.324318, -8.753998, -9.005562, 
    -10.13838, -12.04437, -12.0303, -8.834213, -7.427437, -9.358688, 
    -13.50192, -14.62197, -13.1764, -11.52927, -11.35661,
  -7.449326, -7.606598, -5.123528, -2.886292, -3.529785, -3.941772, 
    -4.934479, -2.854004, -3.268333, -4.74334, -3.509727, -0.299057, 
    0.8678741, -2.577194, -4.303749, -6.863899, -6.672493, -7.976669, 
    -7.782135, -5.010521, -4.44516, -2.368324, -1.707901, -3.243065, 
    -4.12587, -3.94957, -4.645668, -4.381866, -2.988121, -2.779266, 
    -4.185776, -2.885262, -1.068336, -3.686562, -4.188911, -5.405319, 
    -4.46962, -4.014946, -5.00531, -4.060265, -5.86261, -6.350113, -5.086571, 
    -3.165474, -0.669632, -1.291252, -3.371719, -1.680824, 1.122818, 
    1.474648, -0.6693726, -1.899841, -2.067024, -2.893341, -3.82016, 
    -4.110001, -3.650879, -2.802185, -2.935265, -1.703484, 0.4598007, 
    1.04287, 0.7230759, -0.3685913, -0.578743, -0.2133789, 0.1392212, 
    -3.643074, -5.275627, -4.135773, -1.161812, 0.2735901, -3.251671, 
    -5.726669, -6.671707, -5.134995, -3.32093, -3.202705, -2.602959, 
    -3.046455, -2.212082, -3.385262, -4.51886, -7.024849, -8.011826, 
    -10.62927, -12.09515, -11.99567, -9.658699, -7.961304, -6.16156, 
    -4.337868, -2.650352, -2.095932, -1.375618, -4.044113,
  0.7756882, 2.158501, 0.1691818, -0.4644089, 0.818924, 1.784019, 3.441055, 
    2.884285, -1.618057, -5.792801, -6.074562, -0.4154587, -0.07274628, 
    -0.6990509, -2.607124, -1.187073, -0.8904572, -2.07431, -2.581856, 
    1.345482, 3.323868, 1.717613, -0.3750916, -1.613373, -5.44957, -6.323265, 
    -4.398262, -2.642281, -1.439934, -3.003212, -4.598007, -2.924568, 
    -1.430817, -3.191231, -6.156082, -4.370926, -2.230034, -3.155815, 
    -6.428215, -3.108421, 1.615791, -1.880035, -5.315453, -4.417015, 
    -1.065453, -0.2461853, -1.943573, -3.646698, -0.7480011, -2.093323, 
    -3.784988, -3.150871, -2.942795, -0.4555664, 0.8363724, 0.1264725, 
    -1.264153, -4.702171, -2.221184, 0.2863693, -0.7756042, -3.380295, 
    -1.063629, 0.2806396, -0.6847305, -0.9513855, 1.762146, 2.589233, 
    0.4923477, -3.583946, -7.034981, -7.036026, -3.954521, -1.435242, 
    1.418404, 2.161369, -2.041756, -3.133942, -3.127693, -0.4000931, 
    0.5897522, 0.2741318, 0.7499084, -0.2537384, -0.7105103, -1.52092, 
    -2.406082, -2.857903, -5.076393, -4.879776, -3.695145, -3.480293, 
    -0.3961792, 1.649651, 0.2629318, -0.08602905,
  -1.893311, 0.2637405, -3.077133, -1.403725, 1.021538, 0.488205, 2.143921, 
    4.285583, 4.551491, 0.9713058, 2.142387, 2.45697, -1.050331, -1.152687, 
    0.1100845, 1.179634, 3.604355, 1.139511, -0.3935623, -0.1909561, 
    -0.07794952, 1.39653, 2.724678, 1.379631, -0.6461487, -2.729485, 
    -2.831047, 1.357994, 1.891319, 0.9267273, 0.3251724, -0.680542, 
    0.02440643, 2.27076, 0.4408112, 1.175713, -0.2456284, 0.4410858, 
    0.09759521, 0.3947144, -0.02845764, 0.5489044, -0.9518814, -1.391479, 
    -2.1157, -3.524811, -2.799004, -0.9709091, 0.4569702, -3.58625, 
    -0.357605, 1.45356, -0.1141205, -0.5719376, 0.7895126, 2.287704, 
    1.255409, 0.755928, 4.368675, 3.759041, 2.742653, 0.5788193, -0.4459076, 
    0.4119263, 2.353836, -0.4073639, -2.912285, -2.738586, -1.361794, 
    3.023621, 5.297081, 2.336128, 2.875694, 2.693657, 5.825714, 4.201736, 
    2.043922, 2.358765, 2.695221, 2.579102, 1.305153, 0.8434296, 0.6986237, 
    0.1368942, -2.842247, -3.970657, -4.156342, -5.532898, -2.737045, 
    -2.392265, -1.794884, -4.531593, -4.448257, -1.264931, 0.559021, -2.080551,
  -5.783928, -2.006577, 1.268692, -0.03548431, -1.740173, -3.405525, 
    0.208786, 3.522331, 1.095268, 2.063499, 2.683258, 2.358261, 1.077805, 
    3.191864, 0.2960358, -1.030792, 2.702011, 0.5452423, -1.032623, 
    -1.153732, -0.6909637, -1.37561, -1.196442, -2.460495, -1.365448, 
    -0.947464, 2.919724, 0.8527832, -1.294357, -0.7169952, 1.863205, 
    -0.4607544, 1.812698, 6.078583, 3.582214, 4.10878, 4.69812, 3.786911, 
    3.598633, 3.034576, -2.47377, -1.312302, 3.133514, 3.174393, -0.04173279, 
    0.08222961, 0.3077393, -0.4987793, 0.8067017, -0.1789856, 2.962677, 
    1.294968, 1.067627, 2.729599, 3.864777, 3.865036, 1.096283, 2.128845, 
    7.846291, 6.232224, 3.848099, 2.017914, 4.665298, 2.389267, 6.984039, 
    5.956955, 4.831192, 2.509323, 7.746552, 8.149139, 6.568939, 5.472076, 
    5.436119, 0.5973206, 3.125717, 4.134834, 2.87204, 0.5548477, 4.250183, 
    4.696808, 5.012177, 2.632477, 0.552536, 0.06163025, 3.51712, 2.467117, 
    -0.8487549, 0.4025269, 2.956177, 4.529091, 2.794983, 1.408264, 3.037453, 
    3.767914, 3.972061, -2.198257,
  -2.505798, 0.09655762, 2.588745, 0.3788452, -3.035995, -3.34668, 4.55957, 
    5.694214, 3.200714, 6.030151, 6.880936, 2.41713, -0.4281769, 2.576233, 
    1.722336, 0.578064, 0.158783, -2.655014, -1.476624, 2.407227, 
    -0.07923889, 1.447845, -0.3716736, -2.087036, 2.145508, 4.508789, 
    5.490295, 5.627808, 2.80957, 4.353058, 5.904358, 2.67337, 3.953583, 
    4.733536, 2.723892, 7.690033, 12.63536, 5.425461, 5.638214, 7.522858, 
    2.671539, -0.1565704, 3.37207, -0.08444214, 6.301498, 11.92988, 8.504883, 
    6.605423, 5.779373, 2.781448, 3.680145, 2.282227, 1.835342, 4.22728, 
    4.272079, 3.60878, 0.7452393, 1.728058, 6.461395, 9.027542, 2.91478, 
    2.656708, 5.601761, 9.973877, 9.931702, 5.567123, 6.509033, 7.563995, 
    5.533524, 7.779343, 2.206955, 2.840302, 2.583267, -1.999283, 3.327545, 
    1.407211, -0.8047791, 10.40774, 9.502792, 7.431198, 3.574432, 2.318954, 
    1.87886, 3.892639, 8.365829, 7.505661, 5.09552, 7.687698, 6.550705, 
    4.494217, 3.473114, 1.755142, -0.2662048, -1.158142, 1.272598, 0.8462982,
  7.027039, 6.282242, 9.709061, 11.91766, 7.95932, 6.899689, 4.301254, 
    2.32782, 3.654892, 6.945007, 5.143967, 3.271561, 1.822083, 6.156982, 
    4.560623, 3.885635, 5.196045, 5.046051, 3.806198, 2.678589, 6.101257, 
    7.280426, 7.054901, 6.362976, 9.274429, 9.152039, 7.253342, 8.973648, 
    8.698898, 7.232498, 6.559326, 4.768967, 3.134323, 1.446045, 4.971558, 
    4.576782, 1.841629, -2.737045, 0.5463104, -0.5492859, -6.017517, 
    -0.5859985, 0.7124481, 2.777817, 5.822083, 11.17444, 15.66608, 10.75047, 
    4.029358, 2.455688, 10.81453, 7.593445, 3.012192, 3.253342, 1.239532, 
    5.579895, 6.871826, 8.60437, 7.995514, 4.267654, -2.141998, 1.321564, 
    7.534592, 8.172867, 5.253067, 3.768188, 5.336151, 6.906204, 3.320511, 
    1.990829, 4.022095, 2.59552, 0.5090637, 3.657242, 6.915573, 7.817398, 
    21.52313, 31.27884, 17.13354, 1.30722, -2.082886, 0.5705109, 2.666351, 
    1.676773, -2.754486, -0.2297363, 0.5043793, 1.548645, 5.174942, 5.106461, 
    4.187439, -0.04536438, -2.557617, 4.621826, 4.930161, 7.282761,
  1.584061, -2.07193, -0.3198547, -1.100586, -1.88913, -0.8701172, 0.7611389, 
    0.04679871, -0.01881409, -5.454742, -2.813095, 1.327805, 4.890823, 
    3.42363, 0.6366577, 4.53067, 5.453064, 3.516083, -0.9310608, -0.8766327, 
    -0.2055359, 2.417648, 3.583267, -0.3011017, 1.89447, 5.718933, 3.990036, 
    3.71582, 2.842392, 1.060089, 2.861908, 0.880661, -2.443298, -3.843033, 
    -4.210739, -4.83548, -8.457367, -2.481842, 5.357224, 3.656189, -5.593811, 
    -6.099289, -5.180283, -4.556061, 0.2551422, -0.8018951, 2.789261, 
    10.13979, 1.485352, 4.642899, 4.857498, -0.3498077, -3.218292, -5.878448, 
    -3.006577, -2.465958, -0.434433, 0.6293793, -1.709183, -6.370895, 
    -4.106583, 2.062698, 5.470016, 3.613739, 1.918945, 4.545517, 2.012177, 
    3.625458, 6.760376, 7.765564, 11.50227, 10.21817, 8.229889, 7.381439, 
    2.93718, -0.6813202, 16.17155, 20.59161, 9.150986, -1.987823, -8.378189, 
    -10.21152, -5.974274, -5.720383, -6.271164, -6.404739, -2.468292, 
    1.23613, 3.452011, 4.515564, 0.5462799, -0.01257324, 1.186386, 2.617645, 
    2.385086, 4.51503,
  -0.3180237, -1.211517, -3.530533, -2.107361, -2.800568, -5.141464, 
    -6.017487, -0.7154236, 1.026001, -1.696426, 3.334839, 3.370773, 1.68457, 
    1.164001, -5.991211, -10.66647, -15.05397, -14.03236, -5.125061, 
    -4.21907, -1.054489, -0.5318298, 0.9436951, 0.1509705, -0.08027649, 
    2.336655, -6.646423, -6.778442, -4.52298, -2.227402, -4.728714, 
    -10.42947, -12.65889, -13.82635, -12.12323, -6.525833, -5.338852, 
    -5.269592, -0.3484802, -10.22766, -24.84744, -16.5761, -14.6433, 
    -8.331573, -5.055527, -7.318817, -1.423767, 3.225464, -1.794861, 
    -3.764908, -5.422729, -8.732361, -1.444855, -2.319077, -4.14563, 
    -5.489136, -6.091995, -5.097473, -3.87793, -3.38913, 1.32962, 3.457489, 
    -1.060226, -2.492264, -1.55658, -4.540161, -0.5159607, 0.3988953, 
    0.8403015, 3.315811, 3.993423, -3.378983, -4.606323, -1.914383, 
    -3.541977, 4.090317, 4.821289, 3.920288, 0.372345, -15.14043, -11.67923, 
    -7.505264, -7.145905, -3.78183, -1.213089, -0.2985077, 1.26503, 
    -1.477936, 1.840042, 1.329895, 3.089767, 5.347855, 4.249405, 1.406708, 
    -2.463348, -2.329498,
  -6.441193, -4.539368, -5.987289, -2.220093, -2.235748, -2.997955, 
    -2.304749, -1.610733, 3.462173, 1.238754, 1.991623, -1.069061, 
    -0.8898926, -2.284424, -6.058136, -5.153961, -7.559967, -2.207092, 
    -3.169083, -5.557877, -3.360748, -0.8195953, -0.03234863, -1.248245, 
    -7.045639, -9.996674, -8.907867, -6.681839, -3.659958, -4.854736, 
    -9.793518, -12.60916, -14.78285, -17.05188, -11.61047, -11.19847, 
    -12.61723, -13.92062, -12.43286, -19.51256, -22.73885, -7.776611, 
    -7.638336, -8.455521, -4.662033, -3.47142, -3.931046, -1.289917, 
    -7.348511, -4.108658, -7.422455, -3.976624, -0.5341797, -7.93158, 
    -7.566208, -4.117508, -2.756317, -1.378967, -1.912048, -2.92247, 
    -1.532883, 1.112167, -2.551102, -0.2617798, -1.651108, -1.79747, 
    4.312958, 4.334045, 0.02026367, -0.5266113, -5.25058, -9.27739, 
    -7.341705, -1.834946, -1.950836, -2.118256, -1.554474, -2.286011, 
    3.096802, -4.739655, -4.725845, -0.8240204, 2.00592, -3.846405, 
    -4.411255, 3.453323, 5.252014, 3.867386, 3.516861, 3.37233, 4.991074, 
    3.983795, 3.212189, -1.943268, -0.223999, -4.222183,
  -7.338074, -5.948746, -6.285217, -9.691193, -2.664917, -1.394562, 
    -0.7068176, 1.578049, 1.480423, -5.250046, -1.151093, -2.395874, 
    0.5207825, 2.916885, -4.891739, -2.42012, 1.955933, -1.90657, -0.4391327, 
    0.6783447, -1.650818, -0.7870331, 1.295258, -6.764114, -8.928955, 
    -5.707367, -3.789124, -2.350311, -0.3453522, -4.553192, -8.342743, 
    -12.69275, -19.67896, -21.65526, -15.16492, -10.89145, -8.750305, 
    -12.12143, -13.29692, -11.17712, -7.450562, -1.28389, 2.069489, 1.812714, 
    -2.290939, -3.981567, -6.260223, -8.493546, -10.20786, -10.01411, 
    -9.340164, -4.735474, -4.669601, -4.265671, -7.892761, 3.118164, 
    1.329102, -0.7424927, -2.60759, -2.265945, 1.811142, 4.433273, 2.679901, 
    4.536407, 1.724426, 0.1502228, 2.660889, 0.4309387, -3.668808, -1.924789, 
    -10.45032, -3.998489, -2.522705, -2.465149, -6.122971, -4.79953, 
    -0.5222168, -3.551361, 8.334045, 5.943695, -6.886002, 8.271545, 4.285095, 
    2.902786, -2.613327, 1.112717, 3.406708, 0.903595, 5.642914, 6.357498, 
    6.128067, 4.321823, 3.720001, -5.763855, -1.744843, -8.17244,
  -5.789108, -5.100067, -3.219574, -0.2498169, 1.087982, 4.953323, 1.920258, 
    1.298889, -2.191452, -1.984161, -5.12973, -12.16074, -13.45891, 
    -0.3266144, -1.103439, -0.2935333, 9.184601, 0.7059326, 0.2892761, 
    -1.190414, -1.758652, -0.5260925, -2.623749, -5.093796, -4.320358, 
    1.778336, -2.781815, -0.6773834, 2.778625, -2.681549, -9.554474, 
    -16.87038, -20.39748, -16.57819, -15.48965, -15.33289, -15.77844, 
    -14.5347, -13.7477, -12.59978, -3.071411, 2.840317, 6.471573, 1.216354, 
    -0.9849396, -6.238846, -6.727921, -12.37636, -19.45891, -18.68677, 
    -11.9102, -2.783386, -0.2870331, 2.518448, -0.7331238, 3.270264, 
    0.5476074, -4.542496, 2.033295, 6.272079, 3.690308, 3.821045, 1.959595, 
    -0.9797363, 4.239273, 1.966354, -4.924271, -3.787552, -6.579468, 
    -5.755249, -6.670883, -4.122971, -8.043533, -2.476608, -3.08783, 
    -2.233398, -2.61908, -3.868835, 8.991364, -1.582092, -7.570892, 15.45905, 
    9.952301, 8.403595, 2.349152, -2.84198, -1.469315, 2.257507, 2.796829, 
    1.27182, 3.907761, -2.048492, -3.992767, -6.209686, -5.732849, -10.83598,
  -5.323486, -3.324799, -6.950043, -4.222717, -4.699799, 3.616898, 4.802826, 
    2.338745, 3.264526, 6.872864, -7.796127, -12.58755, -18.54251, 
    -0.1292114, -1.55603, -6.115677, 1.731979, 6.946823, 0.4483795, 1.990311, 
    1.349442, 6.358292, 1.719742, 5.801514, 7.838226, 4.334854, 0.1371918, 
    -0.06932068, -2.114624, -4.87558, -15.16125, -17.47559, -20.48993, 
    -16.62323, -17.08679, -19.64825, -13.5563, -7.202942, -7.217224, 
    -6.787018, -6.712814, -6.89328, -2.032089, 1.859589, 3.618439, -4.789886, 
    -11.35422, -15.74692, -15.22505, -13.92297, -5.125305, 3.299957, 
    4.427567, 3.913498, 4.072083, 1.627548, 3.584076, 0.2121887, 1.334839, 
    3.333282, 1.721832, 2.786926, -3.517242, -5.463348, -5.263855, -8.702911, 
    -8.930786, -9.035461, -11.69041, -3.765152, -4.363068, -5.460983, 
    -6.014114, -3.473999, 0.8710632, -10.49825, -2.218292, -2.086273, 
    18.48431, -2.806061, -2.189636, 14.35828, 7.913757, 10.07858, 9.054886, 
    12.73613, 2.545013, 3.303345, 3.745514, -0.5560303, -0.658371, -8.019318, 
    -4.952652, -7.26828, -3.304214, -4.653168,
  -2.551605, -3.530273, -2.132874, -2.055267, 3.261658, 6.462952, 7.232483, 
    1.237213, 6.447083, 10.27858, 0.3702545, -4.499527, -4.088593, -2.686005, 
    0.4483948, -8.04068, -2.643799, 4.738495, 6.793945, 2.197876, 2.588242, 
    -1.683899, -0.4031677, 3.190842, 0.9744263, -2.78598, -2.944061, 
    -4.990662, -8.499542, -12.48392, -14.31046, -11.30865, -12.76935, 
    -10.86279, -19.3761, -18.58575, -8.611755, -10.6037, -5.008652, 
    -3.804733, -0.3182831, -5.210464, -0.7888489, 5.136154, 6.320511, 
    -0.05838013, -9.645615, -4.072189, -12.09041, -10.67192, -5.679993, 
    4.967651, 4.523392, 2.017136, 4.343704, 1.368973, 2.965836, -1.45787, 
    -2.630508, -1.446136, -4.378967, -9.415161, -7.796661, -7.242508, 
    -9.020889, -2.794586, -7.113068, -3.566193, 0.1022949, 0.7124634, 
    -3.807602, -2.542496, -3.335983, -4.998489, 3.348648, -1.869598, 
    -1.605804, 6.23822, 16.33455, 3.572601, 1.938751, 4.669205, 0.4012604, 
    5.87207, 10.0377, 12.59657, -2.760468, 0.06402588, 0.08432007, -3.907867, 
    -5.056046, -7.830505, -4.918274, -2.657074, -3.594055, -3.176346,
  2.813751, 2.402313, 3.118713, 5.541885, 19.36218, 10.40645, 3.517639, 
    -3.359161, 1.525223, 3.450485, 3.176758, -2.243271, -5.758118, 4.220779, 
    8.347351, -2.857605, -3.337799, -0.6531677, 0.5762482, -1.264374, 
    -4.304474, -6.432877, -2.38623, -1.944305, -3.236237, -2.195862, 
    -1.969574, -0.9912109, 1.605438, -5.830811, -7.18808, -8.581573, 
    -6.782867, -4.299805, -9.03363, -22.22427, -9.934174, -12.92999, 
    -11.67921, -14.06332, -9.604477, -0.5646362, 0.1796265, 1.264526, 
    0.1374512, -5.04953, -6.228943, -4.080002, -4.333633, -11.21098, 
    -0.8490143, 2.133026, -8.445892, -3.727386, 0.297348, -1.163589, 
    1.296051, -2.042236, -4.209412, -3.315674, -1.462555, -6.426605, 
    -5.457855, -2.712296, -5.066452, 0.6202698, 0.9533386, 4.392395, 
    4.275986, 11.0786, 7.777557, 8.185379, 6.922058, 4.511414, -2.574005, 
    -7.1409, -6.001892, 9.816574, 11.6067, 4.341339, 0.08978271, 1.623871, 
    -0.4768982, 10.03484, 13.51192, 8.421799, -7.178955, -5.33287, -3.855499, 
    -5.152924, -6.097473, -5.561768, -2.344055, -2.036255, -2.55838, -1.302643,
  1.181732, -1.280548, 1.40332, 3.600739, 13.85619, 12.81374, 8.281967, 
    -8.778717, -14.70189, -19.3644, -17.68861, -17.65291, -11.52191, 
    -2.007339, -0.8227081, -5.302673, -0.9164429, -0.5799866, -2.370361, 
    -7.47374, -6.546158, -6.673248, -1.130249, 1.562958, 1.848145, 7.112732, 
    6.670532, 9.578064, 1.876221, -2.374023, -1.771149, -3.406036, -4.576904, 
    0.8424072, -1.055786, -12.41696, -16.13028, -13.6886, -17.98366, 
    -23.72713, -15.02272, -10.51752, -9.849808, -4.971939, -12.02585, 
    -16.72246, -16.70215, -6.59668, -7.743286, -11.47427, -8.665955, 
    -7.085739, -9.390411, -12.92635, -5.787277, -2.503693, -1.394318, 
    -0.4393616, -1.788071, -1.501617, -1.903687, -3.509155, -1.749542, 
    0.6494446, -1.989624, 2.28952, 5.189804, 6.18927, 6.951782, 11.52312, 
    12.01817, 8.768188, 8.541077, 3.204926, -10.72556, -13.32378, -1.326393, 
    4.720779, -4.539124, 1.00853, 1.47908, -4.379242, 1.236923, 5.806442, 
    17.84709, 20.31949, 10.29889, -0.7776489, -1.094086, -5.420898, 
    -1.267242, -2.838348, -0.5873108, 0.3564758, -0.6873169, -1.269348,
  -2.245911, -0.2292175, 2.007507, 7.692108, 22.54889, 17.3968, 14.77104, 
    3.413239, -19.97897, -36.7886, -27.83183, -20.68784, -13.80008, 
    -7.758667, -0.500061, -1.905518, 0.6655579, 7.716339, 4.042419, 1.579376, 
    0.9306641, 0.1179199, 1.337708, 5.001526, 2.616638, 7.588745, 9.968201, 
    5.28537, -2.601624, -5.117752, -1.73938, -4.956573, -3.135986, 6.244476, 
    -0.9985046, -3.04303, -9.195862, 1.661392, 6.67881, 6.831421, -5.914139, 
    -15.05655, -10.81178, -2.628464, -5.514389, -8.594589, -1.94278, 
    -3.563858, 0.8741455, -1.678192, 2.378311, 3.698624, 1.794724, -2.656326, 
    -6.954468, -5.110458, -5.570358, -6.858643, -8.442505, -6.807343, 
    -2.643021, 1.591354, 1.110107, -1.452393, -2.237549, -1.718018, 
    -4.786743, -3.896912, -1.43988, -5.579742, -3.870605, -8.497955, 
    -9.12793, -5.760468, -12.46802, -16.1472, -11.00061, -7.186493, 
    -2.514374, -7.92247, 6.529633, 6.747589, -0.735199, 5.661911, 12.01503, 
    7.347092, 15.78069, 2.257782, 0.4840393, -0.544342, 0.1090698, 
    -0.6925049, 0.3585205, -0.2185364, 0.1806641, -0.6156921,
  -0.4360046, -2.004517, 1.048645, 9.319763, 16.19945, 14.62051, 21.1924, 
    23.87231, -11.95918, -50.00108, -21.20552, -6.044342, -3.734161, 
    0.6642456, 1.268951, 3.016083, 0.5616455, 1.530914, 3.839264, 7.915833, 
    3.808258, -2.832123, -0.6003113, 4.037994, 5.36792, -0.8914795, 
    -4.894348, -8.569855, -0.2399139, -0.2065735, -3.238846, -4.052391, 
    13.17806, -0.2490387, -0.8466644, 1.018433, -3.93338, -11.24954, 
    -7.637299, -13.51857, -19.50972, -14.55138, -5.416977, 3.104645, 1.22287, 
    9.025726, 10.42233, 14.42809, 18.66246, 20.34135, 17.1028, 14.79579, 
    14.52287, 11.11166, 8.474945, 6.503326, 1.452026, -4.559692, -5.44693, 
    -9.032593, -7.462311, -9.237579, -5.31308, -8.345123, -2.204224, 
    -2.106567, -3.862305, 0.1530457, -0.2929993, -8.588867, -1.431305, 
    -10.42192, -18.41983, -18.58078, -10.5295, -6.054489, -12.52974, 
    -3.738358, -15.46281, -15.89171, -10.21646, -4.18988, 0.5515137, 
    15.23015, 10.54735, 1.836914, 1.188477, -3.086792, 2.38562, -3.753448, 
    1.32074, -0.2219543, 1.136414, -0.5297546, 0.3436584, -1.50058,
  1.52652, -1.257355, 2.184296, 20.06844, 23.41687, 13.7554, 14.44579, 
    20.07832, 4.168961, -26.05034, -24.35422, -5.195923, -2.870117, 2.717651, 
    -2.913849, -1.362061, -0.7748108, 1.613464, 1.492401, -1.92688, 1.032745, 
    2.00827, 0.8004456, 0.8720703, 5.968933, -4.99588, -1.046936, 18.53014, 
    1.035339, -0.01596069, -13.07272, 8.220741, 4.665833, -7.272705, 
    -7.114105, -4.851074, -9.265686, -14.99225, -14.11594, -11.11516, 
    -11.5675, -11.0524, -8.282074, -4.968018, -2.414093, 0.9934387, 
    0.3715515, 5.326263, 9.839264, 10.8252, 13.0351, 10.51245, 11.40933, 
    9.279907, 11.16165, 12.01816, 6.483795, 3.188751, 0.6160889, -3.339142, 
    -3.540161, -6.19223, -7.437042, -1.922211, -4.217255, -3.98288, -3.96698, 
    -3.227692, -5.932861, -10.22482, -11.49796, -19.02037, -26.26646, 
    -28.75189, -16.51752, 1.780117, -22.41466, -11.44276, -14.58807, 
    -17.28549, -7.881592, 1.174438, 11.00333, -0.8188171, 1.500458, 1.121796, 
    6.821808, 3.938202, 5.324921, 4.289276, 0.8988953, -1.00528, -3.230011, 
    -1.513855, -1.472717, -1.464142,
  0.4981384, 0.2330017, 5.73407, 12.51193, 12.43744, 17.70726, 11.23849, 
    6.678864, 6.643188, -10.65863, -18.41333, -6.584961, 0.3202515, 8.247833, 
    3.359558, 1.821808, 2.953857, 2.286407, -2.870636, -3.038879, -2.039398, 
    -2.076111, 0.1934204, 2.078339, 3.103851, -1.505768, 13.01295, 17.31531, 
    -5.634949, -0.3630676, -7.398773, -0.2146301, -6.298218, -1.240936, 
    -3.346405, -4.264618, -2.803436, -3.451324, -0.7388611, -1.103729, 
    -2.784698, -2.869049, -2.668304, -5.009979, -4.646149, -4.483154, 
    -2.603943, -1.995636, -4.236755, -5.962799, -0.1104431, 0.3470764, 
    0.3996887, 7.412445, 9.544739, 12.401, 13.96663, 15.33327, 12.2739, 
    11.09578, 8.739532, 6.983826, 8.38147, 8.589783, 3.420258, 1.918427, 
    -0.3875427, -0.6938171, -3.866486, -7.18158, -13.45581, -9.408936, 
    -13.45865, -21.32504, -23.36229, -6.675598, -22.94328, -13.01022, 
    -12.91776, -1.810211, 5.621826, 3.03511, -1.953415, -5.388077, 
    0.04421997, -0.5688171, 1.477814, 2.237427, 1.841339, 3.709564, 3.379883, 
    -2.288605, -10.79095, -5.466217, 0.2939606, 0.2171326,
  -2.85318, -6.039917, -2.25708, 1.31842, 1.397583, 2.417114, 0.7363892, 
    -1.445404, 5.730133, 10.69629, 17.99084, 2.627289, -1.044098, 0.4543457, 
    10.86221, 9.668182, 8.227539, 7.915039, 4.287689, -2.276886, -10.27612, 
    -6.753723, -5.834717, 1.496552, 0.8609009, -4.579254, -2.14328, 
    -0.9508362, -4.402679, -3.882874, -8.457336, -9.32663, -7.337036, 
    -2.760468, -4.29744, -4.132874, -0.07321167, -2.033112, -0.724823, 
    -0.1971741, -0.5750427, -4.783661, -2.305023, -4.448761, -2.666992, 
    -1.717255, -1.599304, -1.653473, -0.6860046, 1.842377, 3.079895, 
    2.609314, -1.24173, 6.620514, 7.559326, 12.37701, 13.06949, 17.40984, 
    16.01401, 14.86946, 15.2536, 10.36298, 7.348114, 9.680939, 8.340057, 
    6.911133, 6.119476, 1.880646, -2.15448, -4.330292, -4.516479, -6.449524, 
    -9.150848, -9.455261, -5.269852, -4.296143, -8.990448, -7.81543, 
    -1.78418, 5.685364, -2.226608, -2.222717, -0.2279053, 3.790833, 
    -1.858643, -2.061249, -0.2445831, 1.184082, 1.50647, 2.511139, 2.778625, 
    -5.070129, -4.534698, 0.0657959, -3.415436, -3.193298,
  0.6791077, -1.970886, -0.250824, 0.879364, 2.375732, 0.2145081, 1.087952, 
    0.7278137, 0.342926, 4.643677, 8.634827, 0.3408203, -1.611542, 
    -0.2932739, 10.12753, 3.750214, 7.67337, 5.109558, 0.7280579, -8.015167, 
    -10.67792, -10.09875, -2.572205, 0.2252197, -1.225037, -3.109436, 
    -11.79822, 2.479858, 6.141876, 2.839783, -5.292236, -8.155792, -7.259949, 
    -4.14563, -3.77478, -3.414124, -1.78183, -0.9823608, 1.27832, 2.078033, 
    -0.5253296, -1.438873, -2.90448, -3.214111, -2.845123, 3.32312, 3.840851, 
    3.933533, 0.986145, 1.503326, 4.496826, 3.356201, 3.315826, 5.13797, 
    4.988754, 9.877563, 3.95282, 8.229385, 12.11476, 11.05696, 13.90096, 
    14.92157, 14.81949, 14.87912, 14.40021, 10.63403, 8.24707, 3.373352, 
    -1.545624, -6.43808, -8.742493, -8.609955, -8.705017, 5.366608, 4.43277, 
    -6.335983, -8.47583, -11.4097, -1.08078, 7.388229, 0.2746887, 3.137192, 
    0.8692169, 3.64917, 2.063232, 0.6504669, -0.05654907, 3.863739, 3.177795, 
    2.337677, 1.373413, -1.787781, -0.2492676, -0.2601929, -0.1365356, 
    -1.151642,
  1.420258, 1.985077, 3.773346, 5.704102, 4.647369, 2.046814, 3.30777, 
    1.899933, 0.9499207, -0.9735107, 2.877014, 1.278839, 4.473877, 3.03717, 
    0.6803894, 4.832764, 5.991364, -1.638885, -3.799561, -10.22012, 
    -13.76855, -10.53888, -11.28625, -9.083679, -1.793274, -6.208649, 
    -8.516998, -6.610199, -1.667755, -10.59879, -11.27609, -1.007874, 
    -0.1716919, -1.862305, 1.389771, 2.242645, 4.489532, 2.033264, 2.036682, 
    -3.518555, -4.894318, -4.816711, -1.859436, 0.1444702, 0.807251, 2.36087, 
    0.3377075, -0.6867676, -0.03234863, 0.5848541, 0.9259949, 0.7548981, 
    -2.671921, -3.51619, -0.6443176, 3.044998, 0.9723511, 1.270264, 8.223373, 
    0.3889771, 5.227798, 14.57338, 17.14915, 14.04709, 14.49292, 13.5838, 
    8.371307, 4.028839, 5.304352, 5.460632, 4.077301, 11.27209, 17.59889, 
    1.197861, 0.9267731, 3.19162, 1.371048, 2.725204, 2.764511, 2.95697, 
    1.086411, -0.2932739, -3.863861, -3.00708, 0.7113953, 2.197876, 1.888748, 
    5.499176, 3.873901, 5.524414, 2.960083, 1.562469, 2.012451, 0.5218506, 
    -0.3081055, -0.942749,
  1.943695, 1.303558, 1.809814, 2.162689, 3.275726, 3.655914, 2.592377, 
    3.264526, 1.196014, 0.7580261, 2.604614, 3.507202, 9.366089, 6.402802, 
    5.449951, 4.832245, 0.7973328, -6.793549, -1.870636, -3.944885, 
    -9.859985, -12.18939, -10.74667, -11.65033, -9.620636, -16.62585, 
    -20.91595, -19.50967, -18.01228, -20.29407, -4.166718, -2.811523, 
    -5.335724, 2.706207, 3.906982, 5.431976, 4.509308, -1.713318, 2.301239, 
    0.7538452, -0.9450989, -7.810974, -1.160736, 3.166107, 1.189026, 
    2.704117, -0.3646393, 0.3848572, -3.816452, -4.751877, -2.633377, 
    -5.15448, -2.764374, -0.7669678, -1.068802, 1.81662, 2.973648, 0.6416016, 
    2.948105, 2.292114, 3.145767, 3.575974, 8.020264, 11.46974, 7.842377, 
    6.900726, 4.426208, 6.855652, 8.244995, 14.86011, 15.0036, 23.37105, 
    23.90384, -1.411514, 2.888229, 5.189255, 1.41011, -0.6333771, -5.257599, 
    -4.560471, 0.8517761, -7.08754, -5.608124, -5.281311, -6.569839, 
    -3.147446, -0.05084229, 2.199173, -1.753448, 4.972595, 1.976257, 
    1.683807, 1.918427, 0.5072327, 1.652008, 3.712677,
  -1.291229, 0.8613892, 2.909821, 1.404083, 0.416626, 1.478058, 2.545013, 
    1.184052, -0.2872925, 0.4179077, 1.81897, 1.926758, 3.672058, 8.302795, 
    11.20929, 8.326233, 6.366333, 4.812164, 0.8965454, 0.4832764, -0.8240051, 
    -7.074554, -6.12558, -10.62949, -10.22897, -13.6011, -15.63989, 
    -18.60135, -27.33704, -18.72351, -10.60294, -7.96907, -5.38002, 
    -4.632874, 2.589005, 4.003326, 7.735901, 3.070267, -1.466461, -4.869568, 
    -6.363602, -1.770615, -2.075043, 0.1048889, -1.652924, 3.927551, 
    2.804642, 0.6986542, 0.2947388, -3.334946, 1.440842, -5.101608, 
    -1.342484, -0.8953705, -2.766983, -3.093277, 0.3957825, 0.6361389, 
    2.575714, 0.3444824, 0.2908173, -0.6963959, 0.405426, 2.353348, 4.221817, 
    1.437958, 0.4590454, 3.582245, 6.720261, 13.23924, 10.01817, 8.118164, 
    4.50177, 4.217651, 4.947342, 5.608795, 0.2437134, -4.381042, -6.908127, 
    -6.873749, -4.697449, -6.651611, -5.201096, -12.50214, -13.1089, 
    -7.976364, -3.907074, -2.48468, -4.088318, -3.414368, -7.122681, 
    -0.7375488, 0.01687622, 0.3535767, 0.6705017, -0.9721985,
  -1.437317, -0.9656677, 0.004089355, 2.766602, 4.917145, 4.668182, 4.392914, 
    3.518158, 3.271301, 3.328094, 0.4462891, -0.5672607, 0.3632202, 6.027039, 
    12.65228, 13.851, 12.23668, 13.24371, 11.47781, 6.294983, 3.873657, 
    0.2835388, -2.416718, -6.463348, -1.756042, -8.247437, -19.44301, 
    -18.76724, -34.32401, -17.78393, -1.670639, 6.219208, 9.075974, 4.367401, 
    2.193176, -0.6060486, 1.452545, -0.3365173, 1.855667, 5.267639, 
    0.4942017, -0.3813019, -2.465927, -4.982071, -7.374268, -5.042755, 
    3.369736, 5.516357, 1.367661, -0.1271362, 0.2226105, -2.844055, 
    0.09318542, 0.7236328, 0.1127014, -0.1920013, -4.632874, 1.004364, 
    0.3608704, 0.4194641, 0.4897766, 1.592896, 6.167664, 7.174957, 3.760635, 
    -0.5987549, -2.759949, -1.106842, 6.695267, 7.950729, 13.2226, 10.42833, 
    5.905411, 5.819977, 5.952026, 2.991333, 0.4619141, 0.5215454, 
    -0.02012634, -4.03392, -3.695114, 0.3757172, -2.888321, -6.906296, 
    -1.753967, -3.671677, -5.399536, -4.697464, -4.76593, -5.00058, -7.77713, 
    -5.091187, -0.59198, -1.831573, -0.4271545, -0.156311,
  1.616089, 1.765839, 1.291885, 4.120255, 7.405151, 6.116348, 14.05463, 
    10.83823, 8.53511, 14.51479, 10.71375, 5.666885, 3.115326, 7.838501, 
    12.01141, 13.78769, 13.30957, 22.24551, 32.358, 20.37833, 15.04996, 
    1.694733, -6.384949, -8.144318, -2.703186, -4.72348, -8.018799, 
    -13.35031, -29.94121, -17.17116, -3.364395, -1.10527, 4.265564, 7.005417, 
    9.423645, 6.738235, 6.98616, 1.136658, 0.9358826, 2.045258, 4.200714, 
    1.326248, 1.941071, 3.119736, -1.812576, -4.884171, -5.17897, 0.08796692, 
    -1.128448, -3.735214, 1.79837, 1.091339, 0.3525391, -1.746429, -1.959961, 
    -0.5789642, 1.058792, 1.59993, 2.835098, 1.054626, 3.379623, 2.304092, 
    1.518433, 4.162949, -0.8872833, -0.7008209, 1.832245, 4.698898, 11.34525, 
    2.950211, 3.827271, 4.443695, 3.354889, 4.130157, 6.530167, 0.3369141, 
    2.011139, 4.899933, 6.291107, 6.879883, 3.388229, -1.058136, 1.843689, 
    5.222061, 6.290298, -0.6795044, 3.534836, 5.833786, 3.987686, 3.674667, 
    5.61322, 4.029099, 0.3121796, -1.372437, -4.407089, -1.25943,
  7.459045, 15.22235, 21.26765, 12.92781, 5.624146, 4.402023, 1.717911, 
    1.556183, 8.505936, 16.39941, 21.15228, 23.42233, 20.02625, 15.18353, 
    7.04422, 8.809036, 13.13718, 10.60672, 6.915314, 3.582474, -1.538605, 
    -9.83728, -9.849014, -8.351868, -13.57271, -10.62531, -2.32843, 
    0.3043671, -14.23575, -15.77611, -4.909424, -4.006317, -0.7878265, 
    1.272842, 5.700455, 1.809052, -1.328995, -0.1011047, 3.130417, 1.314774, 
    -0.343811, 3.37442, 2.048111, 1.572067, 2.959305, -0.3284607, -1.51152, 
    0.4241638, -0.6094208, -3.28157, -4.707596, 0.3486481, 1.396576, 
    2.020798, 1.516876, 3.283264, 2.519974, 4.96817, 0.8663483, 3.660614, 
    1.129364, 1.60202, 2.483795, 0.5502014, -2.078186, -2.004227, -0.3203735, 
    2.807495, 3.089523, 1.160355, 2.878067, 2.196548, -3.200043, -3.881042, 
    -2.519577, -0.9581299, 0.3866577, -3.602386, -2.03157, 4.141342, 
    6.617126, 3.033279, 3.156204, 4.623917, 4.590057, 9.313751, 9.308807, 
    5.460617, 4.230423, 4.304367, 5.256439, 2.049164, 0.343689, -0.1448669, 
    -3.255524, -2.955795,
  4.971039, 4.008804, 2.804382, 3.152298, -2.031311, -2.163849, -6.751114, 
    -6.840164, -0.2094574, -1.118042, -1.652664, -8.714645, -5.072983, 
    -2.487045, 3.478317, 10.07703, 12.19162, -0.2146454, -4.257339, 
    -3.436005, 0.2423859, -7.908401, -12.89848, -11.81412, -7.441467, 
    -12.04564, -7.363861, -0.1826172, -4.006836, -7.297729, -4.667252, 
    -4.531845, -5.102661, -6.400314, -6.423248, -1.48262, -6.061264, 
    -14.91179, -6.081039, -3.314636, -8.141998, -3.96022, -0.5623016, 
    -1.546936, 0.8298798, -2.073517, -3.007614, -1.384445, -1.664124, 
    -2.971939, -8.593033, -5.297974, 2.356964, 1.383789, -0.7664642, 
    0.1689453, 4.087433, 6.181961, 3.092117, 2.973633, -1.168289, -0.141983, 
    -0.1950989, -7.727417, -13.96413, -16.96516, -20.14174, -15.2058, 
    -2.887833, -1.637039, -3.323242, -7.270615, -8.035995, -12.29929, 
    -13.92609, -12.85838, -7.664383, -5.879501, -5.791992, 1.708267, 
    2.049408, -0.09745789, 1.43457, 4.526749, 6.825195, 2.212967, 2.316605, 
    -0.1914673, -0.1651764, 0.8546448, 1.073639, -1.999268, -1.878967, 
    0.5858917, -0.5354767, -2.773239,
  -5.184708, -6.697723, -6.969315, -12.76363, -13.71959, -11.41623, 
    -17.29044, -17.29591, -19.04355, -10.95087, -10.56075, -19.9084, 
    -21.63287, -0.08964539, 3.882492, -9.256317, -12.3123, -10.61829, 
    -13.13756, -13.62401, -8.871429, -10.44589, -14.91518, -12.90422, 
    -8.064377, -8.863617, -8.349548, -5.870117, -7.255524, -6.556839, 
    -8.759445, -8.053192, -5.823242, -4.682358, -2.439117, -1.482086, 
    -3.500076, -5.648239, -14.31437, -8.501633, -6.62793, -3.656052, 
    -3.758392, -0.9565735, -5.406311, -5.805038, -1.774292, -2.32872, 
    -8.475327, -4.633148, -1.629517, -2.780289, -2.840439, -0.09797668, 
    -3.055283, -4.604492, -3.643311, 1.162155, -0.8151855, -2.365433, 
    0.9408112, 0.6767578, -2.36908, -12.75007, -28.72948, -28.00945, 
    -20.77663, -11.59435, -11.45657, -9.409164, -11.8438, -11.87506, 
    -9.716202, -12.86803, -7.984436, -15.0782, -12.64616, -11.25945, 
    -6.656845, -6.323242, -0.4245453, -0.1946106, -3.287048, -3.472992, 
    -2.737579, -2.228729, -0.3183136, -0.5756073, -6.297974, -5.966217, 
    -6.870636, -9.010483, -2.065689, -5.827667, -10.28731, -4.193825,
  -12.88707, -13.92428, -24.85215, -28.37299, -17.1451, -18.05447, -18.16776, 
    -18.86076, -21.17429, -21.07246, -18.97325, -21.9584, -14.55475, 
    -10.39357, -13.58313, -16.51959, -11.43497, -10.2795, -13.0472, 
    -13.11752, -11.79642, -13.49849, -9.646683, -11.17609, -13.03574, 
    -10.36125, -8.949295, -6.832336, -8.677139, -6.935471, -4.451355, 
    -3.978699, -4.149002, -5.060196, -5.745377, -3.756836, -0.8464203, 
    1.208801, -4.144333, -10.88704, -8.145386, -1.905273, -0.4032135, 
    -0.8612671, -2.516724, -4.620361, 1.896835, 3.316078, -4.719864, 
    -6.526894, -2.94799, -1.003967, -3.048767, -2.943039, 2.064247, 
    -1.249283, -4.743301, -4.745377, -1.525856, -0.5636139, 0.09289551, 
    -0.4873199, -1.452927, -8.21389, -22.98549, -15.44176, -18.4321, 
    -16.82741, -13.22794, -7.680283, -9.909698, -6.185211, -6.575836, 
    -26.67245, -9.312332, -3.221176, -4.370911, -4.447189, -4.920639, 
    -7.806564, 1.249664, -0.5990295, -3.878708, -4.831841, -0.4459, 
    -1.173225, -2.902649, -6.947197, -4.40242, -2.546944, -2.181061, 
    -3.631592, -6.391983, -8.745911, -9.447739, -9.479507,
  -5.020134, -7.863365, -13.13187, -16.42271, -13.90266, -14.96984, 
    -16.38885, -12.93652, -15.0545, -15.37298, -15.73055, -17.02691, 
    -14.77952, -12.32922, -13.03235, -10.36334, -5.567261, -8.817001, 
    -10.9157, -9.716736, -9.649033, -11.74695, -12.95943, -14.8459, 
    -8.932892, -5.221939, -8.363083, -10.62871, -11.44904, -8.205261, 
    -5.985992, -7.850845, -7.145126, -4.733658, -4.680801, -3.65033, 
    -2.571671, -5.331055, -15.32533, -33.77011, -16.56102, -10.61672, 
    -4.128716, -2.150589, -1.602417, -1.287315, -3.742783, -3.488365, 
    -1.472717, -3.676086, -2.272209, -1.420135, 0.1897888, 1.361664, 
    1.607231, 2.028839, 1.186386, 1.180672, 1.64032, -0.7438126, -2.659981, 
    0.4595413, -3.851662, -8.448784, -12.14645, -14.31986, -15.19928, 
    -8.134705, -2.458405, -4.704224, -8.404495, -4.826904, -0.4605103, 
    0.8853455, -1.562057, -3.39772, -5.228455, -3.263351, -1.565437, 
    -2.620392, -13.27766, -2.708672, -21.24903, -8.47377, -5.72197, 
    -2.780296, -1.102173, 0.5704803, 2.063713, 4.708504, -0.4904404, 
    -2.895119, -1.844078, -4.036797, -4.360207, -3.784424,
  -3.818588, -1.027954, -5.518845, -11.30764, -12.09853, -11.4777, -7.989906, 
    -6.161003, -7.035233, -8.931061, -6.063873, -5.627167, -6.246681, 
    -7.240181, -7.545128, -9.545624, -7.082619, -7.048767, -8.103455, 
    -6.586266, -4.66153, -7.97847, -10.35242, -13.80371, -9.633408, 
    -10.17663, -11.35763, -9.793037, -8.154495, -7.312813, -8.278702, 
    -5.864136, -4.681061, -4.829239, -6.049805, -3.534195, -4.780807, 
    -3.043297, -11.14146, -29.96465, -25.4532, -15.83731, -7.558167, 
    -6.946434, -0.7112885, 1.574913, 1.260063, 0.09156799, 1.634026, 
    1.316582, -0.0003509521, -2.752693, -4.925621, -1.727959, -1.013115, 
    -0.9927979, -2.690453, -2.292534, -0.4865494, -1.267792, -1.98394, 
    -4.772766, -4.20974, -3.550873, -6.536026, -9.668297, -11.19772, 
    -8.956306, -3.147469, -0.8055344, -2.340431, -4.830795, -1.518555, 
    -2.291451, -1.200577, -6.428452, -8.138618, -9.658401, -7.934189, 
    -7.888618, -5.900337, -14.53966, -21.00085, -9.560768, -8.538895, 
    -2.748787, -2.393837, -3.701653, -2.198273, 1.929863, 0.496788, 
    -3.565979, -5.064148, -4.898796, -4.01963, -4.535774,
  -1.041237, 2.055901, 1.310326, -5.380302, -7.233162, -1.08004, -1.570663, 
    -0.1417542, -0.7863007, -3.324043, -0.6964417, 1.096008, 0.0105896, 
    -2.684204, -3.715195, -3.243324, -3.87561, -3.963104, -5.058144, 
    -7.771957, -9.369354, -8.882637, -7.925339, -8.157646, -7.336548, 
    -8.647743, -9.101395, -5.005806, -4.412582, -4.384201, -6.619621, 
    -5.866745, -6.695381, -7.315437, -6.985237, -5.067268, -2.648506, 
    -5.276894, -10.70188, -19.6459, -16.54694, -8.947723, -4.970139, 
    -7.717812, -16.8381, -7.262871, -3.322495, -4.834984, -6.595413, 
    -4.667549, -2.319359, -3.93499, -4.191238, -2.492279, -6.184738, 
    -2.947227, -3.707123, -2.273277, -0.3907318, -1.969376, -4.22509, 
    -2.378479, -4.906609, -8.149063, -6.297745, -4.318314, -0.2964325, 
    -0.4308167, -0.5055542, -2.115974, -2.745132, -2.343575, -5.601883, 
    -7.916229, -6.880814, -8.095657, -8.388878, -7.425865, -5.417015, 
    0.1548615, -0.01412964, -6.679497, -9.968575, -2.637329, -3.799835, 
    -5.413651, -8.136559, -7.193329, -4.973274, -1.535782, -2.234474, 
    -5.146202, -2.97094, -1.159477, -2.686813, -4.097481,
  4.802513, 4.902779, -1.461555, -5.03056, -6.691238, -9.850365, 1.166565, 
    0.8131866, -2.271446, -1.510513, -0.9034805, 0.7751617, -1.509727, 
    -4.276909, -3.871452, -4.418076, -8.029007, -8.521202, -7.708954, 
    -4.811546, -4.251396, -3.982903, -4.757652, -4.717819, -5.001671, 
    -4.316254, -4.441505, -5.338127, -5.45713, -4.625351, -7.227951, 
    -9.63707, -10.5829, -8.148788, -4.663895, -3.97821, -4.859207, -6.455299, 
    -7.456596, -8.153732, -9.575874, -12.44437, -12.08525, -11.1527, 
    -8.940201, -10.29723, -15.21598, -26.88239, -27.09984, -23.25687, 
    -21.64542, -21.67249, -12.41598, -6.736809, -4.433174, -1.913124, 
    0.1668396, 1.14106, 1.151466, -1.894882, -1.975342, -2.145142, -2.425369, 
    -4.929268, -4.623543, 0.3347931, 2.538704, 1.043655, 0.04677582, 
    -1.215973, -0.6956635, -3.540184, -6.497208, -8.211006, -8.455544, 
    -7.80085, -5.94854, -3.913887, -2.538612, -1.170403, 0.935585, 1.173347, 
    -1.13707, -3.745926, -4.188385, -6.326653, -5.165977, -3.662323, 
    -1.187599, -1.703468, -2.792015, -2.874557, -0.3201447, 1.947037, 
    2.379341, 2.996521,
  2.076473, 3.68689, 1.075691, -2.872746, -3.515461, -1.780827, -2.458427, 
    -2.122486, -2.921185, -1.268578, 1.723614, 0.2702217, -2.323528, 
    -3.869102, -1.859993, -1.245911, -1.730812, -4.449047, -6.021446, 
    -4.240974, -3.078735, -3.007118, -3.501656, -4.08239, -4.443054, 
    -4.827431, -5.664406, -7.084721, -8.202171, -7.177704, -6.221718, 
    -8.665199, -9.274826, -7.764412, -5.728485, -5.83213, -6.454269, 
    -7.988907, -9.624329, -9.289948, -10.49541, -12.46156, -11.26806, 
    -9.663109, -9.905304, -12.12483, -15.47691, -16.21103, -15.23681, 
    -11.61702, -9.051399, -7.269096, -6.896202, -6.784485, -5.446449, 
    -4.742012, -4.131332, -1.533157, -2.608162, -3.375881, -3.906078, 
    -2.801388, -1.407124, -1.537071, -1.858162, -0.4271774, 0.3720551, 
    0.5400085, -1.816246, -3.207397, -2.718857, -4.579018, -4.487343, 
    -6.345673, -7.115204, -4.35009, -1.283684, -1.462349, -2.714943, 
    -5.582657, -6.059204, -6.472748, -7.220413, -8.531342, -9.709465, 
    -10.273, -9.672226, -10.56389, -6.853737, -5.789932, -6.837852, 
    -6.003464, -2.575871, -1.982384, -2.988369, -1.903736,
  -0.3685722, 0.1668434, 1.25539, 0.6129417, -1.033939, -2.779251, -5.091755, 
    -7.053471, -8.201389, -6.007378, -3.257122, -5.129265, -5.593327, 
    -5.714413, -7.133408, -5.888371, -5.748009, -5.901131, -6.150871, 
    -4.982643, -4.553478, -4.753994, -5.091751, -4.572472, -3.581326, 
    -3.876652, -4.318317, -5.863373, -5.456337, -4.638111, -5.55608, 
    -7.553474, -8.122223, -8.27483, -7.697742, -8.608681, -10.85374, 
    -11.14149, -11.71154, -12.57248, -12.65295, -12.11884, -10.97405, 
    -9.511288, -10.0355, -11.66858, -12.19437, -12.48239, -11.35582, 
    -11.24828, -10.73031, -10.59358, -10.86285, -8.299309, -6.279255, 
    -3.79332, -3.673519, -3.499561, -2.114666, -0.6042557, -0.6602478, 
    -1.208946, -0.8162346, -1.234203, -1.372223, -1.409725, -2.517548, 
    -4.207394, -5.980831, -7.888893, -8.123531, -6.263897, -4.071712, 
    -3.566765, -4.980816, -5.567551, -5.768589, -5.242546, -4.017548, 
    -3.783157, -4.106865, -4.171974, -5.79644, -8.602165, -11.19566, 
    -12.67639, -12.67743, -12.86728, -10.60739, -8.867798, -9.111294, 
    -9.755035, -11.61883, -10.97534, -3.657116, -0.633419,
  -2.414925, -1.462847, -0.09045029, 1.019966, 1.548872, 0.9564285, 
    -0.2628441, -2.954252, -6.518053, -8.837845, -9.003204, -8.099041, 
    -7.026909, -5.989929, -5.197742, -5.759712, -6.304775, -6.017014, 
    -5.135765, -4.165447, -3.654507, -3.268051, -3.12352, -3.45842, 
    -3.653469, -4.08316, -3.924564, -3.753731, -4.050865, -4.760242, 
    -5.80946, -6.212318, -7.371178, -8.099819, -7.621956, -8.058159, 
    -7.788628, -7.257381, -7.199043, -7.91024, -7.346703, -6.920925, 
    -7.138367, -7.562847, -8.042534, -9.05191, -9.233158, -7.613892, 
    -6.211288, -6.527431, -6.620922, -6.227692, -6.185246, -6.221184, 
    -6.018841, -5.221706, -5.404774, -6.045135, -5.912838, -5.730034, 
    -5.760506, -6.356339, -6.643059, -5.051128, -4.227951, -4.29071, 
    -5.325085, -5.861023, -7.188099, -7.321705, -6.310753, -5.571693, 
    -4.862328, -3.913879, -3.149826, -4.114929, -3.553211, -2.713371, 
    -1.978996, -2.499832, -3.520142, -4.853725, -6.706337, -8.280819, 
    -8.662849, -7.792274, -6.86311, -6.992538, -6.464935, -6.734718, 
    -5.86441, -5.265965, -6.581856, -7.622742, -6.07534, -4.717529,
  -2.794096, -2.680557, -2.470659, -3.101389, -3.720922, -5.105034, 
    -5.574306, -5.904768, -6.252686, -5.462582, -4.430815, -3.375084, 
    -2.24774, -1.728207, -1.608936, -2.106853, -3.02873, -3.927948, 
    -4.563885, -4.241488, -3.700344, -2.795918, -2.433678, -2.406855, 
    -3.228991, -3.83264, -4.199045, -3.759983, -3.846964, -3.668835, 
    -3.72196, -4.051384, -4.1355, -4.130812, -4.489145, -4.688364, -4.710239, 
    -4.67873, -4.595917, -4.394875, -3.819096, -3.783417, -4.237846, 
    -4.603729, -4.389668, -4.040447, -3.592266, -3.456852, -3.253471, 
    -3.093052, -3.078728, -3.263885, -4.404251, -5.138885, -5.527687, 
    -5.439407, -5.190453, -4.894096, -4.636543, -4.730293, -4.322479, 
    -3.808159, -3.712837, -3.541222, -3.209972, -2.257898, -2.389145, 
    -2.697477, -3.263102, -3.873518, -4.136801, -3.778988, -3.614927, 
    -3.408154, -3.285238, -3.079765, -2.763359, -2.784191, -2.53706, 
    -2.193054, -2.493053, -2.971703, -3.4105, -3.269085, -2.884712, -2.59409, 
    -2.097214, -1.740181, -1.827168, -2.498001, -3.21727, -3.302946, 
    -3.463364, -3.570658, -3.519096, -3.418837,
  -2.990973, -3.043057, -3.012589, -2.945662, -2.27613, -1.808159, -1.564152, 
    -1.38238, -1.233419, -1.081076, -1.046963, -0.8263893, -0.5625896, 
    -0.7920151, -1.754253, -2.668839, -3.10738, -3.222223, -3.225609, 
    -3.041233, -2.910765, -2.817797, -2.635244, -2.743837, -3.019358, 
    -2.912066, -3.279774, -3.956078, -4.00712, -4.20035, -4.195139, 
    -3.948265, -3.480293, -3.175606, -2.982899, -2.837326, -2.75321, 
    -2.365711, -1.994356, -1.845659, -1.899303, -1.932379, -1.992016, 
    -1.912067, -1.808681, -2.113367, -2.45295, -2.605553, -2.651648, 
    -2.473263, -2.49618, -2.832117, -3.060762, -3.054514, -2.911804, 
    -2.656336, -2.67795, -2.613628, -2.495659, -2.633419, -2.869356, 
    -2.855555, -2.89019, -2.983158, -3.225605, -3.364408, -3.188887, 
    -2.509722, -2.240713, -2.088629, -2.286808, -2.293839, -2.143316, 
    -2.02092, -2.21545, -2.185762, -1.962847, -1.822222, -1.751127, 
    -1.844095, -1.883158, -1.795918, -1.615971, -1.339411, -0.9529533, 
    -0.7498264, -0.8818588, -1.295919, -1.407118, -1.345139, -1.205034, 
    -1.488632, -1.866234, -2.097225, -2.595144, -2.803736,
  0.4801273, 0.511899, 0.4290867, 0.3277836, 0.2168465, 0.1639824, 
    0.09366989, -0.03263187, -0.1821108, -0.3563309, -0.5826321, -0.7615385, 
    -0.8102369, -0.8737783, -1.008935, -1.114404, -1.133414, -1.271173, 
    -1.449039, -1.635237, -1.745132, -1.787841, -1.707372, -1.571434, 
    -1.484977, -1.455289, -1.289403, -1.160236, -1.082893, -1.069872, 
    -1.054507, -1.027425, -1.102424, -1.158935, -1.195914, -1.1993, 
    -1.149039, -0.9852371, -0.916749, -0.8029461, -0.7349777, -0.7607594, 
    -0.8016443, -0.8328934, -0.8628426, -0.8649263, -0.890708, -0.8453951, 
    -0.7633638, -0.8000822, -0.9469576, -1.018312, -1.187843, -1.303988, 
    -1.355551, -1.417271, -1.527686, -1.686801, -1.709718, -1.729249, 
    -1.670655, -1.787843, -1.922739, -1.956073, -1.932374, -1.859717, 
    -1.839405, -1.812322, -1.697219, -1.594875, -1.492534, -1.343575, 
    -1.422742, -1.632898, -1.791492, -2.063628, -2.132378, -2.159202, 
    -2.217013, -2.158941, -2.067534, -1.95868, -1.737586, -1.551649, 
    -1.392534, -1.312586, -1.229252, -1.055293, -0.8034706, -0.5084181, 
    -0.2258654, -0.02742863, 0.03377151, 0.1551266, 0.3095541, 0.4199705,
  -0.2368019, -0.2295103, -0.2545104, -0.2493019, -0.2599788, -0.2808123, 
    -0.306854, -0.3417499, -0.3761246, -0.416229, -0.4662287, -0.5159688, 
    -0.5524273, -0.5683134, -0.5498238, -0.5016463, -0.4459171, -0.4006045, 
    -0.3722191, -0.3586774, -0.3076358, -0.2451358, -0.1920104, -0.1618023, 
    -0.1612816, -0.1618023, -0.1435733, -0.1360216, -0.1115417, -0.07378149, 
    -0.07143784, -0.0961771, -0.1115417, -0.1157088, -0.1269064, -0.1529484, 
    -0.1688337, -0.2042503, -0.250865, -0.2719588, -0.2935734, -0.2982607, 
    -0.2972188, -0.3013859, -0.3357611, -0.3769064, -0.4232607, -0.4683127, 
    -0.526907, -0.5732608, -0.5951357, -0.6172714, -0.6243024, -0.6209168, 
    -0.6302919, -0.6331568, -0.6250834, -0.6349797, -0.6430521, -0.636281, 
    -0.631073, -0.62925, -0.6477394, -0.6474791, -0.6612811, -0.6597185, 
    -0.6659684, -0.6784682, -0.6951356, -0.6808124, -0.6657081, -0.6758647, 
    -0.6823745, -0.698781, -0.7141457, -0.7164893, -0.7081561, -0.7058125, 
    -0.68576, -0.6802912, -0.6633644, -0.6472187, -0.6222181, -0.5974793, 
    -0.5985212, -0.5888855, -0.5818546, -0.5644062, -0.5214372, -0.4644058, 
    -0.3982604, -0.3659687, -0.3344586, -0.3058128, -0.2922711, -0.2573748,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.009374999, -0.005989581, -0.002343751, 0.002864584, 0.004427083, 
    0.002343751, 0.0002604127, -0.00416667, -0.01666667, -0.02760417, 
    -0.034375, -0.03515625, -0.03906251, -0.04088542, -0.04036458, 
    -0.03723958, -0.03567708, -0.03619792, -0.03020833, -0.02500001, 
    -0.02187501, -0.02135417, -0.01718751, -0.01588543, -0.01848958, 
    -0.01822916, -0.01901042, -0.01822916, -0.02317709, -0.03411458, 
    -0.03854166, -0.04401042, -0.05208333, -0.05833334, -0.05598958, 
    -0.05390625, -0.0515625, -0.04765625, -0.04453126, -0.03958333, 
    -0.03671876, -0.03515625, -0.02864584, -0.01848958, -0.02005209, 
    -0.02161459, -0.01770834, -0.01197917, -0.009635419, -0.0125, 
    -0.01171875, -0.009895831, -0.008333333, -0.00755208, -0.009635415, 
    -0.01015625, -0.01067709, -0.01041666, -0.009635415, -0.0078125, 
    -0.005468752, -0.004427083, -0.002083335, 0, 0.001041669, -0.001041666, 
    -0.004687499, -0.001562499, 0.0005208328, -0.002343751, -0.005989581, 
    -0.007031247, -0.004947916, -0.00416667, -0.0007812455, 0.001562499, 0, 
    -0.001302078, -0.000781253, -0.00390625, -0.006510414, -0.005989589, 
    -0.009374999, -0.01510417, -0.02083333, -0.01614583, -0.0171875, 
    -0.01380208, -0.008593746, -0.009895831, -0.01223958, -0.01041666, 
    -0.01328125, -0.01223958, -0.0140625, -0.01015625,
  -0.06510425, -0.0531249, -0.05234373, -0.06875002, -0.1117188, -0.1796875, 
    -0.2109375, -0.2028646, -0.2236979, -0.2783854, -0.3393229, -0.3882812, 
    -0.3768228, -0.3171874, -0.2742188, -0.2520833, -0.2421875, -0.2419271, 
    -0.2963541, -0.3354166, -0.3106773, -0.3140626, -0.3070314, -0.2796874, 
    -0.2432292, -0.198698, -0.1898439, -0.1434896, -0.1442709, -0.1523438, 
    -0.188802, -0.2101562, -0.2528646, -0.3260417, -0.395052, -0.4390626, 
    -0.4614584, -0.4596355, -0.3382813, -0.2502605, -0.2036458, -0.1934897, 
    -0.1682291, -0.1268229, -0.1054688, -0.08697915, -0.08333325, -0.0645833, 
    -0.08255208, -0.09296882, -0.07395828, -0.03932285, -0.03854162, 
    -0.04609376, -0.01380205, -0.0213542, -0.01197922, 0.01223958, 
    0.02369791, 0.005729198, -0.01015627, 0.01953125, 0.02656245, 
    0.004427075, -0.01953131, -0.0205729, -0.006250024, 0.01015627, 
    0.02447927, 0.02005208, -0.02395833, -0.0164063, 0.02161455, 0.0283854, 
    0.0432291, 0.02734375, 0.0354166, 0.05130208, 0.08255208, 0.1044271, 
    0.09479165, 0.1440104, 0.1221354, 0.07369781, 0.05286455, 0.01744795, 
    -0.0484376, -0.09505212, -0.0588541, -0.04505217, -0.05234373, 
    -0.06015635, -0.06015635, -0.05442703, -0.04036462, -0.05052078,
  -0.205729, -0.3447919, -0.4747396, -0.5773439, -0.6281252, -0.6536455, 
    -0.7013021, -0.7523441, -0.8859372, -1, -0.9911456, -1.125, -1.172135, 
    -1.059114, -1.011458, -0.9338541, -0.6752605, -0.5510416, -0.5236979, 
    -0.645833, -0.7294269, -0.8796873, -0.882031, -0.8677082, -0.6963544, 
    -0.7148438, -0.7111979, -0.7054687, -0.6140623, -0.7039065, -0.7791667, 
    -0.6875, -0.7046881, -0.6911459, -0.5820317, -0.5330734, -0.4442706, 
    -0.5716147, -0.5757813, -0.448698, -0.4249997, -0.4049478, -0.341146, 
    -0.3789063, -0.3700519, -0.4802084, -0.5257812, -0.6976562, -0.8125, 
    -0.5455732, -0.2151041, -0.04817677, 0.0447917, 0.1549478, 0.2679687, 
    0.3479171, 0.3804691, 0.3804688, 0.09375, -0.1481769, -0.4927082, 
    -0.7867186, -0.9450519, -1.014844, -0.8726563, -0.6096356, -0.4023438, 
    -0.2333336, -0.1520834, 0.0348959, 0.1403646, 0.2575521, 0.3218751, 
    0.4247398, 0.4328127, 0.4559894, 0.4820313, 0.4731774, 0.2763019, 
    0.08619785, -0.05546856, -0.1325521, -0.1307292, -0.2010417, -0.2971358, 
    -0.4065104, -0.5645833, -0.6312499, -0.6505208, -0.4640627, -0.3161454, 
    -0.2130208, -0.2463546, -0.3330727, -0.2734375, -0.2286458,
  -1.265885, -0.8528643, -0.5544271, -0.660677, -0.8677082, -1.082553, 
    -1.242969, -1.31927, -1.482813, -1.347656, -1.301561, -1.319011, 
    -1.413802, -1.820572, -2.066406, -1.856251, -1.485417, -1.169271, 
    -1.001822, -0.859375, -1.038542, -1.00026, -0.744791, -0.6645832, 
    -0.6408844, -0.7341156, -0.7210922, -0.8776035, -0.7854156, -0.5950527, 
    -0.608593, -0.6263027, -0.7263031, -0.9442711, -1.130209, -1.111198, 
    -1.107031, -0.9023438, -0.4208336, -0.463541, -0.6760406, -1.131771, 
    -1.20625, -1.186459, -1.00573, -0.3880205, -0.1921873, -0.3369799, 
    -0.2335939, -0.2265625, -0.3119783, -0.9075518, -1.161458, -1.382552, 
    -1.295052, -1.171614, -0.9671879, -0.9000006, -0.9343748, -0.9833326, 
    -1.504427, -2.013542, -2.325521, -2.189063, -1.877344, -1.878386, 
    -1.730208, -1.571875, -1.373698, -1.259895, -1.133594, -1.326041, 
    -1.241145, -1.082552, -1.212761, -1.054948, -0.7059898, -0.4013023, 
    -0.2268229, 0.004687309, 0.05260372, -0.09557247, -0.2046871, -0.3656254, 
    -0.8125, -1.272917, -1.815365, -1.927865, -1.958073, -1.69323, -1.426824, 
    -1.340625, -1.678125, -1.95599, -2.079948, -1.672656,
  -3.540886, -3.654688, -2.429167, -2.073698, -1.920834, -1.765625, 
    -1.151823, -1.113281, -1.439062, -1.86875, -1.974218, -1.141405, 
    -1.345833, -1.902605, -2.696095, -3.054688, -2.820833, -2.219271, 
    -0.9648438, -0.1945305, 0.09401131, -0.7893219, -1.046875, -0.8731766, 
    -0.7934895, -1.203384, -0.7604179, -0.002605438, -0.1929703, -0.7307301, 
    -1.410938, -2.449478, -2.925781, -3.663803, -3.74375, -3.665886, 
    -2.93203, -2.372917, -2.141405, -2.215364, -2.358593, -2.22578, 
    -2.269011, -1.93047, -1.529165, -0.816927, -1.119009, -1.20521, 
    -0.08958244, 0.5997391, 0.6442699, 0.4875011, 0.02031231, -0.2132816, 
    -0.5184889, -0.396615, -0.7757816, -1.191667, -1.355729, -1.372917, 
    -1.638542, -2.55547, -3.00677, -2.917707, -2.743751, -2.030208, 
    -1.533072, -0.6789064, -0.2731771, -0.5848951, -1.564844, -2.786199, 
    -2.952604, -2.657031, -2.636198, -2.748177, -2.394011, -2.140104, 
    -0.7885418, -0.542448, -1.044009, -1.509115, -1.208855, -0.6760426, 
    -0.686718, -0.9893227, -1.649479, -1.520573, -1.108334, -0.7942715, 
    -0.9229183, -1.481249, -2.058073, -2.485416, -2.985937, -3.330208,
  -5.595314, -5.703125, -5.548437, -5.789324, -5.670313, -5.009897, 
    -3.916407, -3.797396, -3.978125, -3.98802, -3.598438, -2.730989, 
    -2.647396, -3.653126, -3.956249, -4.306511, -4.008854, -4.309376, 
    -4.302084, -3.825001, -4.167448, -3.877083, -3.725, -3.56953, -3.225521, 
    -2.43203, -1.070053, -0.002864838, -0.03463745, 0.261198, 0.6158848, 
    -0.04166603, -1.354687, -1.760418, -2.966667, -3.438282, -4.373959, 
    -3.798958, -3.842709, -3.832031, -4.432814, -3.069792, -1.776043, 
    -0.5335922, 0.8466129, 1.596354, 0.6372395, -0.4429684, -0.3098965, 
    -0.3848953, 0.05546761, -0.604948, -0.9927082, -1.140366, -0.6330719, 
    0.002344131, -0.3450527, -1.340887, -2.514584, -2.125, -1.472918, 
    -0.8958321, -1.206772, -2.19323, -1.909897, -1.585938, -1.022917, 
    -0.3833332, 0.3057289, -0.1911449, -1.162239, -1.176302, -0.6611977, 
    -1.174219, -1.369009, -1.502605, -1.312239, -0.7200527, -0.3177071, 
    -1.192186, -2.410156, -3.545053, -3.997135, -3.500261, -3.101563, 
    -3.328384, -3.664583, -4.325001, -4.228127, -4.628647, -5.175001, 
    -5.268749, -5.96302, -5.998438, -6.666147, -6.29974,
  -1.759634, -2.178646, -0.8380203, -0.7953148, -1.182032, -2.946877, 
    -2.135677, -1.388542, -1.984112, -2.090105, -0.3354187, 0.2903633, 
    -0.06015587, 0.4416656, 0.3125, 1.165104, 1.579948, 1.196615, 
    -0.01171875, -1.373178, -2.590624, -2.751043, -1.584373, -0.4932289, 
    0.3822899, 0.1927071, -1.15469, -1.846096, -1.219532, -0.4606781, 
    0.848175, 1.319271, 1.198957, 1.151302, -0.8609371, -0.4690132, 
    -0.4627609, -0.874218, -1.095573, -1.088022, -0.9109344, -2.226303, 
    -2.539583, -2.43099, -1.603645, -0.06692886, 0.05937195, -1.089844, 
    -1.607031, -1.55677, -2.754946, -3.464844, -2.433334, -1.107552, 
    -0.0236969, -0.3372383, -0.7453117, -0.642971, -0.514843, -0.01041794, 
    -1.143749, -1.287762, -1.4625, -1.807552, -0.8320313, -0.9765625, 
    -1.590626, -0.994009, 0.0546875, 1.1138, 1.510418, 1.370575, 0.6299477, 
    0.4526062, -0.7624969, -1.113022, -0.455471, 0.1403656, 0.3669281, 
    -1.355728, -1.98151, -2.451302, -2.190104, -1.683332, -1.639843, 
    -2.438801, -2.778645, -2.482292, -2.641405, -2.500261, -2.653387, 
    -2.311199, -2.335678, -2.966404, -2.616407, -1.592449,
  -0.5924492, -3.063019, -3.609375, -3.371353, -1.56953, -1.222656, 
    0.5473938, 1.040886, 1.152344, 1.95208, 2.451561, 1.788803, 0.9656219, 
    0.125, 0.6333351, 0.2062492, -0.971096, -1.841145, 0.07968903, 1.083073, 
    0.8216133, -0.5161476, -1.178123, -1.288803, -0.6203156, -0.6203117, 
    0.3171883, 0.1403656, -0.9414063, -1.573437, -1.528122, -0.6598969, 
    -0.9755211, -0.9260406, -1.346092, -1.394531, -0.1515656, 0.1591148, 
    -0.6520805, -2.070313, -1.765362, -1.42318, -1.017189, -1.649998, 
    -0.6393242, -0.3567734, -1.433857, -3.327602, -0.9283867, -0.004947662, 
    -0.4794273, 0.02656174, 0.6875, -0.4903641, -1.684372, -2.188541, 
    -1.673439, -0.3062477, 0.3203125, 0.8489571, -0.5450516, -1.584114, 
    -0.6216164, -2.222916, -1.479427, 0.9036446, 0.4739571, 0.6653671, 
    0.1635437, 0.6158867, 0.3507805, -0.05521011, -0.6393242, -0.01614761, 
    0.7697906, 0.4244766, -0.4208336, -0.7471352, -0.3531265, 0.2414093, 
    -1.232292, -0.7075539, -1.379166, -0.2859383, 0.6653633, 0.5598946, 
    -0.5635414, -1.357552, -2.645313, -3.510677, -1.527866, 1.074997, 
    -0.7083359, -4.240887, -4.272137, -1.022915,
  -0.4559898, 1.851563, 2.458332, 1.410934, -0.1565094, 0.5591164, 
    -0.7778625, -0.90625, -1.572395, -0.5903625, -0.1976547, -2.740105, 
    -4.476563, -1.751823, 1.997398, 1.823177, 0.8606796, 0.0234375, 1.920311, 
    2.634117, 1.467186, 1.292709, 2.919533, 3.323696, 0.3994789, -1.265884, 
    1.396614, 1.513283, -0.6976585, -0.08853912, 2.283855, 0.8130226, 
    -0.5528641, -2.170315, -1.590103, 0.8729172, 2.614063, 0.3622398, 
    -1.122654, -0.6507835, -1.494011, -0.5200539, -0.4434891, 0.5921898, 
    -0.9888039, 0.6166649, 1.278908, -0.65625, -0.02760315, 1.498436, 
    2.437763, 2.330208, 2.654686, 2.843491, 1.346352, 1.637764, -0.8294258, 
    -1.371353, -1.429428, -1.379425, 0.5234375, 0.6122398, 1.58802, 
    -0.0942688, -2.429947, -0.3963509, -1.646873, -2.561977, -1.182034, 
    1.239323, 1.379425, 1.681252, 3.802864, 3.83672, 3.853127, 1.239063, 
    0.02057266, 0.3252602, -0.3531265, 0.2583389, 0.5992203, -0.5835915, 
    -1.218491, -0.3208351, -0.6437492, -2.695572, -1.416405, 2.126823, 
    0.3736954, -0.5651054, -0.296875, -0.009895325, -1.522137, 0.2416649, 
    -1.027344, -1.95026,
  3.221352, 2.589844, 3.279427, 2.19323, 3.617447, 3.07058, 2.126556, 
    1.006508, -0.2703171, -0.1841125, 0.5505219, 0.9252625, 0.6395798, 
    -1.245049, -0.2583313, -0.007553101, -0.4351501, 0.2505188, 0.4263, 
    1.412758, 3.362755, 1.311722, 1.258072, 5.721878, 3.390625, 1.240105, 
    2.00573, 0.1054688, -2.055473, -0.609375, 1.654427, -0.1429672, 
    -1.408073, -1.351044, -3.011459, -0.4380264, 0.208847, -1.861717, 
    -2.901558, -0.1281281, 0.7674484, 0.6231766, 4.252342, 4.61615, 2.801826, 
    2.066925, 2.423958, 3.017189, 3.578644, 4.515366, 2.394531, 3.143227, 
    4.851822, 2.72448, 2.482292, 2.15313, -1.301041, -1.449738, 1.629166, 
    1.148178, 0.674736, 0.9221344, 0.1901016, 0.1687546, -0.9523468, 
    -2.212761, -0.5481796, -1.246353, -1.921356, -2.000267, -2.502342, 
    -0.4924469, 1.078392, 0.8979187, 1.119011, 0.8804703, 1.03828, 3.59948, 
    -0.04088593, 1.076828, 3.389328, 1.773697, 0.1052094, -1.054428, 
    -0.1299515, 1.488541, 3.329689, 3.683327, 1.790108, 1.847656, 0.6875, 
    -1.508331, -0.6966171, 2.801041, 1.827347, 1.428902,
  2.465103, 0.6046829, 0.9502563, 1.949219, 1.699478, -2.1763, -0.2950516, 
    3.147133, 2.78125, 0.6145859, -0.3015594, 1.545837, 0.2869797, 1.206772, 
    0.4914093, -1.34687, 1.239067, 4.513016, 3.233589, 1.587502, 2.631248, 
    1.419533, 1.581512, 1.387238, 2.277603, 0.5197906, -2.294533, -2.19088, 
    -2.29792, 2.601563, 3.364059, 0.9523392, 2.149216, 4.332291, 2.307816, 
    -0.8507843, -0.2864609, -0.3692703, 1.017708, 3.678391, 5.053902, 
    1.731766, 2.627083, 3.805466, 0.9906311, 1.649483, 5.628387, 5.753647, 
    2.940628, 3.316925, 3.224998, 4.128906, 7.07135, 4.303131, 0.2070313, 
    2.225006, 0.8395844, 1.873695, 3.525261, 0.4187469, 1.933334, 3.983856, 
    3.065887, 2.081512, 2.508591, 0.8486938, -2.962502, -0.6002655, 
    -0.5585938, -0.2622375, -1.188278, 2.734894, 3.054688, 1.149742, 
    -0.04505157, 1.548172, 2.335938, 2.650002, 0.9440079, -0.6458282, 
    0.07239532, -1.002609, -0.5901031, 2.91198, 5.832291, 3.291145, 4.821617, 
    5.274734, 3.559898, 2.292709, 2.076302, 1.977348, 2.436722, 0.7624969, 
    0.8953171, 4.949745,
  -4.75547, -2.06485, 3.356247, 3.71328, 0.6645813, -0.8247375, -0.5999985, 
    1.435158, 2.216667, 4.216148, 4.983078, 1.899734, -1.173698, 0.4312515, 
    0.6351547, -3.213539, -0.6018219, 1.750259, -1.296875, -0.6565094, 
    -0.3760376, -1.892708, 4.751305, 3.615105, 1.3638, 0.6739578, -0.4885483, 
    1.924736, 2.672653, 3.063805, 2.929947, -0.6398468, -2.263283, 
    0.08802032, 2.464844, -0.2578125, -1.366928, 0.1833344, 3.417183, 
    3.673958, 0.8205719, 1.097397, 1.450516, 2.285942, 3.438019, 3.822136, 
    7.550003, 5.425781, 4.564323, 4.555984, 3.634117, 2.153122, 4.621094, 
    3.587502, 1.579948, 1.827866, 2.407547, 3.277863, 2.770317, -0.731514, 
    1.978905, 3.171356, 0.8166733, 2.850266, 2.836975, 1.613541, 1.592972, 
    1.82135, 0.985939, -0.1080704, 0.1539078, 0.1783905, 0.1888046, 
    0.2721405, 1.253906, 4.841667, 9.63385, 13.51511, 7.012756, -1.737762, 
    -5.738548, -1.8125, 1.162498, 0.9494781, 0.6372375, 3.542969, 2.833855, 
    3.669273, 2.61692, 2.028122, -0.3812485, 1.044792, 5.021355, 1.540359, 
    -0.4570313, -2.042709,
  -0.5208435, 2.329956, 0.7913971, 0.8799438, 3.003906, 1.011978, 1.715881, 
    -0.9250031, -2.869263, -0.2010345, -1.968491, 1.317703, 4.115097, 
    2.846878, 1.014572, 0.6968689, 2.182816, -0.0466156, -0.3255157, 2.5513, 
    1.113541, -1.420578, -2.643219, -2.056, -1.434891, 0.7622375, 2.655197, 
    3.224731, 2.6474, 1.375778, -0.3538971, -0.4403687, 1.044022, -0.4492188, 
    0.1221313, 0.7239685, -3.114578, 2.088272, 3.512512, 3.060158, -2.1698, 
    -3.292709, -2.123169, -1.553909, 0.8010406, 1.047134, 1.071609, 
    -0.3807297, 1.665894, 4.265625, 3.502075, 2.454941, 3.907288, 5.229172, 
    3.426048, 2.095581, 2.295044, 2.915367, 3.184639, 3.14193, 7.962502, 
    5.520828, 3.764839, 3.601563, 3.669014, 2.014061, 1.731255, 2.234894, 
    4.099998, 4.312759, 0.2520828, -1.019272, 4.102608, 5.480988, 3.29245, 
    7.25885, 14.82213, 19.08593, 5.4086, -5.5849, -7.640106, -4.424988, 
    -2.752869, -4.342712, -5.525261, -0.653656, -0.01171875, -2.279175, 
    0.8585815, 2.209633, 2.650269, 1.8078, 0.4768219, -2.209122, -1.434906, 
    -0.7421875,
  1.01355, 2.440887, 0.2867126, 2.673691, 1.063812, -0.8013, 1.879944, 
    -0.8143158, -1.730209, 2.359375, 6.008347, 3.115891, 7.553116, 4.350006, 
    3.041931, -1.590363, -3.124207, 0.759903, -1.678131, -4.412766, 
    -3.653122, -4.114059, 0.4499969, 3.379425, 4.270309, 3.157547, 2.426819, 
    0.5179749, -1.462509, -1.625519, 0.9541626, 2.346344, -3.088806, 
    -2.02916, -7.465637, -6.017715, -3.355194, -2.523178, -5.909897, 
    -5.234375, -10.36458, -9.675003, -6.452591, -2.714844, -1.348434, 
    -0.9953156, 2.833862, 1.95546, 1.986206, 4.226563, 1.507294, 3.657288, 
    3.376053, 4.938553, 1.924484, -0.5231781, -0.2854156, 0.1065063, 2.94635, 
    -0.2786407, 3.752869, 1.880981, -0.3377533, -1.396088, 0.9098969, 
    3.17395, 1.183853, 1.171097, 3.7388, 3.638275, 3.784897, 0.8164063, 
    2.210159, 3.133331, -1.280472, 7.969269, 10.57968, 8.028397, -4.279953, 
    -16.75781, -15.1599, -7.080994, -8.274994, -6.161209, 0.4523315, 
    2.904953, 1.210159, 1.876831, 2.171616, 3.438538, -0.5382843, -1.207809, 
    0.1059875, 2.90834, 2.681259, 1.694794,
  1.386978, 2.364319, 4.263031, 2.561203, -3.014847, -1.907028, 0.6187439, 
    0.1635437, 0.04139709, 2.461716, 2.154419, 0.6890717, 2.770309, 1.596619, 
    5.505203, 7.615356, 3.935425, -0.3000031, -1.817184, 0.6026001, 
    -1.258331, 2.075531, 1.235428, 0.22995, -1.630219, -5.994797, -5.040894, 
    -5.578903, -1.578384, -0.7335968, 0.5604095, -6.63385, -13.57005, 
    -10.7112, -7.806778, -8.714584, -7.282288, -9.822922, -11.27605, 
    -10.36197, -14.76953, -10.925, -2.422653, 0.1851501, -0.1414185, 
    -0.03125, -1.217178, -2.454956, -0.3091125, -2.282028, -0.4182281, 
    1.865891, -1.084381, -3.57605, -4.638794, -3.762497, -0.09375, -2.095047, 
    0.3862, 1.7211, 3.121353, 1.24324, -2.45755, -1.913025, -2.155472, 
    -1.277863, 0.5658722, -0.8203125, 2.948181, 3.171097, -0.4221344, 
    1.324997, -2.44426, -3.058334, -2.707291, 1.548691, 2.213547, -1.009903, 
    -4.016663, -16.09036, -14.4073, -6.171616, -5.909897, -4.462769, 
    -0.4833374, 3.658066, -1.884628, -0.3614655, 4.779694, 3.52681, 3.344543, 
    1.287231, 1.368744, 4.583069, 2.467972, 0.2575531,
  -0.05755615, 1.573959, -1.026306, -10.63515, -1.581238, 4.788803, 4.465363, 
    4.779694, 4.296097, 3.392715, 0.4067688, 0.7054596, 6.702087, 9.140625, 
    2.98204, -0.591156, 4.177078, 1.686981, -0.2640686, 1.984375, 4.567719, 
    3.878387, -1.348175, -3.58905, -5.492706, -1.207291, -4.705994, 
    -5.722916, -2.782547, -4.404694, -6.068481, -9.362762, -16.18463, 
    -10.77136, -6.052078, -9.809906, -9.996613, -10.25755, -9.552353, 
    -10.6151, -11.37917, -1.507034, -1.601303, -1.118484, -5.046616, 
    -3.730469, -6.045563, -5.237762, -2.284378, -0.3768311, -5.755478, 
    -3.959366, -7.794281, -2.721603, -1.755203, 0.9950562, -0.4848938, 
    0.0403595, 1.025513, 0.6828156, 1.614075, -0.2726593, 0.6981812, 
    2.348969, -0.08308411, -0.7859344, 1.335678, 1.487762, -1.296875, 
    -4.434387, -5.597916, -0.05259705, 0.6015625, -1.533844, -3.203384, 
    -0.9039154, -2.700516, -2.901825, -1.818741, -3.372925, -4.23645, 
    7.603394, 6.774994, 2.558853, 1.123703, 3.596878, 2.845306, 4.231262, 
    4.148438, 6.156784, 6.189072, 0.285675, -0.7731781, 1.647919, 1.084625, 
    -2.070313,
  0.4820404, -0.7447968, -2.648956, 0.006515503, 3.440628, 1.001038, 
    -5.429947, 1.74791, 6.495316, 6.151825, -1.303909, 0.245575, 0.4617157, 
    -3.577606, -1.741409, -3.338287, 2.847397, 3.422913, 6.842194, 5.204422, 
    5.076035, 0.8346405, -1.553375, -0.6385498, -4.060669, -1.253387, 
    -3.795303, -1.965897, -0.9528656, -3.015625, -9.769012, -11.40208, 
    -11.85495, -7.525253, -5.781769, -9.853134, -9.645844, -9.075256, 
    -7.926575, -7.00444, -1.223434, 4.329422, -3.839584, -7.563538, 
    -7.633331, -7.228394, -8.446091, -2.245834, -4.837753, -5.042969, 
    -6.481247, -6.392975, -5.272141, -2.306259, -0.4479218, -2.342697, 
    2.307816, 2.030457, 0.8632813, 4.234634, 4.915878, 7.2724, 6.851822, 
    4.060425, 5.359375, 2.565887, -4.756775, -0.89505, -4.069534, -10.42319, 
    -2.783325, -0.8632813, -2.690109, -5.206253, -2.824738, -1.494797, 
    -5.654434, -2.724472, -0.1164093, 3.782806, 4.333328, 7.409103, 3.273697, 
    9.133331, 5.469528, 5.043228, 6.789841, 3.464325, 1.555725, 2.358841, 
    2.790878, -0.8859406, 0.6109467, -3.7724, -0.8351593, -4.991669,
  0.1447906, -3.838287, -3.608597, -2.404175, -2.687241, 0.0627594, 1.995575, 
    2.474731, 1.514847, 5.082809, -4.370834, -2.768738, 1.4552, 0.5880127, 
    3.579941, 0.4700623, 2.829163, 1.239578, 4.875, 2.061966, -0.1572876, 
    0.4015503, 3.153137, 0.1492157, 1.532303, 2.461975, -0.1302185, 
    -0.3541718, -2.88855, -3.786972, -9.673691, -8.842453, -6.686462, 
    -4.950531, -6.10704, -8.291397, -7.423447, -5.005997, -0.3257904, 
    4.390884, 2.748444, -5.731766, -9.133331, -5.9776, -4.123428, -6.832031, 
    -5.879425, -1.944534, -6.090622, -9.462509, -5.533859, -7.012497, 
    -2.779694, 0.4666748, 3.909119, 2.824219, 6.089844, 2.972656, 6.348175, 
    5.535675, 8.371353, 8.489319, 8.772659, 0.6778717, -2.307037, -7.134903, 
    -5.532028, -12.756, -8.860687, -3.688538, -5.892715, 0.4395905, 
    -2.448441, -1.335159, 3.834625, -4.520584, -2.008331, -0.7979126, 
    -4.693237, 1.929688, 2.843231, 1.289581, 0.5505219, 10.47527, 16.59949, 
    16.4651, 7.948959, 7.954941, 7.888275, 1.025253, -4.440353, -1.859634, 
    -5.903381, -5.6698, 0.1458282, -3.670578,
  0.2023468, -0.1687469, -2.858582, -0.8414001, 1.181259, 10.0724, 2.872147, 
    8.564072, 10.25052, 11.49115, 2.395584, -8.689072, -8.855988, 2.263535, 
    2.148438, 1.325775, 1.809891, -1.367706, -1.980209, -3.184647, -1.584122, 
    0.8986969, -4.14296, -3.106522, -0.9973907, -1.048447, -0.5369873, 
    -1.807037, -2.794006, -4.207565, -7.310425, -9.191666, -7.013275, 
    -7.330734, -4.986191, -5.100784, 1.553635, -2.270309, -0.139328, 
    4.197922, -2.976044, -1.663284, -8.295822, -0.09114075, 0.005203247, 
    -8.913803, -8.276291, -7.103653, -10.81509, -7.433594, -2.600525, 
    1.208588, 3.244797, 6.648697, 9.807297, 4.591675, 5.081253, 5.0466, 
    4.607285, 4.695313, 4.605988, -0.1885529, -3.020569, -3.499481, 
    -5.969528, -4.475784, -6.546875, -4.829941, -1.482819, 1.564575, 
    1.351303, 2.203125, 1.320053, 5.888016, 2.253128, -1.178894, 0.2955627, 
    -1.609116, -6.118752, 10.26172, 1.808075, 8.067444, 6.686462, 12.04088, 
    20.31668, 16.19896, 7.517441, 5.714844, 5.220322, -0.0236969, -3.986206, 
    -3.676559, -2.141159, -0.3887939, 1.800003, 1.015884,
  4.101288, -3.882019, -6.82135, -1.510147, -1.830719, 13.22266, 11.93465, 
    12.60625, 20.96875, 12.54219, 10.36693, 0.3929749, -2.949219, 4.181778, 
    2.115875, -1.961975, -7.162491, -8.261459, -3.716141, -4.550262, 
    -3.654419, -4.301315, -3.084381, -3.643997, -5.312241, -1.483597, 
    3.582031, -1.26329, 3.083862, 4.362503, -0.5536346, -0.1411438, 
    -1.433075, -0.5489502, -0.8557434, -0.1195221, 17.57292, -3.375778, 
    -5.875778, 4.130203, -7.302856, -2.958862, -0.6286469, 9.469009, 
    3.036194, -7.382813, -13.92134, -14.80026, -16.95494, -7.885406, 
    -4.188797, 0.3065033, 0.6744843, 7.333084, 7.843491, 6.982544, 2.989059, 
    -2.611191, -2.077087, -1.913284, -2.391159, -0.2960815, -2.307556, 
    -4.683594, -4.050262, -1.057556, -1.127869, 5.117981, 6.460663, 7.520828, 
    10.03671, 9.331512, 8.416397, 7.846344, -1.831512, -6.11171, -4.516922, 
    -11.80416, 8.105469, 13.83749, 9.653656, 15.57422, 13.42239, 12.81224, 
    24.06589, 16.4026, 5.007278, 3.333069, 2.384644, -0.2666626, -2.501816, 
    -1.333847, 2.692703, 1.960159, 2.439056, 3.039322,
  3.034637, -0.9833374, -2.76535, -7.586975, -3.363541, -3.558853, -5.951553, 
    -18.38072, -6.672394, -0.745575, 9.650269, 0.8544159, 2.442963, 4.870575, 
    0.3708344, -3.822403, -7.017975, -6.049744, 0.2885284, 4.915634, 5.0336, 
    2.479156, 2.68515, -2.22084, -3.136978, 1.037491, -0.6656189, 2.7211, 
    3.425781, 1.537506, 6.353912, 4.168488, 0.7596436, 2.558075, 3.745316, 
    6.750793, 9.9198, -6.248444, -1.298706, 8.356522, -1.199219, -3.655457, 
    -1.648697, 2.444, -7.258072, -19.76457, -24.54193, -18.47551, -10.62083, 
    -9.529694, -10.86302, -8.687759, -8.973969, -1.289322, 9.017715, 
    9.904678, 4.535431, 5.032028, 2.750259, 1.212509, -2.093231, -4.435928, 
    -0.6942749, -2.43541, -1.417709, -0.4325409, 2.897659, 4.592712, 
    6.481003, 8.2724, 8.991928, 9.656509, 9.779694, 3.974213, -9.708344, 
    1.231781, 9.933594, 15.58672, 4.97084, 8.45755, 8.21199, 8.080719, 
    13.68228, 11.80782, 23.54662, 16.06406, 5.255737, -3.782028, -3.412491, 
    -4.268234, -6.067703, -7.792191, -4.098953, -0.2502594, 0.07525635, 
    1.177856,
  -0.5437317, -2.640381, -1.173691, 7.495056, 18.73332, 5.789063, -3.021622, 
    -18.7164, -37.32605, -21.47891, -3.492706, -5.404678, -3.665619, 
    -0.5768127, 0.1864624, -2.328888, -1.613556, -1.512756, 0.3278809, 
    0.6513062, -4.348724, -2.038513, -3.532043, -4.112762, -0.8268127, 
    1.433075, 4.149231, 1.482559, -4.125259, -5.597931, -3.360687, -5.520569, 
    -4.045044, 3.076035, 2.550537, 4.006775, 1.353912, 1.471352, 11.04271, 
    4.530991, -7.625, -8.895569, -7.563278, -4.521347, -4.955994, -11.58099, 
    -10.84114, -9.531509, -2.116669, -1.463791, -0.8713531, -3.828125, 
    -5.118744, -2.036728, 0.006240845, 1.553131, 1.955719, 2.489319, 
    1.040894, 5.427597, 2.509369, -3.210144, -2.550003, -2.59375, -0.388031, 
    -1.286453, 1.90416, -3.187759, 0.4513092, -0.1544342, -0.2973938, 
    -3.123184, -4.020325, -4.047913, -3.332809, 2.634125, 5.622894, 8.812241, 
    10.31172, 6.202866, 6.838806, 13.52083, 15.59167, 5.839325, 8.52475, 
    6.345062, 1.430206, -7.000778, -2.798706, -4.231766, 0.7033844, 
    -5.998169, -1.685944, -4.363541, -1.994537, -1.214844,
  -3.095032, -0.9052124, 3.55545, 13.92004, 19.36823, 6.600525, 14.85469, 
    5.019531, -18.43152, -47.70181, -18.21327, -0.5083313, -3.658844, 
    -5.141663, -5.304932, -3.890869, -1.456757, 1.313263, 0.8627625, 
    3.130737, 0.4684753, 2.16745, -0.6882935, -0.6570435, -0.7617188, 
    2.821869, -7.634369, -9.208588, -6.076553, -2.685944, -6.027863, 
    -16.70313, -0.3414078, -1.660416, -0.35495, -7.056763, -17.20052, 
    -19.56068, -10.97838, -20.40027, -18.58801, -13.80989, -8.430481, 
    2.999741, 14.88881, 21.35313, 18.87579, 15.12759, 17.84193, 16.70183, 
    12.95729, 6.269012, 3.17865, -0.3901062, -1.426544, -5.813293, -8.179443, 
    -7.414825, -11.83698, -12.79141, -15.52292, -17.68515, -17.9276, 
    -17.2552, -15.5276, -13.82111, -11.57448, -10.78204, -10.01927, 
    -15.85129, -17.31094, -14.36328, -11.71797, -7.517197, 2.907028, 
    7.623962, 8.180725, 13.13516, 14.74896, 3.255219, 12.79141, 7.166931, 
    -0.3059845, 0.4458313, 2.280991, -4.932297, -5.691406, -0.1026001, 
    -2.048187, -0.2903595, -3.341919, -3.835144, 2.047119, 0.1888123, 
    -1.113281, -3.805725,
  -3.232025, -4.488556, 2.276062, 12.08907, 13.1362, 9.398697, 6.851822, 
    2.713547, 1.635941, -16.85313, -15.74506, 0.7606812, -1.205444, 
    -1.612244, -7.348694, 0.2612, 0.3692627, 1.404175, 0.90625, 3.259613, 
    3.826569, 1.515106, -0.0229187, -1.038513, 1.017181, -5.488281, 
    -21.83231, -7.229691, -2.780731, -5.564056, -16.08281, -8.237244, 
    9.877342, -3.827072, -5.534637, -8.339066, -9.224228, -12.52448, 
    -10.75157, -8.157547, -6.691406, -3.808594, -1.776566, -0.2333374, 
    4.780991, 7.844528, 4.049225, 5.220322, 5.852325, 7.434891, 8.715118, 
    9.527618, 7.454163, 7.937256, 4.795288, -1.772919, -6.057831, -8.313293, 
    -10.20389, -10.38049, -11.79871, -10.24219, -10.80652, -13.30261, 
    -12.12891, -12.99765, -8.752625, -11.48254, -13.39636, -17.02164, 
    -17.72031, -18.49219, -18.63438, -9.091156, -3.143494, 14.27734, 
    13.19791, 7.236984, 10.15547, 4.89296, -0.2645874, 0.5109253, 3.025513, 
    -2.740631, 1.128113, 3.392975, 5.494781, 3.489838, -3.979919, -1.309875, 
    -2.212494, -3.709351, -4.6539, -6.432831, -3.148163, -3.636719,
  7.245575, -2.535919, 4.166138, 18.14375, 12.33646, 7.371613, -3.317703, 
    -1.780472, 0.9776001, -23.32031, -22.00885, -0.7966156, -4.559631, 
    2.958069, 6.547913, 1.878387, -0.06326294, -2.325256, 1.37085, 4.927582, 
    2.960419, 1.087494, -0.9031372, -1.122925, -0.6447754, -8.707275, 
    -10.55911, 11.83333, -6.614075, -7.96405, -8.5289, -1.137238, -9.460938, 
    -7.798431, -5.520569, -6.00676, -3.940887, -6.850525, -2.170822, 
    -1.142731, -6.532532, -5.898193, -10.00365, -8.604706, -8.195587, 
    -5.351288, -5.658325, -7.180725, -4.793488, -5.662476, -2.855988, 
    2.537247, 3.682831, 4.694275, 5.728653, 7.272934, 7.407303, 5.028107, 
    6.018768, 1.056519, 1.271606, -0.2841187, -0.1515503, 0.2669067, 
    -3.232788, -3.234375, -2.642975, 0.001037598, -4.76355, -10.80704, 
    -13.98099, -13.72006, -7.689575, -10.82892, -2.00676, 12.16171, 3.597397, 
    3.174728, 4.993484, 3.902588, -0.4606628, -2.797638, -3.599213, 
    -6.557037, 0.8591309, 1.40155, 2.981781, 0.9265442, 4.67865, 2.080719, 
    0.6825562, -2.284882, -6.252625, -4.890106, 4.255478, 9.303635,
  7.755722, 6.330719, 8.901566, 14.85886, 9.184906, 7.5289, 3.6828, 4.028381, 
    8.768494, 15.7263, 20.01668, 4.795288, 2.023163, 2.320313, 3.249725, 
    5.92865, 7.014587, 3.083099, 3.167175, -2.731506, -7.474762, -7.057312, 
    -3.813538, 2.104431, 1.214325, -2.666931, -5.588806, -0.1575317, 
    -3.129425, -0.6174316, -7.947144, -7.861481, -7.577087, 5.866409, 
    0.6666565, -5.085419, -4.412506, -5.718231, -1.550507, -1.536713, 
    -4.889587, -5.640625, -8.924988, -8.786469, -7.128662, -6.019257, 
    -5.903381, -3.246887, -7.386475, -5.300781, -4.416931, -5.794006, 
    -7.03125, -8, -4.815887, -5.752869, -6.357544, -2.196869, 1.6651, 
    1.481537, 4.997894, 9.764069, 9.307281, 6.117706, 2.189301, 0.0625, 
    0.6828003, -2.1763, -5.424988, -12.02628, -8.996094, -5.354187, 
    -7.299469, -3.506775, 0.8289032, -5.483078, -6.934372, 4.644775, 
    -3.976044, -1.377594, -4.444, -4.144531, -7.822647, -1.0224, 1.908844, 
    3.847137, 3.991669, 7.908066, 2.769257, -6.928131, -2.501282, -19.14063, 
    -10.39481, -5.481506, -1.664612, 2.020569,
  -1.936981, -0.9002686, 0.117981, 2.845581, 3.338013, 3.418762, 5.103363, 
    5.459381, 2.449982, 13.27161, 15.99036, 2.948944, 5.8013, 5.078644, 
    3.18335, 0.2002869, 5.783356, 0.5794373, 0.8471375, -6.717194, -7.680725, 
    -8.354156, -4.063538, -1.915894, -3.589844, 0.1658936, -8.644012, 
    -26.15729, -5.492188, 12.28488, -1.3302, -5.021332, -5.466125, 4.292969, 
    -3.290619, -0.005981445, -9.671631, -6.374725, 1.106262, -1.2099, 
    0.2901001, -0.7692566, -1.0112, -1.918243, -5.083069, -5.995331, 
    0.4966125, 1.36145, -2.843994, -0.1755066, 1.900269, 0.5882874, 
    -3.071869, -10.64972, -8.509369, -7.966675, -1.941147, -2.797394, 
    2.675781, 4.957291, 5.477875, 9.384888, 13.71121, 13.40652, 16.73203, 
    12.74063, 8.275787, -0.4057312, -4.683075, -6.571899, -10.58698, 
    -9.473419, -7.682556, -3.907532, 1.128113, -2.267197, -10.57266, 
    -13.16849, -12.33881, -10.93723, -9.643753, -3.704681, 2.171616, 
    2.915115, 1.915894, 5.730225, 7.689835, 6.676025, -0.473175, -1.217987, 
    -6.572662, -4.449219, -6.104156, -6.045563, -4.477081, -2.786987,
  2.949219, 4.678131, 6.182007, 4.422913, 0.4739685, -0.07550049, -2.3685, 
    -1.766418, -1.363281, 0.1992188, 1.452606, 3.15155, 12.56873, 6.143768, 
    1.505707, 2.123718, 0.3036499, -2.441681, -2.764832, -9.682037, 
    -7.956238, -5.455994, -10.56769, -6.514069, 6.182007, -2.07605, -12.2724, 
    -20.46432, -19.52997, -6.427368, -6.097137, -1.281769, -1.297119, 
    0.7794189, -0.2926941, -0.7156067, -0.7114563, -2.233856, -2.251038, 
    -0.869812, 0.5484314, 0.9580688, 0.06484985, 0.2463684, -4.965881, 
    -5.137756, -3.689301, -2.535706, 0.3502502, 4.621887, 3.21225, 4.722656, 
    -2.874481, -4.779175, -4.934631, -9.687744, -9.735931, -4.340637, 
    3.976303, 5.396347, 8.977356, 12.32344, 17.32394, 15.38101, 11.09793, 
    6.486176, 4.2901, -2.689056, 1.261719, 1.947662, -10.78151, 4.335922, 
    13.40988, -1.0401, -0.7901001, -4.671631, -7.050537, -5.785156, -8.47551, 
    -4.986969, -3.571869, -4.588547, -4.168243, -2.115631, 1.108337, 
    5.068726, 6.77916, 10.41873, 4.874481, 0.7338562, -4.920319, -4.163788, 
    -2.824219, -1.824493, -2.735931, -2.471344,
  0.9286499, 4.428894, 7.407562, 6.877869, 4.934631, 7.780975, 6.155975, 
    2.79245, 2.923462, 6.069, 4.060669, 4.564819, 6.236969, 5.038025, 
    4.286469, 1.049469, 0.6005249, -4.005981, -2.314606, -5.675781, 
    -7.583069, -5.328644, -6.922638, -9.273956, -9.443481, -5.032288, 
    -13.99738, -23.51666, -17.64037, -10.69635, -3.229706, -1.237762, 
    -1.257019, 6.529175, 4.809357, 0.7846375, -0.3744812, -2.889862, -1.4841, 
    1.0112, 2.083862, -1.719513, 0.3351746, -0.1578064, -7.514313, -5.888031, 
    -3.705963, -5.75705, 0.7684631, -2.95755, -0.6804504, 0.1427002, 
    -3.141693, -5.296631, -4.619781, -8.002365, -11.14297, -10.10364, 
    -7.592972, -3.437759, 3.876831, 1.034363, 4.585419, 7.014587, 9.339325, 
    8.82135, 3.06485, -0.1000061, -1.472931, 13.46875, 12.56848, 12.27605, 
    13.97421, -4.033081, -0.5385437, -0.6218567, -0.5513, -2.473694, 
    -5.465088, -4.800781, -4.086182, -6.331787, -0.09817505, 2.533844, 
    -0.8054657, 2.016922, 2.606522, 6.768494, 6.613007, 3.215607, 1.151581, 
    -2.584381, -5.455963, -4.623444, -4.917694, -3.572662,
  -3.488556, 1.771362, 7.466156, 7.859131, 6.880737, 9.462524, 12.72891, 
    7.396881, 5.000519, 6.316132, 7.438019, 8.748962, 8.502625, 5.101837, 
    6.095856, 5.469025, 3.131256, 2.921875, 1.725525, -0.5546875, -3.822388, 
    -5.436981, -5.645844, -8.0914, -10.56198, -13.99924, -8.272156, 
    -16.31799, -27.76822, -20.26016, -7.182022, 2.323441, 1.795303, 
    -1.094009, 4.419525, 2.853638, -0.0942688, -1.478119, -1.798187, 
    -2.232819, -2.476837, 0.9645996, -2.735657, -4.179962, -6.234375, 
    -7.953918, -3.453918, -6.55365, -2.024994, -0.9138184, -3.143738, 
    -3.798706, -6.569794, -9.291138, -8.689041, -8.398178, -8.224487, 
    -5.88829, -8.919006, -6.920044, -2.108078, -2.585693, 4.480194, 4.085144, 
    7.154968, 6.542969, 0.8127441, 2.966156, 1.479156, 14.40027, 13.50365, 
    2.251282, 5.608337, -0.9862061, -3.52475, -2.615356, 2.420837, -6.016144, 
    -4.457031, -1.576294, -2.950531, -2.387482, -2.145294, -7.052094, 
    -6.303375, -2.309906, -2.098419, 2.166931, 3.071899, 6.470581, 6.804413, 
    0.7260437, -3.07135, -3.836182, -7.470581, -6.952362,
  -6.380463, -2.723938, 2.626038, 3.860931, 3.129425, 4.947388, 5.699493, 
    9.03775, 9.934631, 9.655975, 6.847137, 6.568756, 8.5672, 10.77319, 
    8.997131, 9.166687, 11.15363, 12.25598, 8.290863, 3.499725, 1.481232, 
    1.661469, -4.159363, -5.621613, -6.904694, -23.96901, -34.77551, 
    -22.09271, -21.00546, -8.974747, -9.97551, 1.092194, 4.599747, -3.623688, 
    -1.496613, 6.119278, 5.649475, 2.116928, 6.442444, 4.395828, 1.618484, 
    -1.753906, 0.2307434, -3.188782, -1.813293, -3.476288, -3.594025, 
    -6.930969, -5.5625, -3.221344, -1.738525, -3.3638, -3.502869, -5.012756, 
    -6.890106, -1.462494, -4.535156, -1.915375, -2.988281, -3.624741, 
    -3.506241, 0.003112793, 5.913269, 2.36615, 13.49142, 2.614075, -1.6828, 
    -1.087219, 4.442993, 8.934631, 2.341675, 2.237488, 1.532547, 3.769531, 
    5.551834, 2.903381, 2.734619, 0.4669189, -0.4070435, 3.9953, 5.070038, 
    -0.589325, -1.175507, -1.803894, -2.196594, -5.677887, -7.406769, 
    -0.2132874, -2.830963, 2.680725, 11.16977, 2.570831, 1.121368, 
    -0.8091125, -5.950775, -7.934631,
  1.544281, 1.964325, -0.0880127, 3.095825, -0.3682556, -1.296082, 0.3736877, 
    5.880463, 3.678131, 6.397888, 12.55832, 6.8927, 6.532288, 11.9487, 
    19.17502, 16.08127, 18.97342, 26.58881, 26.67291, 11.60312, 8.271606, 
    -0.1112061, -15.38306, -8.742462, -7.647919, -21.25208, -31.10077, 
    -25.32005, -17.32474, -5.590103, -3.889069, -1.291672, -3.373962, 
    -5.410675, -3.492188, 0.3578186, -0.4153748, -0.8364563, 0.04219055, 
    4.007813, 3.246353, -2.844528, -3.019012, 0.8179626, 7.294281, 4.257553, 
    0.2565155, -0.2127533, -3.801544, -4.546356, -3.505707, -6.64035, 
    -8.496628, -5.277344, -7.124481, 0.7200623, -2.479416, 1.835159, 
    1.505737, 0.5783691, 2.050781, 1.073944, 4.579437, 3.213806, 3.669769, 
    4.359894, 3.582031, 4.526031, 2.439575, 6.05365, 8.875244, 11.02708, 
    8.814056, 7.370834, 2.9039, 5.144531, 7.078903, 9.145828, 7.090881, 
    4.194016, 7.395309, 6.550522, 6.303391, 2.712753, 0.306488, -3.741913, 
    -2.039078, -2.149475, -3.664337, 0.6955566, 4.154144, 2.286194, 5.282288, 
    5.649994, 11.29324, 11.62473,
  16.64427, 21.45886, 22.46484, 6.386719, 0.3679504, -1.240112, 4.117706, 
    1.3685, 4.420837, 8.971893, 14.83438, 16.98517, 23.93439, 31.26068, 
    30.85027, 23.86433, 33.1203, 32.6599, 23.36275, -0.06509399, -12.56668, 
    -22.77057, -26.78201, -16.93698, -24.16852, -12.34375, -1.188568, 
    -6.805206, -18.89738, -17.48671, -7.852859, -14.83932, -10.39609, 
    -7.443741, -11.1987, -12.5177, -11.41145, -8.332291, -5.299484, 
    0.2179718, -0.45755, 1.643738, 2.668488, 6.590622, 5.748962, 4.071625, 
    2.952072, 5.356522, 8.820572, 5.796616, -0.974472, -5.619797, -1.798447, 
    -2.074997, -2.547134, 0.6867065, 1.448425, 8.232285, 7.875, 2.189331, 
    2.603638, 4.595047, 4.749985, 2.373688, 6.181519, 9.809631, 10.64481, 
    12.5979, 20.19037, 12.47684, 11.27083, 4.526291, 8.844269, 5.435165, 
    -1.983597, 0.2523346, 0.4846344, 5.725006, 7.867706, 7.552338, 3.367447, 
    6.804428, 5.361465, 5.320572, 3.830475, 8.548447, 2.833084, -1.264053, 
    2.170044, -1.381256, -0.3255157, 3.151566, 0.8489685, -1.337738, 
    10.90417, 20.07422,
  18.77969, 11.08932, 11.04401, 12.63568, 5.181244, 4.280991, 11.73099, 
    8.460419, 10.95677, 4.924484, 4.788544, 10.86952, 15.2047, 14.93073, 
    8.447144, 20.56953, 26.00311, 16.72162, 14.43021, -14.10782, -11.30704, 
    -16.77213, -17.86276, -10.30392, -8.524216, -14.131, -7.862228, 
    -4.849213, -9.382553, -11.15704, -12.79688, -14.06509, -7.248703, 
    -6.067963, -9.008591, -9.405716, -2.886719, 1.645844, -5.855209, 
    -2.761719, 1.823425, -2.057816, -1.077347, 3.651306, 2.604172, -3.026825, 
    -0.3703156, 1.516144, 4.354691, 8.540634, 1.588272, -1.217194, 0.9377594, 
    -1.601044, -1.166931, 0.514328, 5.436203, 3.815369, 6.305984, 7.403915, 
    5.117188, -1.860672, -6.546875, -10.98386, -8.137253, 6.502335, 
    -0.9138031, -1.009369, 18.77682, 21.75235, 15.43541, 4.894531, 7.468216, 
    -0.657547, -8.893753, -4.671341, -2.920837, 2.215378, 3.9599, 4.31015, 
    4.416916, 2.210938, -4.933853, -5.203125, 0.671875, -0.8653564, 1.438019, 
    0.0630188, 1.311981, 2.88829, 1.746353, 5.827866, 8.703644, 9.657303, 
    11.6414, 15.56563,
  8.871353, 1.442963, 6.682281, 13.33307, 3.484894, -1.190887, -3.437241, 
    7.785416, 10.56354, 5.161194, 0.6169281, -16.4086, -9.865112, 4.754166, 
    7.920822, 7.433334, 9.352097, 11.93854, 2.747925, -3.346344, -3.295044, 
    -10.83673, -12.02708, -3.864304, -3.764587, -6.669525, -8.206512, 
    -8.789337, -10.93152, -11.75911, -13.30754, -3.641922, -4.137756, 
    -4.730209, 1.885666, -1.639847, -1.866669, 3.747391, -3.970062, 
    -9.577866, -3.454941, 0.07759094, -2.015106, -0.9739685, -0.7976532, 
    -2.821609, 0.3119812, -3.133331, -9.691147, -2.836716, -1.680481, 
    -5.093491, 1.216415, 0.65625, -1.200775, 1.07605, -2.325775, 0.5762939, 
    3.963028, 2.152603, -2.101303, -1.263275, -5.863281, -17.42317, -27.4052, 
    -28.41173, -23.04636, -11.25677, -3.1138, 3.740097, 2.638535, -5.911453, 
    -11.51355, -10.90234, -3.964584, -5.475525, -12.2599, -8.952087, 
    -1.367706, -6.264328, -8.835419, -10.45494, -9.948959, -8.670303, 
    -3.207031, -3.823441, -2.619003, -1.011978, -5.180984, -1.413284, 
    3.016922, -1.523178, -1.800781, -0.2846375, 11.24739, 16.06406,
  -8.286728, -7.362244, -0.6781158, -10.53046, -10.5013, -14.03958, 
    -19.02057, -8.7323, -0.7565155, 2.735687, -4.721603, -12.63255, 
    -15.36224, -9.489059, -7.443756, -11.39322, -9.681, -2.673965, -5.920044, 
    -8.760681, -12.27629, -11.39375, -6.728378, -7.355988, -11.98412, 
    -15.44376, -12.9276, -12.02631, -5.363022, -2.276031, -0.33255, 
    -1.777603, -4.565109, -5.183075, -3.046097, 0.9979248, -0.9080811, 
    1.520844, -1.366409, -11.66927, -8.47995, 3.281769, 3.284103, -1.722137, 
    -2.415878, -1.130478, 1.086731, -1.680206, -3.4935, -0.7630157, 1.528381, 
    2.513275, 5.048172, 2.622147, 0.4729156, 4.110687, 2.648697, 6.230209, 
    4.886459, -0.14505, 0.6507721, -3.018234, -8.183853, -20.90521, 
    -32.77396, -33.64766, -21.51588, -6.717972, -6.724213, -13.07396, 
    -13.01251, -15.51979, -16.85365, -12.59166, -9.94635, -12.27396, 
    -16.65312, -20.92604, -19.9151, -19.85963, -9.9552, -6.115631, -8.813034, 
    -12.53073, -5.855209, -8.818497, -13.59584, -10.50182, -12.84557, 
    -10.22266, -1.538284, -0.1468658, -2.669266, -5.231003, -4.463547, 
    2.719543,
  -4.889847, -13.4151, -16.8552, -14.30026, -8.003387, -6.555222, -13.91199, 
    -18.55026, -15.93359, -13.51796, -9.40155, -10.41328, -6.181, -5.15181, 
    -9.214325, -7.373169, -3.9039, -3.164841, -1.85051, -1.410934, -4.342178, 
    -10.64844, -18.87891, -17.52786, -14.04871, -13.64453, -12.81094, 
    -12.13385, -6.188019, -2.255737, -7.541656, -9.125, -7.521103, -6.256516, 
    -4.842438, -1.184113, -2.579956, -3.699219, -29.1151, -28.07344, 
    -13.58594, -10.52499, -9.072662, -6.757813, -3.048431, -2.272659, 
    -1.196091, -0.7718811, 4.005722, 1.326035, 1.79454, 1.9776, 1.655472, 
    1.354431, 5.653381, 4.900787, 5.2453, 1.500259, -5.379425, -2.518234, 
    2.977081, 0.3166656, -11.60677, -20.9539, -18.05624, -22.36145, 
    -15.28438, -13.84401, -15.72345, -15.369, -21.45105, -14.49583, 
    -14.08022, -9.091934, -15.90443, -22.49609, -21.36406, -16.25259, 
    -15.24609, -12.75417, -13.22708, -3.639587, -17.30338, -9.944794, 
    -9.762772, -13.41173, -14.12656, -12.36198, -8.901566, -6.395325, 
    -7.62735, -4.320053, -2.226563, -8.173447, -5.773697, -1.734375,
  -1.70105, -8.546875, -9.321625, -16.72499, -18.34427, -17.02318, -11.73698, 
    -15.444, -14.81041, -12.68959, -13.26485, -19.80391, -17.70183, 
    -9.119797, -2.764069, 0.390625, 1.916916, -0.7674408, -2.501556, 
    -5.272919, -4.945831, -8.669006, -9.042709, -11.4073, -13.02473, 
    -10.7448, -8.979431, -12.04765, -11.52943, -8.694534, -7.853394, 
    -9.124481, -4.336456, -3.844788, -5.060425, -2.233337, -6.591141, 
    -7.073959, -27.63672, -28.34686, -10.84167, -10.89818, -6.541672, 
    -2.479431, 0.79245, -0.2960815, 0.9976654, 0.3653564, -3.500519, 
    -4.017456, -2.041153, 1.3125, -2.996613, -0.283844, 4.009125, 7.249481, 
    6.53775, 2.092972, -1.851822, -7.605209, -6.427856, -8.047134, -13.86171, 
    -9.82135, -3.563019, -4.673965, -9.655212, -13.81485, -14.04453, 
    -9.654953, -9.303909, -9.324478, -8.282806, -13.0862, -12.89246, 
    -23.85625, -15.68698, -8.483322, -0.8828125, 2.061203, 4.589066, 
    -13.65416, -17.59401, -1.924469, -6.300262, -1.639328, 0.0700531, 
    -0.005737305, -1.791412, -0.1882935, 1.540359, -4.627075, -10.5125, 
    -8.751038, -3.25, 2.208603,
  -9.296616, -16.62448, -18.75259, -25.09479, -23.47292, -9.936722, 
    -9.092178, -21.75365, -16.85912, -11.76146, -10.92343, -10.56563, 
    -8.793488, -13.58464, -9.022141, -9.775269, -9.418762, -7.424484, 
    -3.17421, -5.495575, -9.713547, -11.14505, -13.25781, -13.20677, 
    -13.49141, -8.652344, -6.716934, -8.003647, -14.02682, -14.13437, 
    -6.665619, -3.803375, -3.911194, -9.269791, -11.76563, -7.328125, 
    -7.428909, -4.113022, -23.09818, -27.42915, -17.77605, -9.391403, 
    -4.682297, -0.0721283, -7.7164, -5.007034, -7.150269, -8.386719, 
    -13.74348, -17.22369, -8.839325, -6.241928, -5.994003, -5.858597, 
    -9.179428, -1.25676, -0.7570343, -2.282562, -6.715881, -8.78801, 
    -15.57708, -10.77448, -6.988281, -4.080994, -1.164322, -3.941406, -9.125, 
    -14.18698, -12.65599, -7.809372, -2.501572, -3.645309, -8.498962, 
    -10.51511, -13.76094, -12.50626, -10.62709, -6.639832, -1.053131, 
    0.1835938, -1.312759, -10.52344, -6.561966, 1.616928, -2.844269, 
    -0.5729218, 1.402863, -0.9033813, 0.7981873, 3.17865, 0.223175, 
    -3.296616, -2.387238, -3.082291, -2.457031, -2.262238,
  -10.42787, -12.06953, -24.19427, -22.71693, -18.72397, -13.90547, 
    -17.97527, -19.31354, -19.30469, -16.03438, -12.34038, -11.72421, 
    -14.5961, -8.146103, -6.574478, -8.010406, -9.308853, -8.34375, 
    -9.069794, -10.01848, -8.807297, -9.786713, -9.563019, -11.27657, 
    -12.51483, -8.999207, -8.244263, -7.663803, -9.042709, -7.537231, 
    -4.996353, -3.879684, -8.875259, -13.95833, -12.98882, -10.19218, 
    -8.916931, -2.933853, -2.369781, 1.542175, 5.851563, 2.904938, 1.1026, 
    1.949219, 0.8825531, -4.052856, -9.664322, -45.60963, -41.18489, 
    -36.59845, -34.79297, -32.6086, -24.38177, -21.79089, -16.58281, 
    -10.38907, -8.329163, -7.326042, -6.277863, -5.457031, -8.859116, 
    -5.694534, 0.579422, 4.448181, 3.057297, 0.6455688, -1.58255, -4.91095, 
    -10.99245, -11.17787, -7.611984, -6.88855, -6.22551, -9.321106, 
    -11.34193, -11.19974, -6.86171, -2.523697, -5.896347, -4.3638, -5.154694, 
    -9.1315, -8.588272, -4.580994, -5.484634, -3.50209, -4.419266, -1.865356, 
    -1.659637, -0.901825, -0.2359467, -2.209366, -4.919281, -4.328903, 
    -4.538528, -8.117447,
  -3.583336, -5.355988, -7.666153, -12.7815, -14.39011, -14.60625, -18.03308, 
    -20.51353, -15.61953, -12.68802, -14.44818, -14.08229, -16.68724, 
    -14.97448, -8.500519, -8.74791, -5.981766, -3.250778, -1.775009, 
    -3.802078, -3.99115, -7.27655, -8.596619, -9.029175, -7.498428, 
    -8.057281, -8.884888, -7.969528, -5.875519, -6.424744, -6.442719, 
    -7.552078, -10.65234, -11.06509, -8.373444, -4.938019, -2.900772, 
    -5.064331, -3.929428, -1.101822, 0.9554749, 1.005737, -0.0398407, 
    -3.083603, -4.451553, -6.717712, -10.27344, -14.05209, -16.12396, 
    -18.41978, -20.61719, -20.97292, -21.82761, -17.20157, -13.70313, 
    -11.65077, -8.588547, -4.4888, -1.219788, 1.020828, 2.434113, 2.603653, 
    5.703644, 3.222656, -1.001816, -2.056244, -0.6085968, -2.561203, 
    -4.304169, -3.414063, -3.564835, -4.869537, -2.443222, 0.3291626, 
    -1.721344, -1.648956, -5.271622, -6.088547, -5.87944, -7.110931, 
    -6.616928, -7.265625, -7.889832, -6.257034, -2.363815, 0.8765564, 
    1.209625, -4.808853, -5.116142, -4.589066, -6.792709, -9.391151, 
    -4.681511, -3.331253, -4.825783, -3.608337,
  -2.256775, 0.2442703, 2.552345, 2.244011, -0.0687561, -3.868225, -7.60495, 
    -10.08881, -9.247391, -8.46328, -10.76145, -17.68385, -13.82396, 
    -10.32344, -7.473961, -8.62162, -3.664841, 1.787491, 3.629425, 0.2445374, 
    -4.226822, -5.6875, -5.780472, -5.428383, -6.402603, -6.515884, 
    -7.667969, -7.2388, -5.237503, -1.899994, 0.3341141, 0.0158844, 
    -3.942963, -4.501297, -5.340103, -8.744278, -9.520317, -10.75703, 
    -10.0849, -8.136192, -6.019279, -4.185936, -3.741402, -6.046356, 
    -11.40808, -14.25859, -16.30833, -16.62031, -15.27265, -14.71198, 
    -16.00989, -16.11328, -16.86928, -11.73126, -8.232819, -4.476822, 
    -1.260422, -1.774483, -1.338287, -1.632813, 2.859909, 2.436203, 1.672653, 
    0.8703156, -1.777863, -5.165619, -7.578384, -6.258331, -3.093491, 
    -6.217972, -7.657806, -12.2849, -11.5052, -8.673431, -6.119003, 
    -4.956253, -5.21666, -5.500778, -4.662506, -3.124741, -2.464844, 
    -3.41745, -2.259109, -0.5078125, -2.892715, -4.300003, -4.428131, 
    -5.698959, -7.103653, -8.93959, -9.511459, -10.56902, -15.91979, 
    -18.82369, -3.319267, -2.392708,
  -7.296089, -5.145836, -2.585938, -1.290367, -1.095833, -1.191147, 
    -3.089584, -6.248177, -13.99062, -21.72734, -24.40573, -21.09089, 
    -12.61797, -6.626312, -4.892975, 0.2052078, -1.217194, -4.733589, 
    -8.712502, -11.81875, -11.9987, -11.07343, -10.52032, -9.942451, 
    -8.612244, -9.498436, -9.647911, -6.959114, -6.530212, -4.096619, 
    -1.738541, -0.8031235, -4.197395, -5.68177, -5.392708, -9.369781, 
    -10.78932, -10.43959, -10.25105, -11.58724, -11.24506, -11.68359, 
    -13.04817, -14.00807, -14.13229, -12.73386, -11.5737, -11.10338, 
    -9.467712, -7.75, -8.719269, -9.813293, -11.17058, -12.11641, -13.08932, 
    -12.20988, -11.38594, -11.50755, -11.82005, -12.24115, -11.09634, 
    -8.853394, -8.946091, -6.482552, -8.869537, -8.500778, -8.133072, 
    -7.430473, -8.802345, -9.452866, -8.638802, -7.999474, -7.431778, 
    -4.424995, -3.090881, -3.537239, -4.96875, -6.033081, -9.195053, 
    -8.700012, -5.498688, -4.340637, -4.167709, -4.299469, -6.718231, 
    -8.350769, -7.9888, -7.692719, -8.271088, -8.943222, -11.26563, 
    -14.67551, -17.43568, -14.64818, -13.69219, -13.40911,
  -12.1961, -9.796875, -8.04245, -8.004173, -8.333595, -12.64973, -14.03307, 
    -12.45235, -12.96068, -13.88932, -14.79453, -13.52213, -11.6823, 
    -8.426819, -7.497658, -6.5224, -5.309113, -5.241928, -5.563545, 
    -6.775002, -7.402344, -8.078384, -7.83802, -7.989326, -7.109634, 
    -4.858856, -5.032547, -4.328903, -5.919792, -6.276299, -5.556252, 
    -5.390366, -5.110153, -4.961716, -4.862755, -5.0737, -6.160934, 
    -6.995834, -7.682549, -7.887764, -7.651299, -8.001564, -7.950783, 
    -7.358078, -6.095573, -5.251564, -4.751823, -5.300255, -7.505219, 
    -10.52735, -12.97838, -14.87734, -16.39922, -16.73516, -15.94296, 
    -15.28907, -15.3974, -15.12396, -14.43359, -14.66901, -15.69245, 
    -17.00755, -16.63515, -15.43671, -13.47657, -7.887238, -6.799225, 
    -7.311981, -10.44662, -13.54818, -14.57734, -13.76563, -12.07864, 
    -9.462761, -6.401566, -4.343239, -3.057281, -2.290359, -1.160942, 
    -0.3953171, -0.1658859, -0.4450531, -0.8531342, -0.4359436, 0.6968689, 
    -0.7640686, -3.086456, -5.953384, -8.809387, -11.44609, -12.93021, 
    -12.94661, -12.23646, -10.84792, -8.713539, -10.05052,
  -6.156776, -7.808853, -10.12526, -12.19453, -10.85989, -10.77422, 
    -10.74401, -10.97448, -10.25104, -9.527603, -9.457031, -9.438019, 
    -9.701302, -9.610939, -9.724739, -9.902344, -10.33489, -10.90755, 
    -11.59557, -12.07214, -12.56823, -13.45964, -13.90912, -13.79297, 
    -13.16406, -13.03255, -12.39714, -11.80782, -10.12917, -8.148438, 
    -6.710159, -5.56797, -4.486198, -4.255211, -4.556511, -5.130203, 
    -6.094269, -6.501045, -7.048439, -7.716927, -8.372658, -9.133072, 
    -9.072914, -8.694534, -8.0625, -7.763023, -8.223183, -9.78125, -10.88021, 
    -11.8263, -12.39817, -12.77734, -13.36641, -13.34193, -13.59869, 
    -13.92031, -14.86589, -15.69479, -15.61328, -15.38881, -15.73463, 
    -15.49661, -13.9513, -12.5086, -10.8888, -9.364059, -8.17865, -7.515106, 
    -6.448174, -6.170052, -6.819275, -6.586716, -5.796875, -4.972397, 
    -3.311722, -2.271873, -0.9893188, -0.6869812, -1.199738, -2.587761, 
    -4.361977, -5.476303, -5.397919, -4.427086, -3.719795, -3.70755, 
    -3.174217, -2.857033, -4.046875, -5.782555, -6.632813, -6.168755, 
    -5.805206, -5.060158, -5.034897, -5.526039,
  -6.484901, -6.569794, -6.722916, -6.721092, -6.43412, -6.036453, -6.23542, 
    -5.960678, -5.037498, -4.533073, -4.288284, -4.38073, -4.508072, 
    -4.732292, -5.634636, -6.707809, -8.046616, -8.810417, -9.085419, 
    -9.418228, -9.415367, -8.967186, -8.296356, -7.522392, -6.658859, 
    -6.054428, -5.330208, -4.616661, -4.143494, -3.930984, -3.97187, 
    -4.392708, -5.148438, -5.981773, -6.571358, -7.367706, -8.516663, 
    -9.554688, -10.64193, -11.57135, -12.55469, -12.97162, -13.17265, 
    -12.86719, -12.06589, -11.25677, -10.35599, -9.511719, -9.115364, 
    -8.797913, -8.522392, -8.718491, -9.254166, -9.852348, -10.66745, 
    -11.68932, -12.89948, -13.64401, -13.97395, -14.28854, -15.3263, 
    -16.47656, -17.37292, -17.46797, -16.93568, -15.73828, -14.66485, 
    -13.31536, -11.99609, -10.94714, -10.35313, -10.14792, -9.85833, 
    -9.762497, -9.564316, -9.224739, -8.980469, -8.642181, -7.9151, 
    -7.589844, -7.739319, -7.888535, -8.265884, -9.001305, -9.31823, 
    -10.23125, -10.52917, -10.03281, -9.597916, -8.862495, -7.540108, 
    -6.500778, -5.927078, -5.933853, -6.188278, -6.40078,
  -8.478386, -8.593483, -8.728905, -8.912506, -9.101044, -9.312759, 
    -9.624474, -9.848175, -9.88932, -9.874481, -9.858337, -9.874214, 
    -10.03984, -10.08334, -10.09661, -10.2151, -10.26406, -10.15755, 
    -10.03385, -9.764847, -9.522919, -9.236458, -9.008072, -8.792709, 
    -8.385414, -8.145836, -8.180206, -8.302086, -8.470573, -8.620567, 
    -8.851822, -9.171097, -9.552605, -9.843224, -10.24792, -10.60078, 
    -10.95833, -11.27891, -11.48385, -11.45729, -11.29375, -10.93776, 
    -10.68984, -10.53958, -10.23463, -9.881508, -9.66198, -9.416145, -9.1474, 
    -8.846611, -8.708076, -8.657036, -8.524483, -8.45443, -8.507813, 
    -8.448181, -8.437241, -8.323959, -8.278908, -8.287758, -8.360931, 
    -8.352089, -8.407814, -8.340363, -8.414322, -8.276039, -7.997139, 
    -7.769531, -7.587761, -7.462234, -7.380203, -7.290619, -7.383331, 
    -7.383339, -7.354942, -7.234116, -6.863281, -6.542969, -6.30912, 
    -6.181511, -6.120308, -6.231773, -6.287498, -6.446358, -6.725517, 
    -6.961197, -7.31562, -7.592712, -7.823952, -8.003128, -8.110939, 
    -8.231255, -8.309372, -8.357292, -8.392708, -8.439583,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.03020833, -0.01692708, -0.01770833, -0.009635419, -0.009375006, 
    0.005468756, 0.01145834, 0.01015626, 0.001041666, -0.009375006, 
    -0.003124997, 0.004687503, -0.007031247, -0.009635419, -0.01197916, 
    -0.007552087, -0.0109375, -0.01666667, -0.01848958, -0.01875, 
    -0.03020833, -0.03723958, -0.03645833, -0.03723958, -0.03385416, 
    -0.01822917, -0.01197918, -0.009635419, -0.003385425, -0.01276042, 
    -0.01015626, -0.006510422, -0.0002604276, -0.01276043, -0.01953125, 
    -0.0203125, -0.01692709, -0.02291667, -0.01718749, -0.01796874, 
    -0.01901041, -0.02500001, -0.0294271, -0.03567708, -0.04713541, 
    -0.03854166, -0.02838542, -0.03281249, -0.03645833, -0.03489583, 
    -0.03359374, -0.03072917, -0.009635419, -0.01015625, -0.01302083, 
    -0.015625, -0.01119792, -0.0109375, -0.002083339, -0.007031247, 
    -0.01145833, -0.01927084, -0.01354166, -0.01328125, -0.008593753, 
    -0.005208336, -0.002864584, -0.0078125, -0.009114586, -0.003124997, 
    0.001562499, 0.009114586, 0.009114586, 0.003385417, -0.000781253, 
    -0.00364583, -0.01041666, -0.01223958, -0.01770833, -0.01276042, 
    -0.0109375, -0.00416667, -0.01119791, -0.007552087, -0.003125004, 
    -0.01145834, -0.02630208, -0.02760416, -0.02421875, -0.02187499, 
    -0.02395833, -0.01197917, -0.004687503, -0.006510414, -0.01536459, 
    -0.03307292,
  -0.1593751, -0.2565104, -0.2127604, -0.1395833, -0.04088533, -0.005989552, 
    -0.003385425, -0.07864583, -0.0830729, -0.078125, -0.0419271, 0.0119791, 
    0.01822913, -0.1354166, -0.2320312, -0.165625, -0.1205729, -0.06562495, 
    0.008072853, 0.01901042, -0.0505209, -0.1101562, -0.1002604, -0.10625, 
    -0.1567708, -0.1296874, -0.09401047, -0.06484377, -0.03880215, -0.048177, 
    0.05026042, 0.04661453, 0.06901038, 0.07786465, 0.04713547, 0.0703125, 
    0.0760417, 0.0817709, 0.07473958, -0.02682292, -0.06588542, -0.02265632, 
    -0.04999995, -0.1091145, -0.0760417, -0.1200521, -0.1158854, -0.08567703, 
    -0.09427083, -0.1101563, -0.08671868, -0.0348959, -0.0197916, 
    -0.04166675, -0.08333331, -0.1338542, -0.1226562, -0.1111979, -0.1257812, 
    -0.1549479, -0.1614584, -0.2093749, -0.2684896, -0.2544271, -0.2872396, 
    -0.2536459, -0.2601563, -0.2518229, -0.3203124, -0.3273438, -0.2817708, 
    -0.2291667, -0.171875, -0.1895834, -0.2572917, -0.2507813, -0.2158854, 
    -0.1692709, -0.1169271, -0.05286461, -0.02968752, 0.03359377, 0.04505217, 
    -0.01510417, -0.05442703, -0.02109385, -0.0966146, -0.109375, -0.1645833, 
    -0.2346355, -0.2497396, -0.2309896, -0.1716146, -0.1268229, -0.1403645, 
    -0.1703125,
  -0.8453128, -1.105729, -1.374479, -1.067188, -0.9502604, -0.686198, 
    -0.7309897, -0.6255209, -1.058854, -1.094271, -0.6507812, -0.4380207, 
    -0.6091144, -0.9679687, -1.339062, -1.250781, -1.103646, -1.182292, 
    -0.9966145, -0.9291668, -0.8375001, -0.8664064, -1.053125, -0.8908854, 
    -0.5877604, -0.7018232, -0.6585941, -0.5947914, -0.4945312, -0.3721356, 
    -0.1304684, -0.1609373, -0.01744795, 0.1403646, 0.1294274, 0.1489587, 
    -0.2247396, -0.3901043, -0.5997396, -0.711719, -0.7132812, -0.5994792, 
    -0.3786459, -0.2687497, -0.120573, -0.151823, -0.5080729, -0.542448, 
    -0.3695309, -0.1455729, -0.1140625, -0.2408853, -0.4375002, -0.5403647, 
    -0.5414062, -0.5341144, -0.6278646, -0.5882812, -0.6304686, -0.514323, 
    -0.576823, -0.5268228, -0.4908855, -0.5601561, -0.5317707, -0.3414063, 
    -0.1135416, -0.06718755, -0.5018229, -0.7794273, -0.45, 0.0789063, 
    0.1544271, -0.153125, -0.05989575, 0.0739584, 0.03671885, -0.1322918, 
    -0.4429688, -0.3419271, -0.2408857, -0.4390626, -0.5661461, -0.4981773, 
    -0.5197916, -0.4057293, -0.5445316, -0.8184896, -1.014063, -1.028906, 
    -0.9828124, -0.9502604, -0.9567707, -0.963021, -1.050781, -0.871094,
  -1.261198, -0.9549484, -1.085677, -0.8380213, -0.6325521, -0.4184895, 
    -0.6335936, -1.000521, -0.8445311, -1.010156, -0.5346346, -0.0119791, 
    -0.03072834, -0.1494799, 0.2171869, -0.07760429, -0.5778646, -0.8374996, 
    -0.7726564, -0.5645828, -0.5216141, -0.9257813, -0.8507814, -0.3726559, 
    -0.07942772, -0.06223965, -0.05546951, 0.02838516, 0.07291603, 
    -0.1617184, 0.002083778, 0.3143234, 0.7333331, 0.8018231, 0.7255211, 
    0.667448, 0.2859373, -0.4914055, -0.5716143, -0.411458, -0.380208, 
    -0.6851563, -0.5992184, 0.1369791, -0.1263018, -0.4807291, -0.3492193, 
    -0.006249428, 0.177084, -0.1557293, -0.7859378, -0.7104168, -0.3708334, 
    -0.2843752, -0.3976564, -0.6507816, -0.9453125, -0.895834, -0.4015627, 
    -0.05677032, -0.202343, -0.9856777, -1.25703, -1.015365, -0.6117182, 
    -0.02916622, -0.1700525, -0.1895828, -0.3585939, -0.369791, 0.5018234, 
    0.5442715, 0.04843712, -0.1223965, -0.1059895, 0.1885414, 0.4718742, 
    0.4744787, -0.04557228, -0.1216145, -0.1195316, -0.08359432, -0.5010424, 
    -0.6388025, -0.04296875, -0.4963541, -0.8708334, -1.178125, -1.71276, 
    -1.21302, -0.9177084, -1.358593, -1.757292, -1.396355, -0.9317713, 
    -1.415626,
  -1.307812, -0.3567715, -0.09322929, -0.9260416, -0.4497395, 0.594532, 
    0.3682289, -0.1968746, -0.09192657, -0.08619881, -0.08437538, -0.6973953, 
    -0.1617184, 0.3322926, 0.7533855, 0.4179688, 0.4578123, -0.03802013, 
    -0.5330715, -0.2708321, -0.4536457, 0.3729153, 0.3283863, -0.04843712, 
    -0.4890623, -0.4442701, 0.3140631, 0.452343, -0.353385, -0.9447908, 
    -0.6184893, 0.1309891, 0.3473969, 0.8242188, 0.3187494, -0.3984375, 
    -0.3963547, -0.9481764, -1.184635, -0.8841152, -0.5671883, -0.6809883, 
    -0.1505213, 0.2713547, -0.2997379, -0.4674473, -0.4971352, -0.2950516, 
    -0.4229164, -0.1421871, -0.4067707, -0.5531254, -0.6960945, -0.2638035, 
    -0.5489578, -0.8192701, -0.5002613, -1.318229, -1.286719, -0.07083321, 
    0.2940102, -0.7830734, -0.6148443, -0.2859383, 0.2562504, 0.6841145, 
    0.6307297, -0.2104149, -1.018229, -0.9338551, 0.04739571, -0.04088402, 
    -0.7669268, -0.8445311, -0.3710938, -0.03333473, -0.04166698, -0.2601566, 
    0.1908855, 0.2174492, 0.1794271, -0.901041, -0.9604168, 0.04817581, 
    0.4197922, 0.1841145, 0.3981771, 0.2789068, -0.3289061, -0.8458328, 
    -0.08229065, -0.2492199, -0.8539066, -0.625, 0.1317711, -0.8791666,
  -0.421093, 0.6104164, -1.193228, -1.220314, 0.4716148, 0.5585938, 
    -0.3223972, -1.375, 0.1252594, 0.3322926, -0.5955734, -0.7044258, 
    0.2966156, -0.7309895, -1.358595, -0.4278641, 0.7367172, -0.5919266, 
    -1.982292, -0.7359371, -0.2911453, 0.07448006, 0.7815094, 1.584635, 
    0.5692711, -0.588541, -0.2635422, 0.1427078, -0.8476563, 0.05286407, 
    0.8867188, 1.021355, -0.3994789, -0.4640636, -0.01067734, -0.6023445, 
    -0.4192696, -0.6854172, -1.012239, -0.651041, -0.4963551, -0.6359367, 
    -0.7796879, -0.813282, 0.2242184, 0.478384, 0.2817707, -0.1291676, 
    0.2885418, 1.239063, 1.550261, 0.3388023, -0.01953125, 0.4666672, 
    0.8153648, 0.6065102, 0.9856777, 0.853384, 1.057032, 2.333593, 2.495834, 
    1.358854, 0.8023434, 0.8208332, 0.7432289, -0.2317715, 0.6171875, 
    0.4317722, -0.5091152, -1.576563, -0.4661465, 0.3867188, 0.6846352, 
    0.4039059, 0.4817715, -0.655468, -0.7510414, -0.5098953, -0.4166679, 
    -0.02942848, -0.2789059, -0.1690102, 1.250782, 1.513803, 0.3041649, 
    -0.1804695, -0.2632828, 0.6489582, -0.636198, -2.06875, -0.6973953, 
    -0.5471344, -0.5523434, -0.573698, -0.4429684, -0.5677071,
  -0.08775711, -0.1445313, -0.5135422, -0.8468742, 0.4179688, -0.3440132, 
    -0.2739563, 1.195313, 0.4565086, 1.352345, 0.8986969, 2.107552, 1.379948, 
    -0.5536461, -0.875782, 0.223175, -1.123436, -2.35651, -1.790367, 
    0.5979156, 1.919533, 0.1804695, -0.467186, -2.38073, -3.097916, 
    -0.9052086, 1, -0.1309891, -0.1583328, -0.06171799, -0.8255234, 
    -1.471615, -0.9927101, -0.691925, 0.5622406, -0.1164055, -0.3208351, 
    -1.050262, -0.9781265, 0.9244766, 0.470314, -0.5973969, -1.044792, 
    -1.29948, -2.531773, -1.150784, -1.141144, -1.444271, -1.037498, 
    1.243488, 3.284374, 1.633595, 2.552868, 3.943226, 2.666405, 0.903904, 
    0.7114563, 0.1341133, 2.877342, 4.03828, 1.841148, 0.1471329, 2.117451, 
    3.311455, 1.383854, 0.8958321, 0.7119789, 0.1161461, -0.2825546, 
    -0.9596367, -1.292709, -1.205471, -0.2388039, -0.1192703, -0.2841148, 
    -0.04426956, -0.1856766, 0.4906254, -1.430729, -0.6434898, 0.2546844, 
    0.1374969, -0.9507828, -0.188282, 1.191666, -1.250778, -1.991146, 
    -0.9981766, -0.3825531, -0.2544289, 1.214844, -0.2317734, -0.04114914, 
    0.598175, 0.5786476, -1.246876,
  2.949478, 1.349476, -1.718227, -1.779949, -1.844273, -1.62318, 0.003383636, 
    0.2473946, -0.8315125, -0.04869461, 0.09140778, 0.6291656, 0.1713524, 
    0.4578094, 1.390366, 1.159893, 1.204945, 0.09192657, -0.0695343, 
    2.352085, 2.290886, 1.912498, 0.8679695, 1.332813, -0.004428864, 
    1.096096, 1.846092, 0.591404, 0.05182266, -0.9281235, -1.048698, 
    0.7333336, 0.5859375, -2.045311, 1.038544, 3.565628, 2.152344, 1.772655, 
    3.342968, 2.950001, 3.650261, 2.673439, 1.127605, 2.750263, 2.261196, 
    0.7619781, 0.3966141, 2.788803, 1.361198, 2.619274, 2.465885, 2.625519, 
    2.78672, 2.608856, 1.125519, 2.316929, 3.018753, 2.498699, 2.336456, 
    4.209896, 5.152081, 1.017189, 0.9505196, 1.197918, -0.2598991, 2.580208, 
    0.996357, -0.4080734, 0.3932266, -0.4742203, 0.4481773, -0.4395828, 
    0.3330727, 0.96875, 0.9757805, -1.834896, -1.943489, -0.5942688, 
    -2.373177, -1.793755, 0.405468, -0.7304688, -0.688282, -0.1744804, 
    0.8854141, -0.954689, -2.20026, -0.9080696, 0.8367195, 2.0513, 0.7989578, 
    0.2106781, 1.693489, 2.484894, 1.324738, 1.800522,
  1.760414, -1.109898, -0.7122383, 1.303909, -0.05181885, 0.1825562, 
    1.145309, 0.8651047, 0.7596359, 4.738022, 4.217705, 1.288803, 1.088799, 
    2.649475, 1.717453, 1.890099, 0.9611969, -0.3489532, -0.6682358, 2.2901, 
    1.398697, 0.2989578, 1.843483, 3.720573, 4.769527, 4.292709, 1.374222, 
    1.386978, 0.6356735, 1.201828, 0.3429718, -1.426308, -1.828384, 
    -0.2156219, 3.067711, 3.595573, 2.115891, 2.981773, 3.430466, 1.926559, 
    1.829948, 3.272652, 1.550522, 2.155464, 4.898438, 4.127602, 2.254948, 
    4.374733, 4.010422, 1.546093, 3.074219, 4.003647, 4.091412, 3.096355, 
    3.586716, 2.066406, 1.939846, 1.450779, 2.186977, 2.158333, 3.929691, 
    1.472656, 1.708073, 4.340626, 3.448433, 2.802864, 0.8010406, 2.142708, 
    3.278385, 0.7317734, 0.4002609, 1.042183, 0.751564, 2.270054, 2.038536, 
    1.497398, 5.04948, 2.304688, 1.249481, -0.001304626, -1.620834, 
    -1.422401, 2.127602, 2.358856, 1.671349, -0.2833328, 0.3411484, 
    0.5661469, -1.704948, -0.4447937, 0.3023453, -0.3294296, 0.5223961, 
    1.18985, 1.390881, 2.29974,
  -1.48333, 2.128128, 4.017448, 2.762497, 1.704422, 2.848961, 2.360939, 
    1.794792, -0.5346375, -1.776825, 0.799736, 4.977608, 3.572136, 3.622131, 
    0.7364578, 0.5979156, 2.606247, 2.162239, 3.153122, 5.372398, 4.975006, 
    4.411461, 4.718231, 1.938805, 1.761719, 1.704948, -0.8502579, 2.414322, 
    2.50573, 2.933853, 1.504425, 2.486198, 3.449738, 4.489578, 5.014839, 
    4.400002, 4.307808, 5.590103, 7.426826, 9.953903, 4.882294, 1.278908, 
    -0.02942657, 3.417191, 2.757294, 1.616669, 3.323441, 2.549217, 3.313019, 
    2.225784, 6.452087, 6.784897, 3.613281, 0.7356796, 3.947136, 2.819534, 
    2.784637, 5.635162, 4.005203, 3.577606, 2.627602, 3.85807, 3.304947, 
    2.407288, -0.2872467, -1.604431, -0.1523438, 0.6036453, 1.544792, -0.875, 
    1.508072, 1.080467, 3.613281, 2.182816, 2.060417, 3.021355, 11.08021, 
    9.437241, 4.455727, -2.254433, -4.871613, -4.386978, -1.312233, -0.9888, 
    0.7916718, 0.9645844, 2.168488, -0.2408905, -2.078644, -3.088799, 
    -1.831772, -0.1828156, 0.2265625, 1.630989, 1.4375, 0.06562805,
  1.835411, 3.047394, 3.047394, 2.453125, 6.498695, 5.921616, 4.003647, 
    3.682808, 3.952347, 6.237762, 8.171875, 8.851044, 8.184631, 4.110153, 
    3.040627, 1.137245, 0.2450562, 1.258072, 1.783073, 3.264847, 1.60807, 
    2.341148, -0.2789001, -0.0687561, -0.6539078, -0.3997421, -0.2281265, 
    2.022911, 2.986458, 4.146088, 6.04583, 8.813019, 8.727341, 4.722656, 
    3.351563, 4.333076, 6.153381, 4.959892, 4.357811, 2.59687, -3.625519, 
    -3.833336, -3.169533, 0.3864594, -0.1013031, 2.31041, 2.169273, 4.058067, 
    4.808067, 5.425003, 2.122398, 3.142967, 0.3937531, -0.9742203, -0.266922, 
    -1.018227, 1.3526, 2.066925, 0.1075592, 0.748703, 0.685936, 1.512764, 
    1.691925, -2.314583, -6.188805, -0.2744751, -1.881508, -1.861458, 
    0.2450562, -1.301041, -1.74427, 0.1153641, 3.805473, 3.383858, 
    -0.9255219, 2.982033, 8.453384, 10.48099, 3.113281, -7.458855, -8.592972, 
    -5.020576, -4.436722, -4.854164, -0.8549423, 0.1708298, -0.9578094, 
    -1.460152, 1.664841, 0.8195267, -1.487236, -1.822395, -0.9072876, 
    -0.7536469, 1.416672, 0.0229187,
  1.862495, 1.091408, 2.704948, 7.092972, 5.09584, 5.655731, 8.594788, 
    6.237495, 5.013275, 4.7052, 6.280991, 2.30468, 3.335419, 3.112762, 
    0.8408813, 1.835159, -3.088806, 0.1325531, -3.341148, -2.553383, 
    0.5742188, -3.019531, -5.044792, 0.7606735, 0.4197922, 2.013023, 
    0.7156296, 0.2093735, 1.829948, 3.323959, 11.79037, 12.52161, 6.847656, 
    5.430206, 2.901306, 3.663544, 9.435417, 2.653381, -4.991402, -10.80964, 
    -13.99583, -11.69635, -0.5523453, -2.151817, -0.5112, 2.946358, 4.595055, 
    3.71302, -0.217453, 0.09036255, -4.166405, -3.175522, -1.432549, 
    -0.6846313, -2.401299, -0.0776062, -2.374481, -2.765106, -2.800522, 
    -2.778908, -3.14193, -1.870056, -2.379433, -2.540627, -2.536713, 
    0.5437546, 0.01979065, -0.8888016, -3.941406, -3.810677, -3.026566, 
    -1.914063, -0.1416702, 0.2393265, 0.110672, 0.4828033, 4.202866, 
    5.043488, -0.8864594, -7.837502, -11.36328, -1.828384, -4.523178, 
    -3.650261, -1.181252, -1.277863, -1.435417, -4.377602, -3.450783, 
    -4.00573, -2.677605, -1.182556, -2.184372, 1.353127, 2.778641, 2.171875,
  -2.331772, -1.359634, 2.141144, 1.439575, 1.282028, 6.373444, 12.03775, 
    6.702606, 1.936455, 2.712234, 2.841675, 3.596619, 4.03125, 3.175003, 
    4.316147, 2.888794, 2.993484, 0.09817505, 4.906769, -0.237236, 
    -0.3299484, -1.360153, -1.947655, -2.623436, -3.827347, -2.278648, 
    1.490891, -0.2940063, -0.6109314, 4.265625, 4.582031, 2.373169, 
    -3.770828, -2.101036, 0.606781, 1.097397, -6.47995, -11.80157, -11.95338, 
    -11.32396, -14.52708, -8.215881, 0.21875, -0.4320221, 2.010162, 3.438271, 
    0.3643188, 1.176308, -0.4773483, -4.121361, -2.155991, 1.012245, 
    -1.95755, 0.9304657, 0.1015625, 1.429688, -0.6572952, -2.627083, 
    -3.480209, -2.799217, -1.601303, -2.785416, -5.17057, -4.320572, 
    -3.648956, -4.085144, -2.157288, -3.519791, -3.056244, -4.738274, 
    -5.552078, -1.591667, 1.21666, 0.359375, -2.788544, -2.694794, -3.175247, 
    -1.415634, -5.441666, -10.79428, -9.179688, 3.063805, -1.179688, 
    -1.504944, 0.4424438, 3.073441, 2.890106, -0.7281189, 2.124222, 
    -0.7848969, -2.243484, 0.7273407, 2.109634, 4.5914, 3.019531, 2.452087,
  -1.909119, -0.2395782, -0.875, -0.2773438, -0.9260406, 6.780457, 8.472916, 
    3.210678, 2.188293, 0.505722, 2.1362, 1.436188, -0.6742096, -1.834641, 
    4.872925, 1.941147, 2.097137, 2.419006, 5.651031, 1.492188, 2.305206, 
    0.004684448, -0.1541748, -2.433853, -1.350784, 6.157303, 2.378113, 
    3.466415, 1.103394, 7.352081, 0.9078217, -3.740112, -9.973434, -7.771347, 
    -14.7211, -15.51405, -17.19244, -15.81094, -13.60495, -14.5401, 
    -8.641663, -1.253387, -2.11145, -4.22525, -2.203125, -3.145844, 
    -1.565628, -2.819, -0.3757782, 0.6385498, 1.303116, 2.243759, 1.432816, 
    3.367188, 3.5448, -0.9848938, -1.1539, -0.3489532, 2.440887, 0.7322998, 
    -2.860153, -5.106247, -4.24791, -4.376831, -2.028381, -0.6408844, 
    -1.546616, -2.529694, -4.376053, -3.410675, -0.8382721, 0.6031189, 
    -0.2093811, -2.545837, -2.950775, -4.744003, -3.652344, -2.648956, 
    -6.732025, -10.97578, 2.168747, 9.519791, 4.010147, 12.19036, 10.8362, 
    5.7677, 3.344025, 3.8237, 4.057816, -0.6062469, -0.1755219, 1.68515, 
    -0.3656311, -0.407547, -4.272919, -1.746094,
  -0.9166565, 1.714844, -0.7945404, -1.118484, 0.2226563, 5.836197, 2.232025, 
    2.906769, 3.800522, -1.510681, 2.806519, 4.890106, -2.526825, 2.199478, 
    -0.7960968, 2.969009, 8.535156, 4.563019, 7.484116, 6.275253, 2.990631, 
    -0.46875, 2.845047, 0.1994934, 0.1304779, 5.930725, 5.018738, 6.332809, 
    4.111465, 6.7211, -2.575531, -8.722137, -9.280472, -13.29713, -12.55417, 
    -10.45105, -11.49454, -8.86615, -10.98723, -5.572647, -0.494278, 
    -0.1468811, -0.3609314, -0.8614502, 1.969009, 4.050003, -2.679169, 
    -3.541931, -2.947403, 0.2937469, -3.668503, -4.525269, -1.216934, 
    -2.325256, -5.591415, -2.733856, 0.05703735, 0.8953094, -1.891922, 
    -0.7463531, -4.125, -3.202087, -2.281769, -2.924744, -4.807037, -2.75885, 
    -1.766403, -4.583603, -2.759109, 0.3377533, 3.195572, 2.187241, 2.623962, 
    4.552872, -1.155212, -10.75781, -3.264587, -3.769272, -8.478119, 
    -5.237762, 7.748444, 9.728134, 2.626816, 6.082031, 15.20911, 13.81067, 
    3.691147, 2.329956, -1.640106, 0.2945404, -2.654434, 0.8203125, 
    -2.184631, -0.7942657, -0.953125, 1.72345,
  0.505722, 7.408325, 0.6065063, -2.581772, 2.52916, 10.18828, 0.7218781, 
    2.768234, 4.918747, 3.634888, 5.249222, -2.296875, -4.452347, 0.8635406, 
    -3.543228, -2.402084, -4.850784, -3.255478, -0.6851654, -2.331253, 
    -3.154678, 1.623962, 3.83725, 0.161972, -2.45079, 0.8541718, 1.679688, 
    -1.185684, -2.091934, 1.593491, -0.2541656, -4.482559, -8.141144, 
    -8.741928, -6.98671, -4.863281, -1.630722, -5.680725, -3.027863, 
    3.890366, 3.387238, -1.672394, -0.532547, 1.769791, -0.2963562, 
    -5.022659, -5.125778, -1.069016, -0.8479156, -4.18515, -1.989578, 
    -0.1374969, 1.854416, -0.1091156, 6.132034, 5.538803, 3.671616, 2.924988, 
    3.960938, 3.897125, 1.11145, -1.034119, -1.7724, -1.232819, 1.662231, 
    3.344269, 4.578903, 2.955215, 4.480728, 5.051559, 5.369019, 8.884888, 
    4.744797, 7.05365, -0.4609375, -0.7536469, -0.5674438, -2.706512, 
    -8.186195, 8.760422, 7.213287, 5.57135, 3.170563, 1.862503, 18.75104, 
    16.51901, -3.350784, -0.1760406, -0.2434845, -1.245575, -2.345581, 
    1.93959, -2.612503, 1.095322, 0.1239471, -0.7747345,
  0.8098907, 1.850266, -6.072906, -1.730469, 1.897659, 10.31458, 1.128113, 
    7.691147, 12.11223, 10.69635, 14.30833, 2.678909, -4.968491, -3.191406, 
    -2.963791, -6.812241, -7.887497, -3.644272, -9.213013, -10.80756, 
    -6.547653, -8.029694, -7.847656, -6.940628, -2.745056, -1.0065, 1.314575, 
    -1.542191, -2.934113, -1.514069, 2.796097, 3.702072, -3.708344, 
    -5.626312, -6.798706, -8.525772, -2.123703, -4.201828, -0.5861969, 
    5.819275, -1.0849, -1.500793, -0.4114532, -0.1151123, -5.071091, 
    -6.97995, -4.135422, -2.954697, 1.478394, 4.784897, 1.962494, -0.8940125, 
    -0.7216187, -2.084641, 2.040878, 4.748688, 6.183075, 4.694016, 5.873169, 
    1.098175, -0.2065125, -0.5513, -0.8377533, 2.491928, 0.5562439, 2.883072, 
    5.015366, 2.998962, 4.141663, 8.494537, 9.546356, 11.52423, 11.06406, 
    10.34634, -2.528122, -4.677612, 8.639053, -0.4390717, 3.670837, 9.31041, 
    7.161728, 6.02005, 9.018753, 3.000778, 13.17813, 13.79011, 3.991928, 
    -1.720047, -0.9458313, 2.348694, -1.078644, 1.899994, -2.604172, 
    2.763275, 2.290359, 4.821091,
  5.585419, -0.3723907, -4.117188, -4.099731, -5.318497, -5.717712, 
    -6.298431, -6.564331, 5.827087, 6.532028, 13.10364, 5.918762, 3.772141, 
    5.157043, -0.3010406, -0.1187592, -3.279419, -1.859375, -8.399475, 
    -8.630463, -12.02605, -15.69505, -10.63803, -9.339325, -1.994797, 
    -1.714066, 0.1692657, -2.135681, -0.1135406, -0.8856812, -1.311966, 
    1.412766, -1.130981, -0.03672791, -2.635147, -3.708328, -4.1474, 
    -6.383331, -8.772141, -0.8770905, -4.153137, -2.433075, -3.108597, 
    -4.925003, -7.780212, -8.876053, -5.853653, -2.740875, 1.485687, 
    4.743744, 2.682541, -1.647919, -5.226563, -3.9599, -0.9583282, 4.149216, 
    5.259384, 4.410416, 2.734894, 2.097137, -0.0302124, 1.480209, 0.5434875, 
    2.191147, 0.3763123, -0.7585907, 0.8341217, 3.407806, 6.268234, 9.617966, 
    9.563797, 10.62604, 11.58438, 5.931259, -1.736206, 1.345322, 12.63594, 
    11.60912, 4.923431, 7.436981, 7.615631, 7.378387, 7.389069, 5.548431, 
    12.03671, 12.66692, 15.72318, -3.086975, -0.6799469, -0.9559937, 
    0.3187561, -8.831253, -1.253906, 0.8752594, -0.005996704, 2.474472,
  -0.5205688, -0.1010437, -2.777344, -2.385147, 0.6817627, -7.245575, 
    -8.802597, -16.68437, -13.74843, 9.944275, 21.46172, 14.19453, 4.918488, 
    9.739578, 9.503387, 5.402603, 8.633591, 6.316925, 1.020844, -4.265625, 
    -7.058594, -5.54245, -6.189835, -0.4684906, 3.021866, 4.099731, 1.396866, 
    -4.080734, 3.68074, 1.552078, 1.186203, 2.403656, 0.8687592, -2.552856, 
    -2.085678, -1.298172, -1.251038, -2.733597, -7.058067, -15.13385, 
    -14.44376, -13.05182, -6.339325, -2.551559, -10.94948, -8.700775, 
    -1.581253, -1.447906, -3.449738, -2.59375, -3.104156, 0.3190002, 
    0.9705658, 2.358597, 2.541672, 3.264847, 1.940109, 2.159637, 2.890106, 
    6.236969, 8.217194, 6.739059, 5.22345, 4.48645, 0.8408966, 1.031769, 
    0.84375, 2.383606, 3.265106, 4.287491, 4.139313, -0.4414063, 0.5966034, 
    1.12265, -2.880737, -3.510422, -2.34375, -0.0249939, 5.664841, 7.18985, 
    6.578644, 14.48386, 13.53386, 4.172913, 5.569794, 5.816925, 7.473969, 
    4.330994, 2.325531, 2.7836, 1.371094, -4.874481, -1.339584, 0.3864594, 
    -1.332031, 1.122131,
  4.748169, 2.399216, 2.579681, 10.49376, 5.63385, -10.39322, -4.829681, 
    -17.48749, -14.47136, -13.1013, 3.159897, 16.93906, 10.89792, 1.072922, 
    1.309906, 2.520065, 1.888016, 0.6364594, -1.157562, -2.849472, 
    -0.6612091, -4.608856, -6.966919, -4.036713, -0.6395874, 2.59375, 
    -0.5320129, 1.646881, -6.876297, -5.063293, -0.3669281, 4.418747, 
    8.422134, -0.8541565, -1.4487, 1.520569, 4.855728, 3.587769, -9.840622, 
    -14.9547, -7.554688, -1.668747, 2.746872, 10.04478, 5.096085, 1.815628, 
    8.495834, 6.332809, 0.1648407, 0.02110291, -4.735428, -4.450531, 
    -3.25209, -4.412247, -7.204163, -6.877869, -7.302338, -6.581512, 
    -8.682816, -7.359634, -6.49765, -5.167969, -2.564056, -4.266418, -3.1763, 
    -2.191406, -3.703384, -3.633347, -3.600266, -1.412247, -1.535675, 
    -5.269272, -10.91145, -8.719009, -3.391678, -2.011993, 10.15546, 12.8065, 
    -0.4367218, -0.453125, 3.728134, 17.86589, 26.10573, 12.94583, 11.98308, 
    11.26068, 4.916931, 4.408859, -0.4739532, 6.193481, 6.411987, 2.82579, 
    2.788528, 0.7156219, 1.546356, 2.975525,
  -1.782547, 0.07395935, 5.682281, 18.47551, 12.85495, 3.725784, 5.896088, 
    -0.6229248, -0.9286499, -21.15756, -9.416412, 6.405487, 14.75208, 
    -0.6580811, -3.433075, 0.7111816, -0.5513, -1.166382, 2.2742, 1.913788, 
    -1.958069, -7.628906, -6.396088, -6.590363, -5.291931, -3.286438, 
    -6.340363, -2.930466, -5.965103, -5.0159, -9.488022, -5.621872, 
    -4.348175, -8.170303, -5.617706, -8.96666, -6.970566, -8.134384, 
    -4.446091, 7.724747, 9.795563, 9.329956, 4.470322, 6.051575, 8.660675, 
    10.45103, 9.221619, 0.5570374, 2.291672, 3.021362, 2.501556, -1.363541, 
    -1.328644, -1.29715, -3.796631, -5.370056, -6.198456, -8.665894, 
    -10.40704, -7.832581, -10.29404, -10.12473, -9.115356, -8.194275, 
    -5.178375, -4.380737, -4.411713, -6.425262, -6.00235, -6.9664, -12.90417, 
    -20.40025, -26.32838, -19.33333, -14.27605, 9.695313, 9.679413, 4.3797, 
    6.888031, -0.6372528, -7.238022, 1.59819, 17.49219, 11.53777, 14.84608, 
    11.70183, 8.093491, -0.5799561, -6.438553, 2.034363, -1.008331, 1.807281, 
    -2.760925, -4.347397, -3.095566, -1.683075,
  9.251572, 3.63385, 5.896622, 10.03255, 14.59766, 0.3679657, 1.109116, 
    17.6427, 13.10599, -9.289581, -9.538803, 0.9997406, 15.69453, -0.177887, 
    -2.979431, -0.2460938, 2.7435, -1.293488, -2.209381, -3.754181, 
    -2.858063, -8.446594, -7.767426, -7.570068, -4.860687, -4.659119, 
    -7.503906, -17.92004, 0.4140625, 2.046356, -6.7388, -6.045059, -3.675003, 
    -0.9885406, 0.335144, -5.817978, -4.338287, -3.72995, 5.394791, 4.092438, 
    3.116669, -0.8265533, -5.252594, -5.365372, -0.02812195, 4.167969, 
    -0.1085968, -0.1763, 0.6171875, 2.797653, 4.401047, 3.470322, 3.672394, 
    3.60965, 0.6153717, 4.776306, 2.583862, 1.045319, 1.0914, 0.3414001, 
    -2.685669, -0.5445251, -1.378662, 0.7440186, -0.0791626, -1.331512, 
    -0.05337524, 1.879944, -0.8046875, -6.859894, -10.17786, -15.20677, 
    -15.65027, -14.13776, -8.847916, 13.8427, 5.639328, 6.418488, 17.78307, 
    5.747925, -1.6698, 0.414856, 2.1138, -0.1171875, 6.300507, 6.302353, 
    6.952576, 2.364319, 4.24765, 6.265106, -0.0947876, 1.398193, -1.666412, 
    -1.136719, 7.978119, 7.892197,
  8.345062, 15.57448, 7.986725, 8.338287, 3.935425, 1.600525, -1.386978, 
    5.994003, 6.803635, 14.46251, 32.48567, 2.305725, 3.732574, -1.410675, 
    -3.920074, -1.560425, -0.2887878, 0.01483154, -1.240082, 2.706757, 
    -3.275269, -17.5289, -15.32864, -9.469788, -7.1427, -0.1625061, 
    -6.777863, -13.32709, -6.963806, -3.826553, -0.6075745, 0.2958221, 
    -0.1177063, 0.15625, -9.869263, -8.425522, -6.597656, -7.826035, 
    -6.661453, -9.0896, -10.35834, -6.931778, -11.25728, -10.52216, 
    -5.986725, -2.596893, -5.589844, -4.911987, -1.356781, -5.145844, 
    -5.982025, -9.262238, -7.039581, -6.119537, -3.656006, -6.07135, 
    -3.130188, -1.408325, -0.9786377, -0.3815002, 5.077087, 6.595825, 
    6.547394, 5.191162, 3.539581, 4.636993, -0.4333496, -0.870575, -6.0336, 
    -9.572388, -11.31561, -7.973175, -8.467972, -7.304428, 10.68021, 28.625, 
    19.89011, 22.08047, 5.847656, -7.327362, -10.25156, -12.37735, -9.135666, 
    -4.648972, -1.485931, 0.7059937, -0.7432404, 0.129425, 1.314301, 
    -3.139069, -2.1474, -10.93542, -3.098175, 10.14818, 9.284103, 17.92735,
  -2.837219, -1.019012, -2.8125, -0.1177063, -1.775787, 4.614319, 7.121613, 
    5.931488, 8.657532, 20.3909, 10.60599, -1.818237, -0.5320435, -2.419281, 
    -3.933594, -1.408875, -3.011475, 1.285675, 1.510956, 0.2583313, 
    -8.802338, -20.79999, -18.01587, -17.58127, -13.05548, -1.204956, 
    6.477875, -4.998688, -20.95599, -7.739319, -1.248199, 0.1023254, 
    -3.446106, 2.153915, -8.869781, -5.867706, -10.40025, -11.3474, 
    -8.694519, -12.38019, -10.78384, -6.033356, -7.671082, -7.30835, 
    -9.447906, -3.309631, -6.886963, -8.198425, -3.510162, -5.903381, 
    -5.957306, -1.858582, 0.5872498, 0.2453308, -4.46405, -1.940369, 
    1.982544, 3.350525, 0.966156, 4.504181, 6.80545, 9.889557, 13.11691, 
    11.54895, 14.45651, 15.30939, 8.548462, 3.812225, 0.7679443, -2.713013, 
    -5.969513, -8.678375, 0.8718719, -1.009384, -2.510147, 5.430466, 
    8.076294, 3.463043, -0.5661621, -14.58853, -12.93698, -8.409119, 
    -6.156509, -5.649475, -1.737762, -0.9510193, -1.514069, 2.572662, 
    -2.620331, -4.175507, -9.780731, -6.625519, -2.348694, 0.1145935, 
    -2.814056, -1.545837,
  -1.969788, -1.078918, 1.630707, 1.616913, -0.3997498, -1.776031, 0.2255249, 
    6.886444, 4.589294, 4.701538, 1.719543, -0.3771057, 7.245331, 1.632294, 
    -4.381744, -6.263306, -4.891418, -4.97525, 0.7953186, -9.936966, 
    -5.419525, -16.06226, -23.6987, -17.72238, -10.5513, -3.308075, 10.05389, 
    -6.314056, -16.47971, 0.2778625, 1.904144, 9.893494, 8.940094, 
    -0.1458435, 4.181519, -0.5223999, -4.934113, -6.867188, -6.335419, 
    -2.560425, 0.1343689, -3.376556, -2.987488, -5.836212, -3.697144, 
    -6.524231, -6.405457, -5.542969, -3.742188, -6.825775, -5.099243, 
    2.219513, 5.7164, 1.804962, 1.050781, -1.634888, -1.266937, 1.550781, 
    2.546356, 5.661728, 8.878143, 13.53438, 17.45703, 18.66565, 20.29688, 
    9.015625, 6.426025, 7.429688, 4.882294, 5.962738, 7.6763, 8.885422, 
    6.136185, -6.987244, -8.166931, -3.497894, -2.969543, -3.337219, 
    -3.301849, -8.667175, -8.179169, -10.74792, -9.40184, -5.0177, 
    -0.3249969, 0.7083435, -0.9450378, 1.847931, 0, -1.585144, -4.166687, 
    -5.991394, -1.600525, -3.02475, -4.176819, -4.997162,
  -1.654175, -1.929443, -0.2174377, 1.08075, 3.977631, 3.096863, 2.610931, 
    1.923706, 1.923157, 3.207031, 3.744537, 4.040619, 5.488007, 1.557037, 
    -0.617981, -4.708862, -7.21405, -8.970306, -3.458862, -6.177612, 
    -3.798706, -9.063019, -11.13724, -12.80704, 1.242706, 8.825241, 5.630219, 
    -14.28152, -12.09164, -5.029175, 2.6651, 1.577881, 4.457275, 9.132538, 
    11.78204, 6.029938, -1.678131, 1.028656, -4.1073, -1.255737, 1.300232, 
    -1.146362, -1.446106, -4.748444, -7.461456, -7.463806, -7.314056, 
    -6.968506, -12.41693, -9.913544, -7.369507, -7.087219, -4.856506, 
    -5.474731, -4.219025, -7.653656, -1.154419, 0.401825, -3.68515, 4.4375, 
    4.258591, 8.187256, 4.919037, 10.56171, -0.2567749, 2.682037, -4.07135, 
    -0.1596375, 7.317719, 18.77969, 10.08907, 8.770569, 5.761993, -6.8172, 
    -5.200256, -1.698456, -0.3768311, 0.06018066, -4.157043, -8.8992, 
    -10.95364, -7.612518, -9.358063, -3.967712, -6.449234, -2.513794, 
    0.2236938, 4.6492, 1.273712, -1.910675, -5.115356, -4.307526, -2.855713, 
    -1.335938, -3.364868, -2.153931,
  -4.082794, -3.251038, -5.952881, -4.549225, -3.564575, 0.7578125, 1.989319, 
    2.630981, 3.141907, 1.283325, 0.8312378, 4.456787, 6.702576, 4.186462, 
    4.559143, 1.3461, -1.092957, -1.865631, -3.084625, -4.250275, -4.371613, 
    -5.760437, -9.858063, -9.921875, -5.749237, -10.07059, 2.239594, 
    4.338806, -3.252869, 3.555984, 2.582031, 4.885941, 7.5625, 8.746094, 
    14.21484, 18.35677, 10.92969, 0.992981, -0.580719, 2.572662, -0.194519, 
    -2.078918, 0.3643188, -2.820557, -6.384888, -9.746613, -9.852875, 
    -9.218231, -9.343475, -8.292969, -9.747131, -4.621857, -12.83463, 
    -5.869263, -8.335938, -6.583344, -5.374237, 0.9526062, -2.732819, 
    -5.994781, -3.612488, 1.168243, -0.7221375, 1.590118, -2.6026, -2.188538, 
    -3.64975, -9.835144, 0.3145752, 9.470337, 2.007294, 2.017181, -1.729431, 
    -2.749725, -1.220825, -5.342468, -2.211975, -1.293213, 2.342712, 
    4.094543, -1.200012, -2.414063, -5.889069, -3.626312, -4.468994, 
    -5.095306, -4.686707, -0.4387817, 0.1395569, 5.099976, -2.634888, 
    -2.027069, -2.348175, -0.5242004, 0.01223755, -2.503906,
  -2.83075, -3.476318, -5.851288, -5.586975, -1.795319, 1.887512, 2.757294, 
    3.487244, 5.509644, 4.117462, 3.444519, 5.403656, 10.40784, 7.230743, 
    8.012238, 9.980743, 4.879944, 1.739594, 1.639587, -0.70755, -3.233856, 
    -3.936981, -8.458069, -7.951813, -11.4422, -5.524231, -8.951828, 
    1.753647, -0.4664001, -0.8914032, 2.719528, -2.1474, -1.221359, -1.96666, 
    6.471878, 7.672134, 5.421341, 4.598434, 4.345825, 0.946106, -5.759125, 
    -10.48203, -5.480988, -3.383087, -3.169281, -6.253662, -9.397919, 
    -12.37057, -8.940369, -7.095581, -1.809113, -1.58725, -4.288025, 
    -0.9960938, -6.249725, -9.010956, -7.145325, -8.816162, -4.223175, 
    -5.134399, -1.3862, 0.1898499, -1.30365, 0.6362, -4.814301, -1.161469, 
    -2.573181, -7.835175, -5.381775, 3.692719, 4.028625, -0.7794495, 
    -4.236969, -4.467712, 2.996094, 1.280731, 2.799469, 8.056519, 5.8125, 
    2.380707, -2.441406, 1.800018, 2.934387, 0.08853149, -1.963013, 
    -4.395294, -2.467957, -2.721893, -2.105743, 3.266907, 4.137756, 
    -3.150787, -0.6791687, -0.6075745, 1.157532, 0.9835815,
  1.698456, 0.5684814, -0.5789185, -4.497925, -1.487488, 2.479431, 2.554962, 
    4.674469, 1.789612, 4.326324, 7.939819, 7.167969, 4.145294, 6.98465, 
    15.40103, 14.76535, 12.95132, 10.03229, 13.83777, 4.935425, -1.930725, 
    2.715118, -21.10809, -7.393463, -6.730988, -8.434113, -12.68282, 
    -5.478119, -3.258072, 7.151566, 5.826813, -6.018494, -7.457031, 
    -8.994278, -7.277603, -6.293228, -5.147919, -2.701828, 0.8487091, 
    7.68959, 2.317459, -1.693222, -3.5802, -5.502335, -4.347931, -3.012756, 
    -3.646362, -0.9377441, -0.6700439, -2.381775, 0.9046936, -0.986969, 
    3.431763, 4.911194, -0.1546936, -1.331512, 0.2877808, -1.441162, -4.6185, 
    -1.469025, -3.019257, -1.954163, -1.8573, 0.3114624, 1.2612, -1.583344, 
    -1.239349, 1.208069, 1.214081, -1.638, -5.433594, -2.132813, -2.593506, 
    -2.340881, -2.270844, -1.263306, 2.857819, 9.73465, 5.612244, 7.221344, 
    10.45679, 5.240631, 2.164856, 3.646606, 0.9609375, -1.408325, -4.846893, 
    -0.1791687, -0.01797485, -0.841156, 2.612213, 1.546356, -4.3685, 
    -0.546875, 4.592194, 7.674744,
  14.98752, 11.33957, 7.686432, 2.344543, -5.943481, -4.238525, 0.7182312, 
    3.489349, 2.331268, 3.968231, 6.94455, 8.694794, 19.39063, 29.34586, 
    24.07968, 11.67343, 11.6698, 22.8013, 28.04895, 13.68256, -5.575287, 
    -29.15442, -25.33386, -24.43619, -40.86902, -18.49841, -5.593506, 
    -1.201813, -5.200256, -2.327866, 5.890625, -1.830978, -6.289581, 
    -6.483856, -8.366928, -9.636444, -5.437241, -1.008347, 1.978134, 
    3.020065, 6.278397, 10.80313, 6.949738, 0.8809967, -1.725266, -0.7182159, 
    -1.871094, -2.302322, 2.388535, 3.040634, 1.608093, 6.600281, 11.82578, 
    10.94659, 11.27472, 4.515106, 4.745575, 5.309631, 2.887238, 1.840118, 
    0.7346191, 4.270569, 1.857819, 4.431488, 4.833313, 4.463562, 5.932281, 
    12.08307, 12.21902, 8.116394, 2.0979, -3.132019, -0.004699707, 6.333344, 
    1.733856, -3.514862, -5.254669, 3.180481, 10.16196, 13.92969, 8.771881, 
    4.192169, 4.529419, 3.79425, 1.665375, 0.1281433, 0.111969, -3.384369, 
    -2.36615, -3.101837, -0.9541626, 3.77005, 4.214325, 4.000519, 16.08594, 
    21.88019,
  26.63124, 1.279938, -0.3161621, 2.632294, 0.1583557, 6.023193, 16.03671, 
    16.19218, 16.53749, 5.671616, 9.959381, 12.41014, 24.89661, 11.59637, 
    8.869293, 15.44141, 16.03543, 8.6362, 10.84949, 0.270813, -14.70132, 
    -6.295288, -5.951569, -10.93933, -16.97812, -13.59897, -15.45364, 
    -2.507538, -2.332581, -3.6474, -5.180969, -6.012787, -8.594818, 
    -1.936218, 0.7645874, -11.92343, -14.50156, -4.396881, 2.300781, -2.6026, 
    -3.671875, 1.261459, 3.034637, -0.6885376, 1.6763, 3.843231, 0.3945313, 
    1.714584, 3.049469, 5.305481, 3.791931, 5.926559, 3.856522, 3.44426, 
    6.048431, 7.49791, 4.599228, 9.268219, 7.681, 4.650787, 8.044525, 
    4.514587, 4.537231, 12.1539, 15.05676, 19.10312, 18.28464, 16.52344, 
    20.8927, 20.83279, 11.92941, 5.5961, -0.2921753, 3.288544, 6.185684, 
    8.110153, -1.215363, -1.787231, 1.055725, 0.7109375, 3.958344, 7.542969, 
    3.263016, -2.088806, -5.912506, -7.725021, -4.921112, -1.976563, 
    -0.3528748, -0.8208313, -0.1346436, 0.2401123, 6.590637, 17.84973, 
    24.40182, 30.27603,
  23.27136, 1.343231, 10.03177, 21.83855, 8.201538, 18.09843, 18.39037, 
    9.487762, 7.471878, 0.7531281, -0.2953033, 10.14375, 12.6862, 0.229187, 
    2.341431, 3.195313, 6.102081, 1.569519, 3.795319, 9.149231, 11.13699, 
    4.017944, -2.6474, -4.15625, -5.56665, -2.714325, -5.069794, -11.60522, 
    -6.916931, -1.078644, -3.046875, -7.092438, -3.982819, 1.609375, 
    8.879684, 0.4460907, -8.671631, -3.875, 6.211197, 0.5502625, -4.669525, 
    -3.432297, -4.79921, -11.68515, -10.44974, -4.517456, -2.469528, 
    -0.1343689, -0.7999878, -3.941925, -0.806778, 1.191925, 3.960159, 
    3.198959, 5.122131, 7.393738, 3.373962, 1.738281, 0.8583374, 4.78801, 
    5.349731, 1.879425, 2.771088, 8.279694, 5.458862, 9.217712, 9.856247, 
    9.58905, 14.29166, 14.38803, 13.86798, 4.797134, 2.913025, 1.199997, 
    -0.9276123, -1.180984, 0.6007843, -4.482803, -6.473694, -7.738556, 
    -11.42578, -8.678909, -2.934128, -2.401306, -5.047913, -11.29375, 
    -9.420837, -3.138809, -5.30365, -4.357819, 0.4635468, 4.067703, 4.293991, 
    9.623444, 26.08151, 44.57448,
  9.734634, 8.238815, 14.64818, 4.880219, 4.690369, 8.090103, 5.731766, 
    6.102081, 4.120056, 2.212234, -5.463791, 0.02993774, 3.302338, -3.213806, 
    -3.782288, -5.889862, -4.507019, -2.679169, -2.453369, -1.83075, 
    -3.885681, -3.030487, -7.251068, -8.893494, -10.58594, -8.696869, 
    -14.23438, -14.60886, -8.712524, -6.276581, -4.799225, -10.86798, 
    -6.967697, -7.574753, -10.73203, -6.123688, -2.19426, -0.71875, 
    -0.9992218, -4.896103, -6.775772, -6.606522, -1.706772, -0.8125, 
    -5.376297, -7.027603, -6.338531, -8.288284, -8.460159, -4.78125, 
    -3.461716, -2.420044, 3.158066, 2.946625, 2.847916, 5.221603, -2.052078, 
    -3.363022, -4.835938, -3.362244, -5.100006, -9.132813, -5.446884, 
    -1.823685, -1.9263, 0.9005127, -0.3578186, -0.6953125, 2.530731, 
    2.668747, -2.010681, -9.229172, -8.655731, -9.670303, -6.142715, 
    -9.646088, -10.48724, -12.13437, -9.755997, -4.948166, -7.237762, 
    -8.401031, -6.401291, -4.720306, -11.60416, -15.52577, -15.67578, 
    -12.2948, -10.73593, -10.82813, -5.847137, -2.501556, 0.4132843, 
    -4.987503, -2.06041, 15.34167,
  2.478394, 2.954681, 1.158066, -0.3153687, 2.333588, 2.731766, -1.493744, 
    -0.4203186, 3.882813, 4.260422, -2.302856, -7.252594, -7.375519, 
    -10.91223, -12.53488, -12.31537, -11.31979, -8.522919, -5.852615, 
    -3.552887, -5.711212, -5.404419, -10.21223, -15.52031, -13.97083, 
    -14.63046, -16.07266, -14.30391, -8.129166, -8.309891, -8.032562, 
    -9.647659, -5.406509, -4.994537, -8.300003, -3.732285, -0.4908905, 
    -2.335419, -11.23201, -3.722656, -0.5364685, -2.315109, -6.315628, 
    -9.758331, -7.170059, -3.813278, -7.840103, -11.56511, -9.478897, 
    -5.890625, -1.304169, -1.421341, -0.8867188, -1.006241, 3.916672, 
    6.359894, 4.263016, -3.273697, -5.606262, -8.72995, -10.50598, -6.188553, 
    -11.94061, -17.32709, -20.84505, -12.32317, -11.96666, -13.74193, 
    -17.34532, -10.29141, -8.149216, -7.587234, -10.59427, -14.24089, 
    -11.19531, -16.06537, -16.37813, -15.12709, -10.81483, -9.568237, 
    -8.222916, -13.10989, -8.503387, -1.305206, -5.549728, -9.822922, 
    -12.77266, -20.92604, -15.88568, -11.86145, -10.89844, -4.835159, 
    -1.113281, -4.522125, -2.209366, 5.608856,
  -0.9013062, -3.605209, 0.5429688, 3.982025, 6.670837, 6.650253, -0.7414093, 
    -3.956253, -3.640884, -2.806519, -10.98489, -15.8638, -10.55598, 
    -13.14713, -14.48412, -17.07265, -14.40677, -18.72658, -19.96718, 
    -19.23515, -14.89088, -11.97762, -16.71562, -14.25078, -10.81172, 
    -4.885422, -3.542969, -7.920044, -8.552612, -7.808594, -12.5211, 
    -13.66797, -9.505203, -8.074478, -7.704941, -3.575256, -2.086975, 
    -6.561981, -19.42551, -2.420837, 0.9828033, -7.716934, -21.62109, 
    -21.41875, -16.66901, -10.07864, -6.292709, -4.355209, -4.1138, 
    -4.961197, -6.024994, -4.582809, -1.454163, 2.114838, 5.208328, 5.820847, 
    1.261459, -2.811722, -5.003128, -7.885925, -12.93881, -16.94037, 
    -27.81718, -23.494, -16.58542, -18.53647, -19.98671, -14.93855, 
    -11.55859, -8.588791, -10.92865, -17.95233, -15.49739, -13.66536, 
    -14.53802, -33.02734, -12.70703, -13.07942, -9.37735, -12.60078, 
    -12.99324, -31.23697, -9.444794, -3.141144, -4.664322, -5.416412, 
    -6.441406, -5.407303, -3.24765, -3.376297, -7.824493, -9.957809, 
    -6.532303, -5.730469, -2.401047, -0.1143188,
  -17.70078, -19.67058, -16.34323, -5.918488, 2.751556, 3.436447, -5.483841, 
    -12.75417, -21.28203, -16.18933, -11.55547, -16.47916, -17.76796, 
    -18.90912, -22.869, -31.15051, -29.26302, -16.07996, -17.00626, 
    -21.49896, -21.2948, -20.04584, -13.34975, -11.77553, -17.97369, 
    -16.76068, -7.365875, -6.44635, -11.25078, -16.18985, -13.59349, 
    -17.35052, -9.176819, -5.561462, -0.5072937, -0.6791687, -4.021606, 
    -5.284637, -21.03101, -5.593491, -5.199493, -8.170563, -17.94376, 
    -23.21094, -17.00963, -11.47343, -6.613281, -2.295059, -2.456253, 
    -2.205734, -0.2463531, -0.4109497, -1.813293, -4.311722, -11.43932, 
    -10.04713, -10.23463, -8.211731, -6.697144, -10.24011, -21.17371, 
    -38.59634, -26.55598, -10.63905, -11.00157, -15.45155, -18.17395, 
    -11.73489, -10.10468, -6.452591, -16.23567, -24.70078, -33.72681, 
    -30.35367, -25.66821, -24.70392, -17.94427, -20.83801, -14.76927, 
    -14.36354, -24.78619, -26.64272, 0.7234344, 4.783066, 3.246368, 3.319534, 
    0.4367218, -6.273178, -6.834122, -5.854431, -4.564835, -3.618225, 
    -1.201294, -0.7013092, -2.865372, -6.277603,
  -7.631516, -9.823959, -9.561188, -13.33879, -5.986969, 0.1679688, 
    -1.666931, -6.980469, -15.39142, -18.99245, -14.94922, -16.17604, -17.5, 
    -15.88698, -19.69505, -20.19922, -18.61356, -17.62735, -18.51172, 
    -23.39063, -24.08749, -21.19583, -17.31119, -11.74791, -11.21719, 
    -14.7099, -16.16953, -12.34245, -9.074997, -11.18411, -18.1138, 
    -18.65547, -19.0948, -16.5901, -7.190094, 1.339325, 5.284637, 8.180725, 
    5.78569, -0.8286438, -1.633331, -5.058853, -10.27605, -16.86771, 
    -18.63281, -21.50157, -20.53621, -39.0461, -14.35808, -11.06433, 
    -14.08385, -20.71458, -15.53647, -19.21901, -22.91927, -31.27083, 
    -33.51692, -27.06641, -25.64531, -20.39246, -17.49713, -14.78542, 
    -9.018234, -2.672394, -4.226303, -12.08125, -16.1987, -15.86954, 
    -20.4362, -21.55365, -22.04713, -26.25415, -24.10391, -12.98721, 
    -11.24609, -19.7565, -21.94376, -19.09479, -20.48645, -16.00027, 
    -18.13593, -18.70209, -4.175262, 5.733063, 5.184113, 7.106247, 5.165634, 
    3.317459, 4.479691, 3.797134, 1.747925, -3.201294, -10.15494, -10.55624, 
    -12.50546, -8.841934,
  -9.836456, -10.83803, -6.769012, -6.373688, -7.321625, -5.754166, 
    -7.367966, -11.5159, -12.1776, -16.11041, -12.37396, -10.92708, 
    -12.14818, -17.32213, -18.3409, -18.24271, -17.88177, -15.35182, 
    -12.49974, -10.82579, -14.26042, -18.39011, -17.84738, -10.44402, 
    -6.981506, -7.738541, -4.636719, -8.694275, -13.36693, -11.25104, 
    -13.03438, -12.54974, -11.05026, -6.857544, -0.4580688, 2.153122, 
    5.28125, 9.648956, 7.799225, 3.499466, -5.124741, -8.391663, -8.082809, 
    -11.00182, -10.87057, -11.40079, -12.29897, -13.66147, -14.47708, 
    -10.38802, -12.44141, -22.89948, -16.60782, -12.3513, -11.90964, 
    -11.04062, -8.052078, -7.960678, -10.71875, -12.14375, -9.049484, 
    -7.596085, -4.625519, -6.276047, -12.21146, -17.92267, -22.09843, 
    -22.52605, -21.65051, -22.90392, -21.91145, -20.00572, -14.08047, 
    -6.733078, -8.600525, -12.52917, -16.05, -18.1862, -21.51042, -19.86328, 
    -18.1013, -18.21979, -10.60834, -6.518234, -3.719269, -2.155991, 
    1.478394, 2.574997, -3.7052, -3.990891, -3.172394, -6.126831, -1.4375, 
    -3.978134, -4.905991, -6.642975,
  -5.532547, -3.187759, -0.433075, -0.2890625, -2.079422, -4.597656, 
    -9.578384, -7.988281, -2.871353, -0.3486938, -2.642441, -13.46745, 
    -13.00131, -15.43985, -7.112503, -13.55026, -19.48828, -20.00572, 
    -17.85078, -12.83958, -7.064835, -5.787247, -7.490356, -10.80754, 
    -13.01563, -6.666931, 0.8726654, -0.6132813, -1.208588, -2.925522, 
    -5.749741, -3.755478, -3.755722, 2.897385, 5.525787, 1.936462, 2.122131, 
    -1.577866, 1.069794, 3.039581, 5.618225, 5.635422, 3.216141, 2.682556, 
    -1.180466, -4.582291, -4.061981, -5.510162, -5.857025, -7.492706, 
    -11.58488, -17.10938, -21.14738, -13.47318, -12.06978, -13.0789, 
    -13.21667, -11.86719, -14.42317, -13.80104, -15.56796, -16.86224, 
    -17.1823, -17.19037, -20.22136, -21.6888, -25.29558, -21.60991, 
    -15.81744, -13.21588, -11.88907, -12.14973, -6.082291, -4.336212, 
    -8.350266, -13.50702, -15.74141, -20.02655, -18.08203, -12.57082, 
    -8.369263, -6.568726, -2.5065, -5.785675, -8.82605, -9.680984, -7.954941, 
    -7.700256, -6.828903, -2.693222, -5.963028, -14.99245, -29.5388, 
    -18.21249, -10.21484, -8.805725,
  -6.012512, 0.315094, 0.8908844, -4.108337, -7.858322, -6.282028, -4.771606, 
    -1.906509, -3.185684, -12.17708, -25.93489, -35.21823, -29.89427, 
    -19.4086, -13.5849, -13.6651, -13.85651, -14.72134, -15.4151, -18.28647, 
    -16.09116, -14.86302, -15.50885, -16.25391, -12.42578, -7.116669, 
    -4.211197, 0.8963623, 1.363541, 0.6158905, 1.531509, 5.478897, 3.281509, 
    0.382019, 0.2289124, -5.436462, -7.33255, -8.348953, -8.378387, 
    -8.094269, -4.807556, -2.648941, -1.301575, -1.428391, -4.157547, 
    -4.657806, -3.7547, -1.873688, -1.1698, -1.9776, -5.150253, -10.62656, 
    -15.60547, -18.62813, -18.30495, -16.84323, -16.56017, -19.68593, 
    -23.90703, -24.32083, -21.34949, -17.00026, -13.05078, -1.791397, 
    4.195053, 3.324738, -1.222397, -1.452087, -1.034637, -6.041656, 
    -4.263275, -6.538284, -8.078644, -11.0914, -11.33125, -13.64192, 
    -14.56902, -13.10703, -8.78125, -6.717194, -6.601044, -2.989594, 
    -3.560944, -7.789063, -12.69557, -16.40208, -15.87004, -14.37161, 
    -13.37161, -11.1922, -8.206512, -7.658081, -13.17004, -28.29245, 
    -37.25287, -17.65103,
  -23.77187, -13.49896, -7.228897, -8.204681, -10.83151, -19.31535, 
    -18.83516, -8.884369, -2.915359, 2.964844, 1.264587, -1.087753, 
    -3.616409, -4.564575, -6.31459, -9.415359, -10.92915, -12.71979, 
    -12.56979, -12.62631, -11.66536, -9.458588, -6.921356, -4.156509, 
    -1.368225, 3.3638, 2.923706, -0.6461029, -5.073441, -7.966141, -5.829163, 
    -6.062241, -4.850266, -6.595825, -7.750534, -6.355728, -6.179688, 
    -5.402863, -5.003632, -3.890884, -2.052856, -0.7197876, -2.236191, 
    -4.431519, -6.695831, -7.549469, -7.126312, -6.89505, -5.699738, 
    -8.358597, -11.10365, -13.98125, -17.90157, -20.49948, -23.43073, 
    -24.24922, -23.71588, -22.97578, -24.22656, -26.06354, -26.6151, 
    -26.18411, -22.69974, -19.02892, -17.38463, -8.449219, -7.708862, 
    -9.429688, -10.4823, -12.38412, -11.62317, -11.38855, -11.05702, 
    -12.54895, -14.46275, -12.88177, -13.60832, -13.02266, -12.18333, 
    -9.090378, -5.442444, -4.090363, -4.457535, -5.849731, -7.637238, 
    -8.39035, -11.18152, -13.18515, -15.7901, -16.04089, -14.05443, -14.5125, 
    -16.25548, -18.84479, -21.03073, -27.72891,
  -5.983078, -8.061981, -12.16458, -18.24113, -15.78125, -17.20103, 
    -17.34038, -18.48541, -15.19479, -12.18098, -10.44427, -9.415619, 
    -9.647125, -9.642197, -11.12318, -12.72551, -15.06615, -17.09634, 
    -17.73698, -18.34973, -17.83099, -15.35104, -11.78828, -8.585938, 
    -4.983597, 4.057816, 4.082291, 0.9604187, 1.419525, 0.8585968, 0.4966125, 
    -0.2911377, -1.446609, -2.703384, -3.398956, -4.286453, -4.510162, 
    -3.283859, -2.338791, -1.494263, -1.808594, -2.979172, -4.458069, 
    -5.898956, -6.726822, -7.215897, -7.763016, -6.557816, -4.509628, 
    -2.428391, -1.773697, -1.819794, -4.315887, -6.989838, -9.115875, 
    -10.30209, -11.30937, -12.07864, -13.0099, -13.00912, -12.63698, 
    -12.08775, -10.99193, -9.683334, -8.786987, -7.634888, -7.294006, 
    -8.602341, -8.87735, -9.142441, -8.763275, -5.096359, -0.7348938, 
    0.8666687, 0.4296875, -0.2786407, -2.492706, -4.988022, -5.623962, 
    -5.670059, -5.681244, -5.988022, -5.744019, -5.51796, -3.821869, 
    -1.179947, 1.584381, 2.517181, 2.224747, 0.6658783, 0.4145813, -1.116394, 
    -3.375778, -3.477875, -3.668228, -4.33046,
  -5.196625, -5.315094, -5.416412, -4.71875, -3.785416, -3.135941, -2.629166, 
    -1.512497, 0.9247284, 4.173965, 7.646866, 9.18959, 9.956253, 10.37683, 
    10.42188, 9.619537, 7.942459, 5.493484, 3.166656, 1.061203, -1.338547, 
    -3.902084, -5.864578, -7.563797, -9.125778, -10.2276, -10.18437, 
    -8.925781, -7.175522, -4.438797, -1.713272, 0.1799469, 1.824738, 
    3.196091, 3.862762, 4.603653, 5.273178, 5.81041, 6.48645, 6.646866, 
    5.396622, 3.354172, 0.9057312, -1.597656, -4.398438, -7.222916, 
    -9.398956, -10.92371, -11.41328, -11.34583, -11.69505, -12.69531, 
    -13.92682, -15.16199, -16.66589, -18.42656, -19.73151, -21.26823, 
    -22.55598, -23.70729, -24.66823, -25.68359, -26.4263, -27.11874, 
    -26.93307, -27.13516, -27.18282, -26.37161, -24.36302, -21.82603, 
    -18.91719, -15.56017, -13.74167, -12.57083, -11.63124, -11.37474, 
    -11.4711, -12.00339, -12.17969, -12.43359, -13.49011, -13.89531, 
    -13.60208, -13.53984, -14.1375, -14.32683, -14.31485, -13.69661, 
    -12.24635, -10.84766, -9.419006, -8.554688, -7.431778, -6.237747, 
    -5.976303, -5.732285,
  -13.82916, -13.73854, -13.68021, -13.89037, -14.12917, -14.51588, 
    -15.31093, -16.21692, -17.05573, -17.98203, -18.8737, -19.85495, 
    -20.92317, -21.50702, -22.16093, -22.68098, -23.03777, -23.56615, 
    -23.78177, -24.00391, -24.29584, -24.55885, -24.48463, -24.09116, 
    -23.34323, -22.12161, -20.48203, -18.78255, -16.69844, -14.56772, 
    -12.85912, -11.08646, -9.378647, -7.791138, -6.297134, -4.721878, 
    -3.579422, -2.50235, -1.482285, -0.5836029, 0.1065063, 0.4765625, 
    0.6927032, 0.9294281, 1.064056, 1.147919, 1.1875, 0.7484283, 0.2067719, 
    -0.0848999, -0.438797, -0.7677155, -0.7770844, -0.8085938, -0.961731, 
    -1.143494, -1.578644, -1.764847, -1.755478, -1.986191, -2.046097, 
    -2.192703, -2.122391, -1.979691, -1.8591, -1.484634, -1.247925, 
    -0.9208374, -0.2903748, 0.0447998, 0.563797, 0.7054749, 0.744278, 
    0.6328125, 0.3927002, -0.0239563, -0.8638, -1.760422, -2.818741, 
    -4.001038, -5.241669, -6.336456, -7.345047, -8.171875, -9.125519, 
    -10.08516, -11.06979, -11.60521, -12.10339, -12.77499, -13.46014, 
    -13.92422, -14.0229, -14.21538, -14.08958, -13.87032,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.08255211, -0.09166667, -0.1226563, -0.09895831, -0.06822917, 
    -0.05546874, -0.07187501, -0.08854169, -0.07135415, -0.06302083, 
    -0.04609376, -0.04531249, -0.06119794, -0.09401038, -0.09921876, 
    -0.09114581, -0.08645833, -0.07395834, -0.07291669, -0.05989587, 
    -0.04947919, -0.02786458, -0.02135414, -0.03281248, -0.03749996, 
    -0.03125, -0.03619793, -0.02343753, -0.03541666, -0.05052084, -0.0830729, 
    -0.06380209, -0.03984374, -0.03072914, -0.04609376, -0.06484374, 
    -0.0908854, -0.08437499, -0.06119794, -0.03333333, -0.03281251, 
    -0.03411457, -0.03593749, -0.01979166, -0.02760419, -0.04427084, 
    -0.02682292, -0.003125012, -0.01145834, 0.002604157, 0.009635419, 
    0.001302093, -0.01250002, -0.03489584, -0.02708334, -0.01197916, 
    0.006770849, -0.01354167, -0.04270834, -0.05885416, -0.04531249, 
    -0.02500001, -0.02005211, -0.02656248, -0.0390625, -0.03203127, 
    -0.03229165, -0.01354167, -0.02968749, -0.02916667, -0.01119792, 
    -0.02005211, -0.01848957, -0.02161458, -0.0234375, -0.0361979, 
    -0.04869792, -0.06588542, -0.06145835, -0.03333333, -0.02734375, 
    -0.07057291, -0.06354168, -0.04505208, -0.05442706, -0.05026042, 
    -0.04739583, -0.06354168, -0.02109376, -0.01744792, -0.02317709, 
    -0.04609376, -0.04921874, -0.0497396, -0.06458333, -0.07760414,
  -0.8182292, -0.7718749, -0.7158854, -0.4947917, -0.5140624, -0.6356771, 
    -0.7601562, -0.7148438, -0.7385416, -0.6122396, -0.3643229, -0.3070314, 
    -0.3468752, -0.4276042, -0.4695313, -0.5914061, -0.675, -0.7466145, 
    -0.8013022, -0.8432293, -0.8664062, -0.8510418, -0.721875, -0.6611979, 
    -0.6122396, -0.5322917, -0.3903644, -0.1703124, -0.188802, -0.3984375, 
    -0.375, -0.1804686, -0.01041675, 0.09843755, 0.02890635, -0.0140624, 
    -0.1765623, -0.2570312, -0.279948, -0.3278644, -0.2091148, -0.09895849, 
    -0.1367188, -0.09479165, -0.1109374, -0.2765627, -0.1171875, 0.2351563, 
    0.2861979, 0.161979, 0.002604246, 0.05494785, 0.07994771, -0.07291651, 
    -0.2648437, -0.1778646, -0.09114575, -0.1557293, -0.0320313, -0.03723979, 
    0.002343655, -0.0625, -0.1546876, -0.2054687, -0.1966147, -0.08437514, 
    -0.05156255, -0.1427083, -0.1130209, 0.02968764, 0.0846355, -0.0263021, 
    -0.0838542, -0.1979167, -0.1351564, -0.1169269, 0.0888021, 0.2294271, 
    0.175, -0.02161455, -0.2713542, -0.4638021, -0.4197915, -0.5309896, 
    -0.3890626, -0.3031251, -0.2846355, -0.4158854, -0.4744792, -0.4104166, 
    -0.4539063, -0.4385417, -0.5851562, -0.5328126, -0.5348957, -0.6341147,
  -1.771354, -1.630989, -0.8039064, -0.9236979, -1.40625, -1.088282, 
    -0.6184897, -0.1927085, -0.1255207, -0.3028646, -0.4367189, -0.7411461, 
    -0.3658857, -0.07682276, -0.2278643, -0.106771, -0.05156231, -0.2929688, 
    -0.4570313, -0.495573, -0.3804688, -0.1106772, 0.01249981, 0.180469, 
    -0.07265615, -0.2252607, -0.1135416, 0.3484378, 0.2744794, -0.3338542, 
    -0.6546874, -0.1184893, 0.276042, 0.1044269, 0.3377604, 0.4013019, 
    0.09036493, -0.4083333, -0.6679688, -0.578125, -0.4627604, -0.2382813, 
    -0.3929691, -0.6265626, -0.7763019, -0.7283854, -0.3317704, -0.2020831, 
    0.03802061, -0.1226563, -0.2906251, -0.1325521, -0.1929684, -0.3151045, 
    -0.755208, -0.3578124, 0.0661459, -0.598958, -0.7401042, -0.2380209, 
    -0.08463573, -0.4932294, -0.5919271, -0.2583332, -0.3041663, -0.5585938, 
    -0.4510417, -0.09322929, 0.02291679, -0.006510735, 0.03411484, 
    0.07656288, -0.1968746, -0.2523437, -0.09401035, -0.1111979, 0.08203125, 
    0.04010391, 0.1859374, 0.2617188, 0.4333334, -0.5916667, -0.7364583, 
    -0.9393225, -0.4127603, -0.2401042, -0.2294273, -0.1906247, -0.6851563, 
    -0.9716144, -0.5210938, -0.1645837, -0.4286456, -0.5416665, -0.870573, 
    -1.515104,
  -1.804688, -1.236458, -0.2419271, -0.4640627, -1.275782, -1.023698, 
    -0.9981766, -1.307552, -0.7401037, -0.3486977, -0.1622391, -0.09973907, 
    0.2442703, -0.7890625, -0.9796877, -0.3127604, 0.2414064, 0.1463537, 
    0.2151041, 0.9911461, 0.8117189, 0.5432291, 0.948698, 1.53724, 1.601302, 
    0.296875, -0.1661463, 0.06510448, 0.01614571, 0.363802, 0.2018223, 
    -0.02005196, 0.8044271, 0.8492184, 0.2317715, 0.2627602, -0.1320314, 
    -0.2221355, 0.008072853, 0.332552, -0.1835938, -0.2945309, -0.3552084, 
    -1.001823, -0.936718, -0.2489586, 0.5257807, 0.3411455, 0.8497391, 
    0.4505205, -0.391407, -0.709115, -0.6645832, -0.3117189, -1.279428, 
    -1.155729, -0.7109375, -1.12474, -1.097135, -0.5653639, -0.8687506, 
    -1.241406, -0.614583, 0.09375, -0.3328123, -0.5049477, -0.1906252, 
    -0.2234373, 0.296875, -0.4234381, 0.01276016, 0.08489609, -0.3963547, 
    -0.1776047, -0.2763023, -0.3927078, -0.3122396, -0.06979179, 0.2080727, 
    0.2513027, 0.9666662, 0.7276039, 0.4541664, -0.2093754, -0.4401035, 
    -0.4872398, -0.05364609, -0.01458359, 0.467968, -0.6028643, -0.848958, 
    -0.5127602, -0.3656254, -0.2809896, -0.629427, -1.291145,
  -0.526041, -0.7786446, -0.3942699, -1.798437, -1.682293, -0.5020847, 
    -0.1765633, -0.8187504, 0.2002602, 0.374218, 0.3398438, 1.003906, 
    0.7273445, -0.002342224, 0.2085934, -0.4669285, -1.167707, -0.7234364, 
    0.3395844, 1.02422, 0.2627602, -0.1812496, -0.421875, 0.250782, 0.515625, 
    1.210938, 0.7333336, 0.2541676, -0.3463535, 0.09088707, 0.4848957, 
    -0.1270828, -1.286457, -0.2640629, -0.4148426, -0.5585938, -0.9276028, 
    -0.4052086, -0.1697922, 0.1466141, -0.4088535, 0.1104164, 0.8106785, 
    1.145573, -0.270052, 0.4958344, 0.2979164, -0.2687492, -0.4963531, 
    0.5908852, 0.1682281, 0.1390629, 0.8661461, 1.422657, 0.7005215, 
    0.3635426, -0.7216148, -0.2184887, 0.1541672, 0.5062504, -0.6059895, 
    -2.057812, -1.90625, -0.7208347, -0.9296875, -0.724741, 0.1283855, 
    -0.1476555, -0.2986984, 0.9697914, 0.4822922, 1.079687, 0.8395844, 
    -0.1411457, -0.4867191, 0.5023422, 1.160938, 0.2658863, 0.6044273, 
    0.5114594, -0.3981762, -0.06536484, 0.05364609, 0.3773441, 0.2895832, 
    1.25703, -0.3361988, -0.7773438, -0.3515625, -0.4627609, -0.6463547, 
    -0.1557293, -0.6820316, 0.1682301, 0.8916664, 0.823698,
  0.3809891, -1.199741, -1.320572, 0.02447891, -0.5343742, 0.06614685, 
    -0.7341156, -0.3252602, 0.5994759, -0.004425049, -0.4307289, 0.1119804, 
    -0.1747398, -0.9710922, -0.7002602, -0.8315086, -0.7127609, -0.7502594, 
    0.1669273, -0.7322922, 0.1156235, -0.3682327, -0.2065086, 0.3460922, 
    1.461201, 0.1549492, 0.2080727, 2.037498, 2.059895, 2.528387, 2.030472, 
    0.5247383, -0.02447891, 0.4460945, 0.7151031, 0.6388016, 0.6752586, 
    1.838543, 2.362499, 1.72578, 0.1861992, 0.4072914, 1.539322, 2.77578, 
    2.436199, 0.8265629, 1.645836, 2.7612, 1.789063, 2.523701, 3.778908, 
    2.402084, 1.313023, 0.6796875, 1.691666, 2.504688, 0.8447914, 
    -0.02968597, -0.5445328, 1.16901, 1.235939, 0.1731796, 0.5406227, 
    1.557034, 1.110935, -0.6096382, -0.7552071, 1.020309, 1.685158, 1.815365, 
    -0.3666649, -0.6414032, -0.1484375, -1.454948, -0.7117195, 1.273439, 
    1.009113, -0.9518223, -1.006767, -0.5369759, -1.543751, -0.7606773, 
    1.074738, 2.78672, 1.893227, 2.469791, 1.343227, 0.6458321, 1.636982, 
    0.389061, -1.691929, -1.459637, -0.01327896, 0.2791672, 0.2843742, 
    0.1971359,
  -0.09218597, -2.11068, -2.176304, 0.4609375, 1.094269, -1.01302, -1.935154, 
    -2.588543, 0.7289047, 2.497395, 2.392971, 1.271091, 2.158855, 0.8020859, 
    -0.2296906, -1.805729, 0.471096, 3.002342, 1.162502, 0.1098938, 
    0.5447922, 0.5354156, 0.5041656, 2.52005, 3.985157, 2.739586, 2.71875, 
    3.030731, 3.622135, 1.047134, 0.359375, 1.401566, 2.103386, 0.4406242, 
    0.842186, 1.45182, 0.7789078, 1.830208, 1.905468, 0.7718735, -0.08020782, 
    -0.4080734, -0.5291672, 0.9882813, 2.360676, 0.9484367, 2.56406, 
    5.417446, 4.248959, 2.686722, 1.815887, 2.894531, 3.28828, 1.465626, 
    2.140362, 1.940884, -0.3174477, 2.928646, 1.407295, 1.114845, 2.33802, 
    1.541668, 1.091404, 2.496616, 1.446354, 0.9796867, 0.2497368, 0.9502602, 
    0.6968765, -0.3434868, -1.108593, 2.723957, 0.830471, -0.6911469, 
    2.175003, 3.134373, 0.6911469, 0.2138023, 0.2580719, 0.3838539, 
    -1.032551, -0.7432289, 1.178127, 1.458591, 0.4315109, 0.3419266, 
    1.439323, 1.644794, 2.599998, 2.092968, 0.4192696, 0.3476563, -0.904686, 
    -0.3164063, 0.8622398, -0.4145851,
  -1.639843, -0.2705727, 2.402084, 1.882553, -0.8343773, 0.2005196, 
    -0.6585922, -0.05416107, -2.171875, -0.6020813, -0.5132828, 2.406509, 
    1.992973, 1.563278, 2.343231, 2.103645, 0.5273438, 0.1138, 0.8492203, 
    1.030727, -1.185936, 3.298958, 4.441143, 3.377602, 5.790886, 6.763283, 
    5.689583, 1.160942, 1.550522, 1.185417, 0.2690086, 2.490887, 3.944271, 
    1.492706, 2.03334, 3.22057, 2.777607, 1.733593, 2.827866, 0.6395798, 
    0.4320297, -0.8255157, 1.227341, 1.313282, 1.295311, 0.4458313, 
    0.3195305, 3.107033, 4.175262, 4.93203, 4.364059, 3.525002, 3.966148, 
    1.702084, 2.08073, 2.924999, 2.936718, 2.513283, 1.720051, 2.237759, 
    3.879948, 3.365887, 3.483074, 4.533073, 3.714062, 3.815887, 3.660938, 
    -0.4869804, -1.011978, 1.185677, 3.403645, 3.569271, 1.31953, 2.205208, 
    2.86953, 0.6164017, 0.3489609, 1.819271, 1.396095, 0.07343292, 0.7341156, 
    0.3151016, -1.699997, -1.460415, 0.07421494, -1.080986, -0.8684883, 
    -1.631771, 1.419533, 2.105469, 3.386978, 4.113277, -0.1479187, 1.159634, 
    -1.269531, -3.504166,
  2.4487, 1.584381, 2.578125, 1.400261, 3.476822, 2.818748, 3.38932, 
    2.743225, 1.094536, 3.071877, 7.070045, 8.240105, 7.511192, 8.025261, 
    8.17318, 6.699478, 6.467712, 4.477608, 3.43412, 2.055992, 3.34375, 
    2.802345, 2.373444, 3.115883, 1.172653, 0.3617172, 1.800781, 2.397133, 
    0.828125, 1.609116, 3.709373, 4.660942, 3.59037, 2.893227, 1.793747, 
    0.170311, 2.704163, 1.112236, -2.281509, 0.7927094, -2.26432, -2.67318, 
    -3.272919, -2.087234, 0.0231781, -1.157036, 1.383072, 7.296097, 3.877861, 
    4.893227, 7.173439, 4.81041, 4.270576, 2.259895, 4.70443, 2.697914, 
    1.731773, 2.521614, 0.9713516, 1.836723, 2.809639, 3.978905, 4.061203, 
    3.385933, 2.759377, 1.362755, -0.2083282, -0.5987015, 0.734375, 
    0.3062515, -1.815109, -1.771873, -2.234375, 0.05364227, -0.6296844, 
    -0.1997375, 2.055992, 3.032547, -1.767181, -3.011719, 1.056511, 
    -0.2932281, -1.75, 0.2354202, 0.2908859, -2.11953, 1.9086, 2.219528, 
    2.396873, 3.241928, 1.850258, 3.379951, 3.639839, 0.9768295, -0.03020477, 
    3.428383,
  3.052086, 1.246872, 1.193748, 4.102859, 4.698441, 0.529686, 3.025261, 
    1.530464, -0.1575546, 3.29557, 7.945572, 6.652344, 6.074738, 5.91198, 
    7.403389, 8.0289, 6.46875, 1.976303, 1.790886, -0.391922, -0.1916656, 
    -0.6026077, 1.22995, 0.4234314, -1.811722, -2.423965, -3.035942, 
    -0.8682251, -0.4408875, 2.300781, 5.315369, 5.158073, 2.078384, 
    -5.214577, -5.201561, -8.717445, -6.719009, -3.046097, -8.608856, 
    -9.515625, -8.184631, -9.303383, -2.573181, -1.016403, -0.8062515, 
    0.8554688, 3.935417, 6.318748, 4.826828, 4.439064, 4.648178, 0.8679657, 
    0.1635437, -0.7223969, 2.785942, 0.9765625, -0.7593765, 1.574997, 
    2.261192, 2.660156, 2.136719, -0.1140671, 1.830208, -0.6513062, -2.5513, 
    -2.513023, -2.967705, 0.9158859, 0.7770844, 1.485939, 1.450523, 
    0.9989624, -1.858337, 2.214844, 0.2463531, 1.41198, 2.5961, -0.6020813, 
    -1.93177, -3.231514, -0.9278641, -1.195572, -0.3226547, -1.608589, 
    3.2388, 1.582809, 5.527344, 2.120827, 5.024734, 1.013542, 2.175522, 
    1.932289, 3.274223, 2.972137, 2.3237, 2.924217,
  1.009377, 1.168488, 1.126564, -0.3575592, 0.8799438, 0.6682281, 6.39843, 
    3.385422, -1.442711, 4.784119, 8.515366, 3.384109, 4.986725, 8.395576, 
    5.015106, 4.657555, 4.170311, 5.980209, 2.781509, -3.032028, -2.529694, 
    -1.328125, -3.454422, -1.466667, 2.199738, -1.214317, -2.157814, 
    -4.133858, -2.20443, 1.867188, 5.262497, 0.3187485, -13.66875, -17.57344, 
    -12.12057, -10.78359, -15.74271, -18.26406, -15.44297, -13.65495, 
    -10.9625, -6.496613, 3.860931, 4.565102, 4.55365, 4.823959, 5.527863, 
    1.680733, 2.960938, -2.245834, -1.947395, -0.4940109, 1.667191, 
    -0.7598953, -2.582817, -4.620567, -3.748695, 1.187241, -0.6632843, 
    -0.2976532, -3.010155, -3.8862, -5.006248, -3.938019, -2.649483, 
    -2.210678, -3.323174, 0.3192673, 1.774742, -2.395576, 0.05937958, 
    -0.985939, -1.90078, 3.159378, 1.580208, -1.571106, -2.489319, -2.933594, 
    -5.507813, -1.992188, 0.1166687, 3.524742, 3.20417, 2.52552, 4.593231, 
    3.267448, 5.360939, 2.29583, 0.8385391, 3.073952, 4.081512, 1.514839, 
    1.625786, 3.194016, 2.281776, 0.8994827,
  1.460938, 0.8460999, -2.774475, -0.8635406, -2.726822, 0.3611908, 3.642715, 
    1.931778, -0.8447876, 1.004166, 3.197662, 5.208328, 1.598175, 0.1882782, 
    3.514847, 5.528641, 3.407036, 1.578651, 2.582558, 2.996353, 0.3515625, 
    -0.7916641, 2.323692, 0.1695251, -0.1544266, -3.089058, -5.823433, 
    1.463799, 5.067703, 3.979172, 1.642181, -0.9651031, -12.35104, -16.28281, 
    -16.36667, -20.22057, -24.73568, -23.65755, -16.69921, -10.06511, 
    -3.588806, 2.358856, 4.299728, 5.313797, 3.754433, 0.1541672, 5.027603, 
    1.279686, 0.5606766, 0.3151016, 2.265884, 2.082817, 1.472916, -2.86953, 
    -5, -1.781509, -1.029953, 0.03020477, -2.596092, -4.768753, -4.064583, 
    -4.28125, -3.336975, -2.290619, -2.921097, 0.4020844, -3.085938, 
    -4.268234, -2.63385, -2.375, -1.939323, -3.440102, -2.342445, -1.591148, 
    -0.2406311, -2.346863, -4.650269, -6.979691, -5.860672, -1.830475, 
    5.058334, 10.50807, 10.21614, 9.215622, -1.473961, 2.078903, 4.664841, 
    3.464584, 4.585159, 0.744278, 0.9148407, 1.342194, -0.6161423, -3.288536, 
    -1.589584, -2.166145,
  -4.005463, 0.3684845, -0.7283783, -2.374222, -2.624481, 1.694519, 5.876572, 
    3.858582, 6.421616, 3.820045, 0.2658844, 5.937759, 0.9203186, 6.845833, 
    1.062241, 1.090103, -1.217972, 2.447403, 3.239594, 1.798706, 1.713806, 
    1.435684, -1.124222, -4.216934, -5.608856, -1.627335, 0.5179749, 
    -0.4994812, 5.585678, 1.787766, -2.388016, -4.4487, -7.14505, -18.39009, 
    -15.49948, -11.55313, -11.76459, -14.12083, -9.061188, -1.474747, 
    4.971619, 2.382553, 1.610168, 3.683594, 2.360931, 1.459885, 1.274734, 
    4.515366, 8.472656, 8.478653, 5.339844, 4.633865, -0.160675, -3.2164, 
    -1.302338, -2.434113, -4.397919, -3.114059, -3.815353, -3.971085, 
    -0.3494873, -0.5697937, 3.082306, 5.027084, 0.07240295, -2.584122, 
    -2.787247, -5.906769, -2.028122, 1.914841, -0.4523468, -0.4304657, 
    1.411209, 2.983856, -0.7401123, -13.66171, -8.023956, -7.000778, 
    4.248703, 6.660942, 9.316666, 13.35991, 9.375259, 12.79036, 7.669533, 
    10.2013, 3.754944, 1.161209, -1.691406, 2.973969, -1.494797, -5.779175, 
    -4.74324, -1.622147, 0.3416595, -1.602875,
  3.22995, 2.075256, 0.6723938, -3.132034, -3.82605, 3.115097, 4.719528, 
    6.455719, 11.31822, 4.455734, 10.77708, -4.121628, -2.624481, 5.014053, 
    0.9127655, -4.436203, -0.6351624, 1.238281, 7.206253, 3.171875, 3.414581, 
    1.654434, -1.676041, -4.387756, -3.393753, -0.1161346, 0.8401031, 
    -0.6869659, 2.079422, 3.835678, 2.426575, -4.497925, -4.914581, 
    -6.758591, -6.877869, -6.182556, 0.5583344, -3.764847, 0.8247375, 
    10.08177, 7.613022, -0.4010468, 3.399216, 7.142975, 6.827866, 1.155472, 
    3.246353, 3.452347, 4.400009, 0.7658844, 0.09817505, -1.56485, -6.417709, 
    -5.289063, -3.140106, -1.255219, -4.289841, -0.3408966, 1.115616, 3.7099, 
    9.081253, 5.660934, 0.6989594, -1.412231, 0.2526093, 0.4382935, 1.253906, 
    0.6026001, 0.6763, 6.831238, 6.09584, 5.846359, 5.69635, 2.9888, 
    -8.369537, -2.811722, -3.980469, 0.6390533, 12.31068, 15.24191, 14.25677, 
    6.996094, 5.873428, 3.033859, 20.24635, 19.54089, 0.5791626, 1.400528, 
    0.1773376, 1.929688, -8.592194, -4.432541, -4.363281, -2.127869, 
    -2.143478, 0.05052185,
  8.590103, 3.679169, 0.401825, -2.945572, -4.785675, 2.244537, 0.4968719, 
    7.822647, 12.71718, 11.03073, 12.15416, 2.385681, -4.279953, -4.12265, 
    4.696091, 5.584106, 1.17421, 4.192184, 1.906509, -1.399475, 1.615097, 
    0.3455811, -2.441666, -2.400269, -1.636459, -3.963806, -4.767441, 
    -4.061203, -2.583069, -2.383591, 0.1989594, 2.140884, -0.7393188, 
    -3.008347, -5.746872, -4.74765, 0.6010437, -3.283325, 3.226044, 8.016144, 
    -0.2622528, 4.15416, 8.516403, 7.297394, 5.540375, -2.674225, 3.304153, 
    2.171356, -0.9666595, -2.375519, -0.6479034, -2.325516, -3.711716, 
    -0.8627625, -2.256516, -1.738541, 0.2028656, 1.421616, 2.495834, 
    3.674744, 3.183334, -0.2841187, -0.129425, -0.6130219, 2.005203, 
    0.1320343, 5.345322, 8.485153, 9.33905, 7.671616, 7.932816, 7.225266, 
    8.096603, 3.88385, -1.534897, -4.376038, 5.952087, 11.36198, 8.990891, 
    15.1763, 14.25911, 3.944534, 4.697647, 0.5112, 17.09662, 13.79584, 
    -1.835678, -3.873962, 2.456253, -2.65416, -4.567444, -1.314575, -4.4888, 
    4.216919, 0.2044373, 6.45079,
  8.960678, 7.218491, -2.21875, -8.604431, -5.389572, -3.605209, -4.996872, 
    -4.254944, 2.741409, -4.608337, 9.091156, 9.232285, 4.649216, 5.812241, 
    3.943741, 8.513809, 4.238022, 3.62709, 7.561707, 9.148972, 9.245041, 
    5.579681, 1.747391, 0.2979126, 1.526306, 4.540619, 3.309631, -1.815369, 
    0.04244995, -2.61171, 0.2249908, 0.4518127, 1.895325, -2.108597, 
    -4.927353, -4.757294, -2.510162, -5.561188, 0.3036499, 1.188797, 0.65625, 
    0.2971344, 5.243759, 0.8278656, 1.808594, -5.501816, -2.083069, 
    -2.458603, -7.624222, 0.3609314, 2.754166, 2.692184, 0.4505157, 2.333084, 
    -0.008865356, -2.3013, 0.2911377, 1.591415, 3.10704, 2.777084, 4.741409, 
    5.60704, 3.093231, 3.194794, 2.895584, 6.286728, 6.186188, 5.760925, 
    6.523438, 3.869278, 6.886719, 7.944794, 9.1315, 8.64296, -3.416138, 
    -4.844528, 10.13048, 15.40521, 4.246887, 9.325775, 7.120834, 3.37709, 
    8.867966, -0.2447815, 5.8638, 10.05391, 12.80156, -5.0672, -6.172134, 
    -7.1138, 0.06381226, 2.096619, 2.082809, 7.630722, 7.577606, 6.881241,
  1.521088, -3.913544, -10.07866, -8.176041, -9.767181, -8.447647, -8.413269, 
    -10.25285, -4.887497, 5.638535, 16.55547, 17.75313, 2.991928, 5.545822, 
    8.409637, 7.103912, 6.522919, 6.958069, 6.232285, 7.578384, 5.753647, 
    4.308853, 0.3744812, 1.523956, 5.806778, 7.536972, 4.365631, 2.514847, 
    11.06641, 4.998688, 0.03489685, 2.511185, 8.038803, 5.947403, 4.734634, 
    3.302856, -4.075256, -16.5302, -4.887238, -0.3562469, -6.969009, 
    -3.708328, 2.564331, 5.489838, 4.564316, 3.223953, 6.905991, 1.575775, 
    -3.988022, -5.345322, -2.536987, -1.040115, 2.150528, 3.361465, 
    -2.449219, 0.0929718, 0.3468628, 2.611725, 4.100525, 4.162766, 5.030991, 
    6.304428, 6.637772, 6.336197, 5.863281, 2.929947, 6.858337, 7.403122, 
    8.3974, 7.906769, 8.566666, 8.615112, 2.729691, 5.310944, -5.295578, 
    2.175247, 12.04506, 5.340622, 14.63855, 15.83308, 12.42056, 8.630737, 
    5.922653, -1.110672, -10.04193, -2.011978, 8.832809, 2.648956, -3.093231, 
    -5.2789, 1.090622, -2.213547, 1.492188, 3.213547, 7.403397, 2.0672,
  0.0252533, -0.7554626, -2.471085, 1.0737, -11.7289, -13.08855, -11.78021, 
    -16.58072, -12.19714, -9.857559, -4.535934, 24.25417, 16.63907, 4.421616, 
    6.933853, 5.199478, 6.126572, 4.106766, -0.1552124, 2.199738, 0.9791565, 
    -3.756256, -4.532547, -1.657028, 1.81485, 4.364578, 6.980988, 11.52995, 
    0.6117249, -1.540634, 6.472137, 14.48021, 20.02344, 3.978638, -1.967453, 
    7.253387, 7.322922, -0.5307312, -3.76355, -6.167191, -4.063797, 
    -1.807541, -2.532822, -5.275513, -4.783081, -1.638535, -4.028381, 
    -8.337234, -17.09453, -25.42787, -28.50363, -23.46094, -20.80183, 
    -13.65547, -12.55052, -12.03542, -9.790375, -6.815887, -3.282288, 
    -1.462769, -0.4388123, 1.223953, 4.590363, 5.470306, 3.692703, 1.615631, 
    6.159897, 2.525528, 3.876038, 4.482819, 4.33255, 1.670578, 2.332565, 
    2.121353, -8.542191, 2.904953, 20.21666, 18.12969, 12.32918, 9.457809, 
    15.41615, 17.99011, 16.18776, 14.51511, 11.95442, 18.67995, 13.88776, 
    2.119003, -2.104156, 1.845322, 6.175522, 1.298706, 3.903915, 2.489334, 
    6.241653, 2.53334,
  -1.952606, 1.359375, 0.865097, 6.118759, -0.2716064, 1.209122, 4.139587, 
    -5.744797, -5.025253, -15.66432, -12.30833, -2.015106, 17.55859, 5.07605, 
    6.082016, 5.109375, 5.196869, 4.248184, 1.311203, 0.714325, 0.2481689, 
    -1.986984, -3.880737, -5.220825, -6.101303, -2.120316, -0.3247375, 
    0.8312531, -7.799484, -7.1297, 1.182556, -7.106247, -18.23958, -12.256, 
    -4.923706, -1.111725, -0.441925, -3.534378, -2.39505, 0.1677094, 6.11615, 
    3.017441, 1.358078, -7.849213, -5.272659, -1.369797, 3.629959, 0.688797, 
    -1.962769, -1.829956, -5.299728, -8.590881, -7.729156, -6.275787, 
    -7.143234, -5.951569, -3.238037, -4.082275, -3.004456, -2.044556, 
    -3.007568, -4.111725, -3.014313, -1.92865, -0.9710999, -1.830719, 
    0.3273621, -0.6148376, 3.016663, -0.2364502, -2.863022, -4.605209, 
    -12.5224, -18.59193, -25.17683, -5.116135, 8.1474, 1.871094, 10.91119, 
    10.73855, 6.105209, 18.75261, 39.54271, 31.97917, 29.8698, 26.57657, 
    16.66849, 4.940369, -1.81041, 2.542969, 11.77266, 12.23125, 9.888275, 
    3.625, 1.994781, -1.78125,
  7.114059, 6.842453, 15.90833, 12.73906, 10.77031, 6.289063, 13.68202, 
    18.19193, 18.50417, 10.45937, -6.574478, -8.140106, 8.525238, 13.23697, 
    4.800262, 4.462219, 8.9888, 4.874222, 2.671875, -3.29921, -4.852081, 
    -6.1828, -10.50002, -8.348694, -10.50389, -2.922668, 0.2166748, 
    -12.77682, -8.163025, -0.1005249, -6.400772, -8.540359, -12.22343, 
    -8.574219, -7.62265, -4.254944, -1.666138, -4.066666, -3.053909, 
    -2.692459, 7.456253, 7.989594, 6.961456, 2.481781, 0.3434906, 4.478897, 
    12.62292, 13.20651, 10.57996, 12.42474, 13.19167, 11.02316, 9.828903, 
    7.015625, 7.009644, 8.126038, 5.286972, 1.592438, 6.280472, 3.807816, 
    4.354172, 2.732819, -0.1598969, 0.6070251, -5.138794, -7.014572, 
    -5.740372, -4.155731, -5.454178, -4.623703, -5.853394, -20.12344, 
    -20.29193, -15.60001, -5.805984, 2.027863, -0.5804749, 2.232033, 19.575, 
    22.98099, 14.94324, 17.81772, 15.07526, 12.675, 13.2823, 4.163284, 
    4.734894, 2.360428, -0.9916687, 3.896103, 3.738281, 6.811203, 5.155212, 
    -2.744278, 8.313019, 8.801041,
  15.24583, 18.88853, 17.09999, 13.87215, 8.044525, 7.569, 6.138809, 
    13.50859, 17.28932, 28.35938, 18.00235, -7.323181, -0.9234619, 2.041168, 
    0.1789246, -2.453125, -1.233093, 1.067169, -3.072403, -2.75235, 
    -1.537262, -8.190628, -19.63022, -13.95131, -11.24818, -8.230209, 
    -5.704681, -2.970047, -10.97891, -16.85963, -9.441147, -4.098175, 
    -5.227341, -3.515366, -6.759644, -4.671097, -5.864334, -5.882553, 
    -9.847916, -9.429688, -0.3880157, 5.706512, 3.796875, -0.96875, 
    -2.128632, 2.458328, 1.891922, 2.237762, 1.118759, 1.813278, 3.666412, 
    3.758072, 1.999207, -0.2914124, -0.7612, 0.6140594, -1.059906, 1.413544, 
    1.588547, 0.4692688, 4.507813, 11.83568, 10.53697, 8.100784, 2.681778, 
    5.170044, 6.124481, 4.027603, 0.3510437, 10.8914, 1.110947, -8.592712, 
    -6.122131, -1.792175, 3.04454, -2.119003, 5.678131, 13.50781, 7.5, 
    9.442719, 3.754669, -0.6729126, 1.1651, 5.629944, 3.765106, -0.6773529, 
    3.34584, 0.4614563, 3.847137, -1.567184, -0.2773438, -1.775009, 
    -3.833847, 13.99609, 15.31561, 18.87917,
  8.483597, 6.897919, -0.9031372, 0.7770996, 2.917175, 5.689575, 0.4221497, 
    1.353668, 5.466431, 6.399994, -0.3221436, -4.059113, -1.625519, 
    -4.549744, -3.808075, -0.6320496, -4.979431, -1.498718, -2.961212, 
    -2.032288, 2.251831, -16.17317, -21.4021, -27.46275, -17.6362, -8.151306, 
    3.916931, 17.91432, -1.697922, -12.29454, -4.952087, -0.5528564, 
    -5.240112, -0.1885529, -3.890106, -0.5117188, -5.807816, -13.63046, 
    -11.13568, -7.555206, -4.470047, -6.074997, -4.246094, -3.400269, 
    0.7674561, -0.4296875, 1.24765, 3.389832, 3.951813, 1.696106, 4.698944, 
    3.194275, 0.5481873, 3.283081, 2.665894, 2.024231, 0.1411438, 3.900543, 
    4.077606, 8.646362, 8.073181, 4.993744, 3.407043, 1.311981, 5.302368, 
    4.555725, 9.012238, 6.269531, 6.631241, 12.91849, 3.856522, 1.982544, 
    9.671875, -3.025787, -15.1552, -13.43961, -10.42682, -7.916656, 
    -6.701843, -13.40314, -7.603119, -1.79454, -2.530731, -4.208069, 
    -1.47995, 2.562759, 2.580734, 4.528641, 2.258087, -0.2320251, -1.871338, 
    -8.676575, 7.4953, 13.50076, 9.3414, 9.79686,
  5.086731, 3.457031, 1.159119, 0.8395691, 0.0078125, -1.517975, -0.8796997, 
    -2.113525, -4.671875, -3.061737, -2.398163, -4.262756, -3.662506, 
    -7.099213, -7.684387, -6.822662, -4.517181, -9.246857, -7.561188, 
    -6.581512, -11.29062, -21.51978, -16.74115, -13.49687, -20.09558, 
    -6.374222, 13.68933, 12.05598, -0.9627686, 1.223694, 7.995575, 11.25807, 
    8.036209, 1.079437, -0.04452515, -2.444794, -9.206268, -12.56691, 
    -6.594788, -3.392181, -0.8817749, -1.749237, -0.4249878, 0.7942505, 
    3.583344, 0.638031, 1.566406, 3.847137, 2.024994, 5.396088, -1.31665, 
    -1.993774, -0.0687561, 4.1698, 3.2836, 4.900772, 5.310425, 6.81041, 
    11.30154, 15.83853, 13.25989, 15.65234, 16.66458, 12.24219, 16.77682, 
    8.059875, 7.062744, 9.074219, 6.578644, 14.15182, 17.68178, 32.99323, 
    27.23021, -3.019531, -9.493774, -15.50729, -12.98019, -12.56796, 
    -11.68204, -4.928406, -3.925018, -9.110931, -8.815872, -3.627869, 
    2.052597, 1.93985, -1.289063, 6.621613, 2.360168, -0.8513184, -2.709106, 
    -2.931519, 3.18045, 12.24924, 12.93777, 8.255463,
  9.309387, 9.87085, 7.142181, 3.101044, 1.451569, 0.5612183, -0.02474976, 
    -2.00885, -3.288788, -3.4216, -3.614594, -2.548431, -5.491394, -6.527588, 
    -11.44974, -15.62524, -13.74088, -2.410156, -10.57266, -10.92578, 
    -10.58646, -18.0672, -24.84531, -13.15938, -5.933594, -6.749222, 
    -1.729691, -15.45547, -6.713028, -1.910934, 4.793472, 5.863022, 9.11145, 
    10.37056, 6.808594, 1.077087, -7.030487, -5.298157, -2.192719, -3.619263, 
    0.8971558, 6.491669, 3.507813, 1.857056, -0.8648376, 0.5161743, 
    -0.234375, -1.792725, -4.100006, -1.373444, -2.224487, -0.6002502, 
    -6.442444, -2.526306, -1.628662, 1.858063, 3.137253, 6.696884, 6.466156, 
    12.3672, 11.04193, 12.91016, 11.9823, 10.8909, 7.703644, 5.135925, 
    6.474731, 2.220306, 7.448181, 17.00626, 28.16849, 20.32111, 17.17136, 
    -2.531769, -2.326843, -8.652588, -5.948151, -5.591675, -7.25235, 
    -10.19662, -7.306244, -3.930206, -1.980988, -6.68985, -1.934906, 
    1.932556, 2.0065, 6.311462, 6.547913, 4.765106, 0.4085693, -1.421875, 
    0.7867126, 9.156769, 15.54529, 12.59247,
  8.558594, 10.91119, 17.35156, 9.021118, 7.274994, 7.972931, 2.509613, 
    -0.0760498, -1.418243, -2.369537, -3.246338, -2.050262, -1.2388, 
    -4.610962, -7.602112, -11.36743, -15.58618, -13.5672, -18.3078, 
    -14.68622, -11.10522, -16.34531, -15.59247, -20.46799, -16.35704, 
    -22.17995, -18.36017, 1.992188, 5.222656, -1.924744, 7.421875, 11.00052, 
    14.54477, 24.44923, 16.33463, 8.658081, 6.216919, 4.609375, 6.98465, 
    4.721893, 7.456757, 3.160156, -2.271881, -4.840363, -0.877594, 1.494537, 
    -0.1268311, -2.553925, -2.020569, -2.202362, -4.206482, -4.619019, 
    -3.48175, -12.13541, -7.090881, -3.160675, -2.79245, -2.239319, 
    -1.049744, 5.383881, 6.11145, 1.029663, -2.433868, -1.499207, -2.2388, 
    -5.855225, -6.063812, -3.766144, -2.164581, 6.658325, 8.510162, 
    0.9494934, 3.0354, -0.2007751, -4.015625, -1.592468, -0.6148376, 
    -3.467987, -1.926056, -2.973175, -5.060669, -5.391663, -7.926056, 
    -7.327087, -2.632538, -4.127625, -5.219269, -1.244019, -1.776306, 
    4.256531, -2.7659, -0.6104126, -0.1755066, 3.029449, 7.493744, 9.992706,
  4.450531, 4.456238, 7.091125, 9.454163, 11.22995, 8.867981, 3.278381, 
    0.4559937, -0.6955872, -1.633575, -2.991394, -2.130463, -1.733063, 
    -2.581238, -4.517456, -6.933838, -6.745056, -7.891144, -8.857819, 
    -11.17059, -10.93176, -18.10156, -30.07083, -18.95206, -19.33932, 
    -20.56511, -8.708328, 10.44115, 20.32213, 10.48151, 6.018494, 5.126556, 
    13.78177, 13.37915, 11.49426, 6.866669, 3.162231, 3.665375, 8.560944, 
    8.897675, 8.802887, 2.963531, -8.278656, -9.047394, -7.301819, -4.2146, 
    -2.83255, -2.008331, -6.773712, -8.443756, -7.268494, 2.601318, 3.687744, 
    -0.7903442, -0.6239624, -2.035675, -5.264557, 0.3890686, -6.2547, 
    -6.020325, -3.865112, 0.006744385, -4.817719, -5.883362, -16.20624, 
    -11.0625, -10.00858, -7.420044, -6.036743, -9.82135, -5.033051, 
    -6.591644, 0.9369812, 0.5031433, 7.809906, 4.140106, 5.455444, 4.988281, 
    1.188019, -4.873718, -2.422394, -2.530731, -3.526825, -1.647675, -1.8508, 
    -5.573181, -5.7453, -4.003662, -7.161194, 1.603119, 3.784637, -6.515381, 
    3.739594, 1.867432, 2.626831, 4.788544,
  2.689819, 5.459106, 7.953888, 4.557037, 7.195831, 4.809113, 6.257813, 
    6.127869, -0.8713379, -1.53125, 2.47995, 0.5255127, -2.380463, -1.152344, 
    -0.4010315, -4.638794, -3.148682, -3.650269, -7.278656, -6.819275, 
    -9.505463, -16.2406, -29.84946, -16.66251, -16.09143, -21.87265, 
    -18.85599, 0.9484406, 8.976044, 10.19426, 6.568237, -4.402084, -9.468231, 
    -5.126556, 0.6744843, -4.246109, -4.581253, -4.751297, 0.8536377, 
    6.342453, 10.16693, 4.9039, -4.701813, -5.570587, -4.902344, -4.056488, 
    2.0849, -1.055969, -5.169006, -6.29895, -4.295837, -2.991394, -0.9536438, 
    -3.602356, -0.9898376, 0.5427246, 1.564331, -0.4070129, -2.4711, 
    -5.65155, -4.650238, -4.73465, -0.9710999, -12.11356, -5.426819, 
    -8.590607, -11.069, -4.987244, -10.94843, -11.72891, -11.20834, 1.7565, 
    1.527863, 1.192963, 7.273712, 0.8335876, -1.826813, 3.441406, 0.3078003, 
    -0.7216187, 1.180725, 3.125519, 3.510925, -1.340637, -0.491394, 0.984375, 
    2.898438, -4.349762, -6.619781, -5.372131, -5.917725, -0.8559875, 
    -9.063782, -0.05807495, 2.562225, 8.3414,
  9.099731, 12.52917, 16.33334, 6.590363, 5.526581, 4.519287, 8.179962, 
    5.665619, 12.91095, 4.845062, -0.2627563, 1.358582, 2.716644, 9.516693, 
    6.179688, 0.6531372, -0.7814941, -2.423462, -7.051056, -1.9888, 
    -0.5770569, -6.703644, -2.142456, -0.3539124, -12.16458, -7.065887, 
    -10.28568, -5.458862, -4.765106, -9.381241, -10.08907, -5.735168, 
    -8.219025, -15.16328, -11.04453, -13.05965, -16.77238, -15.71564, 
    -9.301804, -6.329422, -4.2052, -6.772659, -3.386993, 0.5729065, 
    -1.577866, -2.683838, -3.191925, -1.186707, -5.086975, -4.891663, 
    2.54715, -0.9309998, -2.946625, 3.019806, 1.552368, 0.2614746, 0.7888184, 
    4.147156, 2.159393, -0.1338501, -2.037476, -3.966125, -2.818481, 
    -2.109131, -3.1763, -4.60495, -6.444244, -6.969543, 1.76355, 1.669281, 
    -0.6273499, -1.23645, 3.036438, 4.252075, 5.885925, 2.676544, 4.159119, 
    3.304688, 1.030212, -0.1781311, 1.466156, 0.953125, -1.997406, -5.748169, 
    -3.072144, -2.751556, -6.542725, -7.034119, -1.6922, -5.981506, 
    -3.412231, 4.208069, -0.4080811, -2.871368, 5.418762, 11.5,
  15.68384, -0.09817505, 5.815125, 14.73022, 10.00912, 12.32916, 17.99948, 
    14.04193, 17.15262, 22.46716, 13.54034, 13.34894, 18.67422, 16.75363, 
    2.630463, 5.478912, 4.722382, -2.817963, -7.049225, 3.081512, -5.438293, 
    -1.815613, -2.459106, 1.434113, -1.569794, -5.672913, -3.642456, 
    3.921326, -1.117981, -7.999207, -12.444, -14.81458, -10.03125, -10.68333, 
    -7.908585, -8.759644, -8.594788, -6.943237, -14.18439, -14.77422, 
    -11.16692, -5.34375, -7.302353, -3.683594, -4.163284, -9.149475, 
    -0.7072906, 1.152084, -0.4658813, -1.954163, -4.005981, -1.614319, 
    3.730469, 5.194, 2.564316, -1.121613, -0.870575, 5.683594, 4.428375, 
    -2.270325, 4.164337, 0.5549622, 3.773956, 1.003632, 2.260925, 5.432831, 
    2.761475, -5.802582, 4.385162, 8.623169, 5.108856, -0.2966003, 4.130219, 
    7.285706, 11.71484, 8.633591, 0.8859558, -1.502075, 5.585175, 7.697632, 
    9.035431, 8.980743, 6.959656, -5.088043, -10.96719, -22.63596, -17.07007, 
    -13.18698, -7.4216, -1.610931, -1.6763, -5.038025, 1.764862, 6.730469, 
    8.404694, 16.88281,
  17.07292, -2.085144, 8.82785, 17.20468, 5.000793, 13.49142, 8.624466, 
    -1.708588, -3.188538, 0.588562, -1.613831, 10.29713, 9.8815, 0.9328308, 
    3.885437, 2.961975, 3.179932, -1.998688, -7.037476, -3.897888, -5.561707, 
    -2.757568, -6.020294, -8.437225, -6.67865, -7.113281, -5.783875, 
    -8.12735, -8.025543, -4.328369, -2.374207, -2.750275, -0.2367249, 
    1.766937, 6.052597, -0.4179688, 4.227081, 5.467682, 1.122925, -4.500519, 
    -6.713806, -13.22343, -14.40338, -10.51276, -7.064316, -8.893494, 
    -5.373688, -2.712753, -1.228378, -4.918488, -7.112503, -7.165359, 
    2.48671, -4.83699, -4.999741, 4.679947, -0.220047, 3.496613, 3.496872, 
    3.101044, 3.304688, -2.686218, -0.60495, 5.754974, 11.79034, 15.87631, 
    12.45157, 9.392975, 10.54062, 8.646088, 4.364838, 3.47525, 5.340118, 
    11.09869, 8.349213, 14.1086, 8.307556, 0.2606812, 3.293213, 7.020813, 
    -2.10495, -2.206512, 0.282547, 3.244537, 0.7382813, -10.34505, -13.95337, 
    -9.808075, -8.403381, -0.9724121, 2.974213, -7.1987, -5.079956, 12.67813, 
    26.90417, 41.45026,
  0.7028656, 2.6315, 22.70209, 15.17267, -5.981506, 3.398972, -0.5578156, 
    -10.98959, -0.1611938, -2.236969, -10.82318, -14.50754, -11.08383, 
    -5.242706, -8.294525, -7.735168, -8.969513, -8.375244, -8.619019, 
    -9.553894, -10.07397, -9.604431, -7.874481, -10.33258, -8.929169, 
    -7.653381, -11.04767, -8.81015, -2.714325, 3.074219, 6.208588, 7.623718, 
    5.289307, 0.5523682, -1.697647, 0.03019714, 3.772141, 5.656006, 7.6362, 
    0.0544281, -3.287231, -0.2807312, -2.218216, -9.084106, -8.153656, 
    -8.381241, -6.624741, -6.830734, -1.318481, 4.588547, 0.2484283, 
    -1.805206, -3.030991, -6.542969, -8.605743, 0.2533875, -2.834106, 
    4.394791, 5.538269, 0.1010437, 2.027328, -1.984375, -2.849976, 2.686188, 
    2.921616, 7.971863, 14.20338, 17.24661, 11.82761, 5.991119, 1.409363, 
    4.669281, 3.610168, 1.102875, 9.352341, 11.70157, 9.967712, 5.938278, 
    7.520309, 4.864334, -5.144775, -7.663528, -9.898697, -4.545822, 
    -3.243225, -9.75235, -8.083328, -7.431, -15.65573, -16.19246, -7.56459, 
    0.6455688, 5.3974, -0.7481995, 0.6174622, 10.75807,
  -3.870056, 2.103134, 0.9156189, -2.73204, -11.31927, -5.187225, -4.471603, 
    -4.239044, -3.276825, -1.857574, -5.12265, -9.163025, -9.639832, 
    -6.710938, -6.800262, -7.922913, -6.243225, -2.317474, -1.464325, 
    -1.314056, -6.351288, -8.230469, -6.980743, -13.23935, -7.705231, 
    -8.889603, -12.35884, -10.12579, -5.315887, -4.339066, -2.572418, 
    0.6148682, -4.507813, -7.418488, -10.22316, -3.079697, -5.039597, 
    7.045319, 4.567719, -2.296356, -10.38437, -11.28751, -5.130722, 
    -2.119278, -3.654953, 1.4599, 4.995575, 6.029694, 7.671875, 10.46771, 
    11.92188, 6.069, 3.41095, -1.860153, -1.863541, 0.5744781, -5.829941, 
    -5.050781, 2.949219, 1.0112, -5.839844, -6.718475, -0.2278595, 6.999222, 
    12.54948, 12.51042, 10.23412, 4.672119, 5.267426, 1.916931, -2.851044, 
    0.4914093, 6.847656, 4.663803, 7.094009, 9.504944, 7.964066, 11.75468, 
    19.86406, 15.97318, 8.359634, 8.415894, 1.56485, -6.953384, -4.996353, 
    -2.625259, -11.26744, -16.51509, -16.4724, -13.82135, -15.87943, 
    -10.32579, -0.1867218, -1.790375, -0.3494873, 2.119019,
  -3.923447, -7.879974, -14.31458, -8.506516, 0.4255219, -2.731247, 
    -1.609634, 3.715881, 2.581238, -0.6374969, 2.855972, 3.489075, -3.374481, 
    -3.219543, -3.559357, -3.273163, 2.606781, 1.207031, 3.071869, -2.183838, 
    -7.353912, -10.01901, -8.440613, -11.59479, -15.16251, -10.42369, 
    -8.989578, -12.87526, -15.37733, -16.08438, -12.66275, -13.25494, 
    -24.34843, -22.17499, -18.76563, -17.76459, -13.70416, -9.678375, 
    -12.45052, -12.5909, -11.77864, -16.00729, -17.39662, -11.96407, 
    -8.84375, -7.489594, -8.147919, -2.794785, 1.139069, 2.430466, 5.408081, 
    10.14349, 7.652878, 0.5919189, -6.173431, 0.05104065, 4.358597, 3.776031, 
    -0.407547, -9.227081, -9.601563, -5.272659, -8.150253, -9.138016, 
    -5.176559, 1.6362, 2.503387, -2.110687, 2.254684, -5.248184, -8.305466, 
    -5.953384, -7.996613, -7.949738, -1.765366, -26.83595, -2.903122, 
    -1.380203, -5.273178, -13.06667, -8.348953, -1.890884, -2.633072, 
    -10.44583, -16.13333, -11.71249, -5.293228, -7.889847, -12.16823, 
    -9.166656, -8.482025, -8.611191, -9.251572, -9.546616, -3.674225, 
    0.04428101,
  -0.09141541, -8.839584, -18.49297, -15.35001, -3.941666, -1.70285, 
    -3.32785, 1.079681, -2.281769, -1.370575, 2.523697, 5.761978, -0.7148438, 
    -1.041931, 0.5966187, 3.063538, 2.825516, 0.6575623, -2.70755, -2.983078, 
    -8.248688, -10.01875, -3.540359, -5.64035, -10.00574, -16.40312, 
    -19.69766, -14.15781, -19.49167, -24.25626, -25.96875, -18.58151, 
    -17.32292, -28.53802, -33.76094, -29.31017, -20.47577, -16.42891, 
    -18.30339, -23.85365, -32.86145, -32.09167, -23.34688, -11.24245, 
    -7.185684, -10.33984, -13.85834, -3.941925, 4.555725, 11.52057, 13.93672, 
    14.37135, 10.02213, 6.378647, 11.20052, 9.376556, 3.324478, -2.835419, 
    -9.429428, -17.50391, -21.95494, -20.35495, -15.64218, -9.254166, 
    -14.78229, -9.538025, -11.22864, -19.21484, -17.77682, -11.34818, 
    -10.90625, -17.26407, -37.63776, -38.64246, -34.57944, -30.82291, 
    -11.90208, -13.5789, -23.98671, -32.06406, -37.43567, -17.47057, 
    -11.28308, -13.60052, -14.40051, -3.356766, -0.7346344, -3.39949, 
    -2.574738, -6.345566, -8.629166, -5.430466, -2.255219, -10.89999, 
    -11.11172, -3.960419,
  -10.34349, -12.25494, -8.685928, -10.37604, -8.779175, -12.15312, 
    -2.905991, 2.659897, 1.178894, 4.052338, 5.733337, 0.4749908, -2.848969, 
    2.766922, 8.370041, 6.628647, 1.947144, 1.776291, 2.079941, -4.336456, 
    -9.722122, -10.34323, -8.818741, -10.29323, -13.01694, -18.02058, 
    -15.63933, -20.09949, -21.19113, -23.91563, -19.61015, -16.49948, 
    -12.53177, -12.16093, -17.25989, -22.54947, -19.91484, -23.92787, 
    -25.99767, -28.3362, -29.12787, -32.50339, -25.925, -16.65886, -12.01953, 
    -10.49661, -11.49687, -5.585419, 0.97995, 8.210419, 10.20988, 9.919266, 
    9.433334, 2.06485, -2.228394, -4.967453, -12.78775, -21.11224, -25.75911, 
    -20.56953, -20.22266, -18.18515, -13.97266, -5.142197, -9.603897, 
    -12.19688, -10.94843, -11.00781, -7.565109, -11.03671, -20.14244, 
    -33.81277, -36.9841, -29.57864, -24.35443, -27.60858, -24.97943, 
    -29.72423, -43.00676, -49.27266, -42.49609, -27.50079, -14.81276, 
    -6.06015, -6.603134, -5.279434, -6.258072, -5.971619, 0.1710968, 
    1.350266, -0.8760529, -2.814316, -4.476303, -9.293747, -7.447922, -6.0625,
  -12.42136, -12.4375, -3.990112, -2.882553, -7.498184, -2.499741, -5.482559, 
    2.890366, 7.4664, 6.734375, 1.277084, -2.381775, -1.472916, 3.505463, 
    6.804169, 2.445053, 0.2708282, -3.376831, -7.480988, -11.19948, 
    -8.106506, -5.305206, -5.004684, -8.206772, -13.17786, -17.53438, 
    -18.65547, -25.55806, -27.38203, -25.77812, -22.6823, -19.88438, 
    -16.74113, -15.2711, -16.08307, -18.4151, -24.85599, -28.72188, 
    -26.48932, -23.32265, -14.96016, -20.49609, -20.95782, -31.22084, 
    -36.27188, -32.10469, -20.20885, -14.8078, -14.95468, -1.552872, 
    -0.2450562, -16.29871, -5.55365, -0.4343719, -1.680466, -9.589584, 
    -15.56667, -16.31537, -14.87109, -21.26927, -28.02448, -35.08229, 
    -36.33932, -27.34843, -16.37421, -12.69765, -16.66197, -20.25261, 
    -19.86354, -20.69531, -26.38802, -29.02994, -26.49245, -25.0448, 
    -32.93697, -33.77214, -27.31329, -20.57187, -29.05417, -32.61302, 
    -45.88489, -30.68774, -14.17656, -4.353394, -0.153656, 1.184631, 
    3.677078, 6.655212, 7.766144, 4.457809, -3.655731, -2.885406, -0.7328186, 
    -0.8122406, -1.611206, -3.606262,
  -4.657288, -5.858078, -6.148956, -4.826294, -3.024475, 2.117706, 4.220566, 
    0.06692505, -6.09584, -6.666916, -6.751816, -6.869797, -8.389053, 
    -9.008591, -5.740112, -5.358597, -8.35025, -11.2198, -7.676559, 
    -4.763031, -0.05052185, -1.900772, -9.632813, -15.11069, -20.54636, 
    -28.98256, -27.30833, -23.05728, -17.35495, -16.82057, -15.85547, 
    -23.69817, -24.83203, -22.78384, -23.87187, -23.46484, -24.88568, 
    -34.40494, -33.28151, -27.96667, -23.16354, -23.04219, -29.17397, 
    -32.27553, -34.31537, -31.02864, -28.20781, -30.15886, -27.26068, 
    -19.88725, -21.17058, -30.35963, -32.20808, -17.21536, -13.65573, 
    -15.59193, -17.98671, -21.09532, -27.92474, -30.51485, -35.4888, 
    -35.59634, -34.22058, -30.58958, -27.54245, -25.59036, -21.29323, 
    -17.86224, -19.63515, -35.48543, -26.89635, -35.44714, -38.32266, 
    -38.80885, -25.67265, -25.52451, -19.45183, -22.48021, -30.01328, 
    -46.82916, -47.66458, -37.76276, -26.67163, -16.92004, -11.8638, 
    -9.006744, -4.954437, -0.640625, 2.517975, 2.103882, -14.27682, 
    -21.17343, -19.84792, -4.271606, 2.874741, 0.6695404,
  0.3752594, -0.2450562, 0.1835938, -0.2453156, -1.562241, 0.4309845, 
    2.603394, 1.721878, 2.573441, 3.17421, 1.539063, -7.1026, -22.37735, 
    -28.73985, -26.41068, -19.76172, -27.0383, -22.45259, -17.70468, 
    -12.2599, -15.52344, -13.58647, -15.70026, -16.44922, -19.07916, 
    -21.23802, -24.24115, -25.30495, -26.6638, -25.8065, -24.33568, 
    -25.04739, -24.78697, -26.20235, -24.90833, -23.80339, -27.10963, 
    -28.62944, -26.29713, -25.56798, -24.46173, -25.12135, -28.49036, 
    -32.14609, -35.40338, -35.92735, -33.75598, -30.12372, -27.67499, 
    -22.91614, -17.77681, -14.69061, -16.43672, -18.62709, -20.16145, 
    -20.44194, -18.96512, -19.84792, -20.82343, -23.00443, -25.11198, 
    -25.20546, -20.64818, -9.185684, -7.869278, -7.261719, -7.947128, 
    -7.227859, -10.73203, -22.60052, -22.38985, -25.18594, -27.15781, 
    -18.05989, -13.51797, -9.784897, -10.55339, -19.34116, -28.74011, 
    -34.11902, -31.20444, -26.80026, -20.04819, -19.72473, -17.51041, 
    -18.96823, -20.25, -14.58228, -7.433838, -1.933594, -2.552094, -12.41901, 
    -23.39011, -25.24037, -10.87057, -0.8192749,
  -3.575775, 3.019272, 2.685165, 0.9578247, -4.154694, -10.65103, -28.80782, 
    -36.12187, -35.49922, -26.38905, -24.88098, -23.74324, -24.40886, 
    -24.49998, -24.36928, -25.23828, -23.04063, -22.41902, -24.42267, 
    -28.18333, -28.87422, -27.46979, -24.65938, -21.46068, -21.19609, 
    -24.88255, -24.50052, -20.30208, -19.40729, -18.21068, -17.88046, 
    -11.33698, -8.881775, -7.163284, -8.382553, -9.960678, -13.19948, 
    -17.19922, -19.79688, -18.9086, -17.45755, -16.78725, -15.02814, 
    -15.29349, -18.69218, -23.52943, -25.8927, -27.74741, -29.28177, 
    -29.18437, -29.51511, -29.25026, -27.46353, -27.91145, -29.08099, 
    -29.43204, -29.54688, -27.24088, -22.03751, -16.9901, -11.32552, 
    -5.085403, -0.7648315, -1.603912, 0.5744934, 16.66484, 13.11121, 
    8.861984, 2.789597, -6.846619, -15.4716, -17.77812, -13.09975, -10.82449, 
    -12.09975, -17.23099, -19.11096, -22.49921, -23.21222, -24.61435, 
    -23.68854, -20.25418, -17.37994, -15.24323, -14.72498, -15.15701, 
    -15.80807, -16.36511, -16.48566, -14.45364, -10.60471, -15.28906, 
    -13.16721, -17.31485, -21.4091, -18.41615,
  -10.77943, -14.1539, -18.98386, -22.15286, -6.228119, -7.727859, -8.220825, 
    -18.91173, -15.78098, -13.41223, -13.9875, -15.58827, -18.27708, 
    -20.50807, -21.05339, -21.38905, -19.81615, -17.79558, -15.27318, 
    -14.08072, -13.80469, -12.52942, -11.78673, -10.29974, -7.963287, 
    0.9945221, -1.086197, -12.71379, -13.90808, -14.07761, -14.25626, 
    -13.23308, -12.5573, -12.19427, -12.60754, -12.70807, -12.00259, 
    -10.96275, -11.28595, -12.39088, -15.19792, -18.68906, -21.57214, 
    -24.43698, -26.46016, -27.70209, -27.29036, -25.93933, -23.18697, 
    -20.14662, -16.6763, -13.86876, -12.47632, -11.95522, -11.19194, 
    -10.85493, -11.91641, -13.42554, -13.2448, -13.5862, -12.2211, -11.48541, 
    -10.68593, -11.94531, -12.52917, -12.66667, -13.38672, -16.58386, 
    -18.33179, -19.05704, -17.69141, -17.18437, -15.85078, -6.577362, 
    -9.063782, -12.52213, -15.92941, -19.47034, -23.21716, -26.62891, 
    -27.71875, -28.33722, -26.45081, -22.26743, -16.81485, -11.13724, 
    -4.532806, 0.6471252, 2.202606, 2.217468, 0.9979248, -0.6200562, 
    -9.257294, -8.976288, -9.671875, -10.2052,
  -2.270309, -3.677078, -5.591141, -7.018234, -9.407822, -12.38124, -14.5448, 
    -15.91017, -17.92577, -20.77266, -23.53905, -25.57083, -27.26431, 
    -27.98698, -28.29167, -27.37553, -25.10858, -23.42371, -21.65962, 
    -19.78828, -18.22968, -18.17941, -16.48203, -15.63176, -15.87759, 
    -16.5638, -16.30312, -14.65651, -13.50026, -13.03046, -12.83542, 
    -12.52214, -11.95938, -10.50964, -8.783844, -6.496613, -4.89296, 
    -3.414841, -3.024734, -3.196091, -3.844009, -4.367447, -5.639053, 
    -7.329681, -9.314316, -11.04349, -12.2039, -11.84088, -11.64088, 
    -11.20183, -11.79376, -11.58853, -11.77942, -11.55885, -11.49452, 
    -11.49115, -11.67397, -11.80286, -12.75053, -13.23619, -12.13829, 
    -10.84035, -8.82579, -7.895569, -7.292191, -6.313019, -6.64296, 
    -7.029694, -7.991943, -9.128113, -9.829163, -10.15652, -10.43909, 
    -11.39194, -11.41171, -11.52759, -13.33435, -14.79895, -16.50992, 
    -18.31174, -20.26144, -20.98749, -20.18567, -18.12891, -15.26849, 
    -12.07343, -10.14294, -8.356232, -6.331787, -5.010925, -3.830719, 
    -3.714569, -2.100281, -0.7409058, -0.875, -1.363541,
  -8.231247, -8.003372, -8.20105, -8.642715, -8.996353, -9.39296, -10.14142, 
    -10.67006, -11.67578, -12.95131, -14.00104, -14.52943, -14.93333, 
    -15.50835, -16.06563, -16.20755, -16.42473, -15.7935, -15.61172, 
    -15.55391, -15.46771, -14.82838, -14.56015, -14.14088, -13.63646, 
    -13.47134, -12.66354, -11.49973, -10.45729, -9.452087, -8.715622, 
    -7.958344, -7.584366, -7.245834, -6.570313, -5.711975, -5.672913, 
    -5.809357, -5.788788, -5.603363, -5.720306, -5.54715, -5.599731, 
    -5.698975, -5.875275, -6.545593, -7.016144, -7.356232, -8.138794, 
    -9.234894, -10.40964, -11.45, -12.53491, -13.24818, -14.26848, -14.74507, 
    -14.93646, -14.94843, -14.76118, -14.10051, -13.4375, -12.91745, 
    -12.26953, -11.61667, -10.56041, -9.185944, -8.441406, -7.570313, 
    -6.383331, -5.735672, -5.369003, -4.826309, -4.817184, -4.862762, 
    -5.159378, -5.568481, -6.199219, -6.891922, -7.849213, -8.565872, 
    -9.13205, -10.52242, -11.0979, -11.61562, -11.95052, -11.99791, 
    -11.90808, -11.63905, -11.50546, -11.14792, -10.72475, -10.67084, 
    -10.1151, -9.812515, -9.266159, -8.814316,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.03697917, -0.04244791, -0.03333333, -0.03958334, -0.04010417, 
    -0.04401042, -0.03880209, -0.04375, -0.0408854, -0.03802083, -0.02604166, 
    -0.02473958, -0.01848958, -0.005208328, -0.006250009, -0.01822917, 
    -0.02395834, -0.01328126, -0.0002604127, 0.007291675, 0.01145834, 
    0.007031262, -0.00390625, -0.006249994, -0.0002604127, 0.001041666, 
    -0.008593753, -0.01927084, -0.02109374, -0.02838542, -0.03749999, 
    -0.028125, -0.03151041, -0.0203125, -0.01406249, -0.01666666, 
    -0.02395834, -0.02135417, -0.01145834, -0.01380208, -0.02005209, 
    -0.02760416, -0.0296875, -0.04479166, -0.06354167, -0.05390626, 
    -0.0421875, -0.03255208, -0.02760416, -0.02942708, -0.03697917, 
    -0.03776042, -0.03802083, -0.04192708, -0.04166667, -0.04531249, 
    -0.03671874, -0.02786458, -0.03072917, -0.03203125, -0.02473958, 
    -0.02890626, -0.02890624, -0.02838542, -0.03645834, -0.03802083, 
    -0.04713541, -0.04817709, -0.02994791, -0.01666667, -0.0078125, 
    -0.005468756, -0.01640625, -0.02578124, -0.02838542, -0.03098957, 
    -0.02369791, -0.01901041, -0.01796875, -0.009114586, -0.01041666, 
    -0.01223958, -0.00390625, -0.00338541, -0.00390625, 0.002864584, 
    -0.005729169, -0.0005208403, -0.001302078, -0.002343744, -0.006510422, 
    -0.005729169, -0.01041666, -0.002083331, -0.0078125, -0.02942708,
  -0.3367187, -0.3973958, -0.3583333, -0.3182293, -0.3710936, -0.4135417, 
    -0.3015625, -0.2684897, -0.2802083, -0.2822917, -0.2437501, -0.2351563, 
    -0.1346353, -0.1049478, -0.1335938, -0.1289063, -0.1291666, -0.190625, 
    -0.2281251, -0.2601564, -0.213021, -0.08125019, -0.0640626, -0.08333325, 
    -0.001562595, -0.0184896, -0.1182294, -0.1786458, -0.1916668, -0.2520833, 
    -0.2760417, -0.2210939, -0.09401035, -0.0859375, -0.0872395, -0.03046882, 
    -0.0263021, -0.0320313, -0.04869795, -0.1033854, -0.1380209, -0.1065104, 
    -0.1083333, -0.1755208, -0.2549479, -0.2731771, -0.3098958, -0.328125, 
    -0.3333334, -0.2583333, -0.2130209, -0.1546875, -0.0604167, -0.1484375, 
    -0.2195313, -0.1872395, -0.2002604, -0.3109375, -0.2611979, -0.2739583, 
    -0.18125, -0.008854151, -0.04505205, -0.2830728, -0.4440104, -0.5640625, 
    -0.508073, -0.4786459, -0.3330729, -0.3028646, -0.3710938, -0.4208333, 
    -0.3578125, -0.3447917, -0.3544271, -0.353125, -0.2325521, -0.0994792, 
    -0.0567708, -0.1195314, -0.1276041, -0.1257812, -0.05989587, -0.0234375, 
    -0.002343774, -0.05729175, -0.1838541, -0.2239584, -0.2434895, 
    -0.2046875, -0.2757813, -0.2705729, -0.2302084, -0.2354167, -0.2471355, 
    -0.3385417,
  -0.7747393, -1.079167, -1.429948, -1.426042, -1.217448, -1.034896, 
    -0.8968754, -0.8041668, -0.8757815, -1.193229, -1.610937, -1.464323, 
    -1.039583, -0.7875004, -0.678906, -0.6817708, -0.6317711, -0.6351562, 
    -0.6937499, -0.6713538, -0.5921874, -0.3226562, -0.1820312, -0.6643229, 
    -0.6065106, -0.5679688, -0.5083332, -0.3062501, -0.5101562, -0.4880209, 
    -0.2911458, -0.4273438, -0.2145834, 0.0838542, 0.4653645, 0.4781251, 
    0.009114265, -0.1739583, -0.7249999, -0.8499999, -0.5882812, -0.6213541, 
    -0.5367188, -0.3960938, -0.2627606, -0.2929688, -0.2971358, -0.2609372, 
    -0.1888018, -0.1374998, -0.0718751, -0.1526041, 0.04739571, -0.1695309, 
    -0.1372395, -0.002864361, 0.229948, 0.3096356, 0.04453135, -0.116406, 
    -0.2567706, -0.3161459, -0.106771, -0.1354165, -0.2432294, -0.5348959, 
    -0.492969, -0.2703123, -0.2302084, -0.1265626, -0.2776041, -0.2093754, 
    -0.15625, -0.2914062, -0.3971357, -0.3752604, -0.3966146, -0.06744814, 
    -0.02630186, -0.5044274, -0.6776042, -0.6710935, -0.5018229, -0.488802, 
    -0.5828128, -0.6888022, -0.7648439, -0.703125, -0.7791667, -0.7739582, 
    -1.006771, -1.333333, -1.052865, -0.5471354, -0.6598959, -0.8361979,
  -2.641147, -1.94427, -1.98724, -2.0375, -2.048438, -2.272917, -2.014063, 
    -1.090885, -0.7752609, -0.9651041, -0.7039061, -0.6536455, -0.915885, 
    -1.138021, -0.8822908, -1.063021, -1.529687, -1.621354, -1.520312, 
    -1.747656, -1.758594, -2.008333, -1.690886, -0.848177, -0.573698, 
    -0.7950516, -0.9919271, -0.6783857, -0.97474, -1.042969, -0.5674486, 
    -0.3205738, -0.4065104, -0.5789061, 0.03151035, 0.3466139, 0.2179689, 
    -0.06588554, -0.4546871, -0.535677, -0.08072948, 0.2921877, -0.04635429, 
    -0.1419268, -0.08307266, -0.2442713, -1.078385, -1.311979, -0.6783848, 
    -0.0114584, -0.5684891, -0.5541668, 0.3309898, 0.1002598, -0.6656246, 
    -0.4265623, 0.003385544, -0.2489586, -0.2156248, -0.05911446, -0.124218, 
    -0.4648438, -0.761198, -0.317709, 0.05208302, -0.2070313, -0.198698, 
    0.1622391, 0.2476568, -0.6395836, -1.000781, -0.53125, -0.6882811, 
    -1.01875, -0.6031256, -0.4015627, -0.01770878, -0.01536465, -0.06822968, 
    -0.4255209, -1.028646, -0.604167, -0.807291, -1.144271, -1.197135, 
    -1.473958, -1.828906, -2.117708, -2.333854, -1.733073, -1.556251, 
    -2.124219, -2.144271, -2.150261, -2.410677, -2.749219,
  -1.555729, -0.96875, -2.105207, -1.939585, -0.9617176, -0.9460926, 
    -0.8953133, -0.1596355, 1.252344, 0.7906246, 0.6533852, 0.1463547, 
    -0.07187653, 0.4388027, 1.040363, 0.2885418, -0.2789059, -0.2250004, 
    -0.4273434, -0.8843746, -0.6289063, -0.5276051, 0.1924496, 1.333334, 
    0.5539074, -0.2791653, -0.4481773, 0.7661457, 0.3132801, -0.5033855, 
    0.0627594, 0.7846355, 0.4880199, -0.104948, -0.1643238, -0.6460934, 
    -0.6619797, -0.697916, -0.9713554, -0.495573, 0.04479027, 0.9494801, 
    0.1901054, -1.539583, -1.09948, -0.3976555, -1.139845, -1.578646, 
    0.5830727, 2.137239, 0.4468765, -0.7289047, 0.2885418, 0.5382805, 
    0.4463539, 1.173698, 1.812239, 2.160936, 1.419271, 1.649479, 1.39271, 
    -0.02968788, -0.4007816, -0.4044266, 0.05729103, -0.2255211, -0.4911442, 
    0.3109379, -0.1757813, -1.023176, -0.6950512, -0.03333282, -0.5078125, 
    -1.134897, -1.295834, -1.038542, -0.452343, -0.3247395, -0.7307281, 
    -0.3716145, -0.2312489, -0.3354168, 0.06588364, 0.2015629, 0.104166, 
    -0.1489582, -0.2992191, -0.2630215, -0.1750011, -0.6885414, -1.074739, 
    -0.892189, -0.4192715, 0.229166, -1.027864, -2.128906,
  0.2963543, -0.7218761, -0.4445305, 1.326822, 1.532553, 0.06822968, 
    0.2437496, 1.394009, 1.447136, 0.7380199, -0.547657, -0.6304684, 
    -1.747135, -2.010939, -0.5656261, -0.864584, -1.128906, -1.053905, 
    -0.08567619, -0.895834, -0.4398441, 0.8182297, -0.04140663, -0.1416664, 
    0.8809891, 1.060156, 0.3411465, 0.4255199, 0.9953136, 0.3507824, 
    -0.2721348, -0.5151043, 0.08724022, -0.8252621, -0.8945313, -1.576563, 
    -0.5127621, -0.3179703, -0.4513016, -0.96875, -0.04192734, 0.3825512, 
    1.216928, -0.704689, -1.373438, -0.6174469, 0.8619804, -0.8427086, 
    -1.056509, -0.1666679, -0.4500008, 0.2101555, -0.7315102, -0.01093674, 
    0.9911461, 1.988541, 1.425522, 1.051043, 2.030209, 2.172655, 1.124218, 
    0.2424488, 2.105991, 0.2169266, 0.02395821, 1.185417, 1.28125, 0.2645836, 
    -0.8007813, -0.9765625, -0.2666664, -1.208855, -1.652605, -0.1575508, 
    0.5127602, -1.679167, -1.548698, -0.8604164, -0.7109375, -0.05833054, 
    1.727863, 1.77552, 1.035934, 2.064062, 0.6843758, -0.3028641, 
    -0.05078125, 0.7726555, 0.9807281, 0.7809887, 1.277082, 1.065365, 
    -0.1197929, -0.8018227, -1.008854, -0.5934906,
  0.5635414, 0.2208328, -1.152863, 1.254948, -0.8390617, -1.989323, 
    -0.7414055, -1.335674, -2.297134, -2.804428, -3.46146, -2.27578, 
    -1.790363, -3.135414, -2.161457, -1.646877, -0.9213562, -0.5523415, 
    -1.74453, -1.524738, 0.7156219, -0.5729141, -1.121876, -0.717968, 
    0.8466148, 2.22578, 0.8356743, -0.7815132, 0.1458321, 0.7197914, 
    1.203907, 1.104168, 0.5375023, -0.3026047, -0.9562492, -0.4036484, 
    2.929947, 1.073959, 0.6145859, -0.0471344, -2.174999, -1.914845, 
    1.076565, 1.098698, -1.891148, -0.1968727, 0.842186, 0.6875, 0.2262993, 
    -0.4369774, 0.4476585, 1.01432, -2.382294, -2.493752, -0.4223976, 
    0.421875, 0.5065117, 0.8752594, 3.277344, 2.03854, 2.029949, 2.871876, 
    1.41901, -0.1520844, 1.271873, 0.6151047, -0.157032, 0.186718, 
    -0.1768227, 0.08463669, -0.3031235, -0.4177055, -0.9424477, 0.3809891, 
    -0.2755203, -2.724998, -2.407553, -1.771093, -0.7703094, -0.2455711, 
    1.521355, 1.213543, 0.3997383, 0.7369804, 1.907814, 1.365364, 0.7299461, 
    1.171093, 0.2966118, 0.6203117, 1.277863, 2.472397, 2.352341, 0.515625, 
    0.7765656, 0.2315102,
  -0.09531403, -0.9302101, -2.481251, -1.146873, -0.1770821, -1.50573, 
    -3.288021, -3.511459, -2.045055, 0.7098961, -0.4221382, -1.590885, 
    -1.850517, 0.0544281, 0.2164078, -0.6716118, -0.2992172, -0.5299454, 
    -1.651302, -0.5822906, -0.1377602, -1.938541, -0.7192726, 2.30521, 
    2.39167, 3.184113, 5.025002, 4.765106, 1.81094, 2.147919, 3.898956, 
    4.386459, 0.9033852, 1.60651, 3.143486, 0.2072945, 0.828125, 1.485939, 
    0.7184906, -0.3244781, -2.202343, -2.880989, -0.04322815, 0.985157, 
    0.6244812, -0.7791672, -0.2559891, 0.9580727, 2.974998, 3.058334, 
    1.164063, 0.6854172, -0.4979134, 2.066406, -0.9466133, -0.264843, 
    1.916409, 1.508331, 0.3502617, 0.4937477, 0.6338539, 1.930992, 1.058594, 
    0.7091141, 2.336716, 0.9653625, -1.546616, 0.9346352, 2.647396, 1.151825, 
    0.25, 0.8669281, -1.729946, -2.992966, -0.2861977, -1.369274, 
    -0.07526398, -1.334373, -0.5880203, 1.333069, 1.615364, -0.2458344, 
    -1.787498, -0.4713516, -0.4223976, -0.2908859, 0.6455727, 1.195572, 
    -0.5703125, 1.326565, 1.671093, 1.776043, 1.380207, 0.4666672, 0.8901024, 
    0.2526016,
  1.276299, -0.5255203, -2.047394, 1.821358, 2.311981, -2.830467, -4.02813, 
    -3.0849, 0.27005, -1.689323, -3.082031, 3.447395, 5.923958, 5.019012, 
    4.683334, 3.454948, 1.802864, 4.190887, 2.417709, 1.648178, 2.570313, 
    4.299995, 8.464325, 8.338806, 5.594009, 3.844788, 4.809891, 4.08567, 
    2.651825, 2.346611, 3.655731, 5.509636, 2.268745, 2.060936, 3.494011, 
    2.855469, 0.5713501, -1.07214, 1.025002, -1.331512, 1.133591, 1.245575, 
    -0.3604126, 1.701042, 2.054428, -0.422142, 1.052345, 3.616146, 5.408592, 
    2.433598, 3.431252, 4.091408, 1.153908, 2.909637, -0.8565063, 0.7937546, 
    2.13047, -0.5112, 0.2674484, 0.672142, 0.7072906, 1.629951, 0.7653656, 
    0.1127625, 0.2697906, -1.432293, -1.574478, -2.540367, -2.675522, 
    -2.098175, -0.5270844, -0.6557274, -1.44297, -0.171608, 0.4794312, 
    2.660416, 3.399483, 0.6804695, -0.8515625, 0.155983, -0.5812531, 
    -0.1257858, -1.678902, -2.615891, -3.416664, -3.875519, -2.496094, 
    -2.069267, -4.01432, -3.022919, -0.3015594, 0.6721344, -0.9929657, 
    -2.003639, 1.609116, 0.8049469,
  1.100006, 3.533333, 6.173958, 2.550255, -0.0158844, 0.9742203, 3.293747, 
    4.137505, 3.436195, 4.929169, 8.522133, 15.09141, 14.05235, 10.38906, 
    9.544792, 8.436203, 8.1987, 6.227867, 7.888535, 11.00755, 10.05807, 
    9.878647, 9.104164, 3.984901, 0.9179688, 4.054161, 3.63047, -1.299484, 
    1.718224, 1.487762, 3.479942, 1.455475, 3.998177, 3.32135, 0.9041672, 
    -1.585159, 0.5539017, 1.004684, -0.9268188, 0.8695297, 2.36042, 
    0.3070374, -6.74453, -2.026825, 0.9679718, 0.05364227, 1.360153, 
    4.050781, 2.264061, 6.012756, 7.051048, 4.831253, -0.6200485, 0.4263, 
    0.7255173, -1.567192, -0.1549454, 0.1804733, 3.307808, 1.702599, 
    2.060936, 2.400002, 0.3143234, 0.3799515, 0.7307281, -2.346619, 
    -3.767448, -2.098701, -0.01822662, 1.288803, 0.6958389, 1.888023, 
    0.171875, 3.915627, -0.0942688, -0.3572922, 1.81797, 0.6187515, 
    -2.927345, -1.651299, 0.862236, -1.113022, -5.461197, -3.351044, 
    -0.5354156, -0.8255157, -0.9598923, 0.127861, 2.541672, 3.836464, 
    1.772659, 1.234894, 2.024483, 4.186455, 2.779945, 1.859894,
  3.773438, 3.866661, 3.624481, 1.882545, 1.590881, 3.595314, 6.484375, 
    3.472397, 3.713799, 3.975266, 11.75521, 7.087761, 7.373695, 12.2401, 
    11.20287, 7.720314, 8.415359, 6.623962, 5.615883, 5.926308, 5.004433, 
    -0.2976532, -0.4075546, 1.818489, -2.037506, 0.1479187, 1.127083, 
    -3.176819, -1.324478, 1.099739, 4.805733, 0.1773376, -4.684639, 
    -2.331253, -5.086723, -6.427086, -4.415108, -2.914841, -5.358856, 
    -4.082291, -2.492455, -2.950005, -2.343491, 0.7518234, 2.62735, 3.704948, 
    5.064583, 6.2612, 5.879692, 3.684113, 5.209114, 2.383072, -0.3247375, 
    -0.2612, -2.107292, -1.944794, -1.021355, 1.836716, -1.554169, 0.1476593, 
    2.8125, 1.523438, -3.891403, -2.591141, -2.285156, -6.669533, -4.9375, 
    -6.329689, -2.467194, -0.8723984, 0.1520844, 2.3862, -1.901825, 
    -2.143227, 0.159111, 1.673965, 0.4487, 0.6856766, -3.01355, -3.706772, 
    -2.385162, -4.196869, -3.933594, -1.759636, 5.774734, 4.448959, 5.147133, 
    4.706512, 2.249481, 0.6039047, 2.730469, 2.981514, 3.086716, 3.087761, 
    2.066666, 0.3559875,
  1.504173, 1.514069, 1.037247, -0.05130005, 2.498962, 5.385147, 10.51146, 
    14.1823, 5.898697, 3.275772, 6.995567, 6.92865, 5.839844, 10.73933, 
    7.075783, 5.045837, 8.794014, 10.82943, 6.543228, 0.9679718, 1.99115, 
    0.1992188, 1.284897, 4.737762, 1.085678, -1.670311, 0.778389, -3.736717, 
    -6.710159, -1.840881, 3.576569, -1.038803, -7.189056, -9.555984, 
    -4.453384, -2.501038, -9.367195, -7.352859, -7.28125, -10.23567, 
    -10.62943, -1.801826, 7.017189, 6.172653, 8.706512, 4.369789, 2.85807, 
    1.66172, 3.811714, 4.120049, 0.06771088, 3.754684, 3.111458, 3.902863, 
    3.632286, 2.33828, 2.4263, -0.0776062, -4.490097, -1.734901, -3.867966, 
    -5.494537, -5.402603, -6.016411, -2.158073, -3.741661, -4.113281, 
    -6.141144, -1.566406, -4.77578, -1.872139, -1.307289, -2.118744, 7.46328, 
    3.309906, -0.954422, -3.303131, -4.080475, -5.099747, -1.873169, 
    6.065628, 6.825523, 7.075783, 4.578651, 4.779694, 2.862244, 5.109642, 
    4.900787, 2.174217, 2.060677, 3.98307, 2.859901, 1.870834, 2.176308, 
    2.256508, 3.239067,
  0.6809998, 1.017181, -2.507813, 0.348175, 0.9171906, 7.004425, 10.07266, 
    10.47501, 7.326569, 5.560944, 8.079178, 4.967712, 2.908066, 1.451035, 
    3.216156, 7.520309, 5.162506, 5.066406, 5.527344, 5.973953, 1.632034, 
    2.790627, 0.1583328, 0.8828125, 0.703125, -1.938278, -3.143219, 
    -5.253906, -4.290359, 0.3252563, 5.047928, 3.058334, 0.146347, -4.394791, 
    -5.944519, -13.23177, -17.96719, -8.073959, -8.334641, -8.491669, 
    -5.184898, 1.859116, 6.483597, 1.244263, -1.486206, -1.423965, 0.9039001, 
    3.192703, 6.529678, 5.607025, 4.160156, 4.0737, 6.215622, 3.259109, 
    3.517448, 2.635681, -3.392448, -3.044014, -2.098434, -8.135681, 
    -8.842186, -9.077866, -6.667969, -4.875519, -7.729416, -5.178909, 
    -5.822128, -5.730988, -4.119537, -5.635422, -3.998184, -4.214066, 
    0.4552002, -2.764069, 1.301559, 1.543488, -5.551315, -7.585938, 
    -4.539581, 0.1929779, 10.76067, 8.768234, 6.165115, 14.12813, 6.513802, 
    0.1695251, 2.807556, 0.958847, -2.264328, -2.507813, -2.237762, 
    -1.148438, -2.21537, -1.783066, 0.6526031, -0.4148407,
  -1.606506, 2.240891, 0.6901093, -1.597656, -1.035675, 6.672394, 8.417191, 
    5.288544, 5.483582, 0.3346252, 0.2166595, -2.410156, 4.293747, 10.35208, 
    -1.108063, 4.873962, 6.54454, 3.882813, 7.8237, 5.820053, 0.6539154, 
    0.04348755, -0.4804688, -0.8153534, -2.802872, -3.58725, -2.351563, 
    -3.744019, -2.070572, -0.8513031, 4.204178, -0.1533966, -4.272141, 
    -5.995834, -10.14244, -10.87735, -9.905991, -7.526566, -6.000519, 
    -4.496353, -2.551559, 1.438278, 0.2921906, -3.750519, -2.166931, 
    -0.5575562, 4.2453, 6.567703, 1.615372, 0.2638092, 3.285156, 4.198441, 
    4.382553, 2.007294, -5.564056, -3.349747, -4.213287, -2.027863, 
    -4.717697, -4.590622, -3.186707, -5.702606, -5.284119, -4.416916, 
    -1.610168, -3.671616, -2.142441, -0.879425, -2.276306, 1.101044, 
    0.7635345, 1.162247, -3.772141, 2.853119, 3.6474, -8.586716, -5.903381, 
    -6.21875, -1.645828, 8.48671, 11.55939, 6.482025, 5.493484, 12.46172, 
    10.22707, 3.702858, -2.947403, -4.248962, -2.4263, -1.512772, -4.739578, 
    -4.227097, -3.836716, -1.697403, 0.4804688, -0.9656219,
  4.630981, 8.500778, 1.577347, -2.902344, -2.216415, 4.703125, 0.141922, 
    0.7736969, 5.773697, -0.1635437, 1.916153, -6.667435, -3.828384, 
    0.7666779, -0.9976501, 4.048431, 6.470047, 3.616409, 2.358322, 2.390106, 
    1.084122, -1.903656, 0.4570313, -1.66954, -3.495834, 0.8559875, 1.592697, 
    1.594269, 5.733337, 6.670319, 3.260941, -2.958862, -7.498169, -5.983063, 
    -6.018753, -6.286713, -2.886978, -2.639847, 2.368759, 5.533844, 
    0.7208252, 1.064575, 0.4450531, -1.120575, 3.385406, 3.831253, 5.246094, 
    4.230469, 5.818237, 2.480469, 3.867722, 3.513809, 4.183594, 3.82579, 
    3.2211, 1.059891, -3.384888, -1.866135, 0.3721466, 2.847656, -3.566147, 
    1.694778, 5.147919, 2.627869, 5.044022, 5.333588, 2.232803, 0.8986969, 
    0.2898407, 5.579163, 0.2562561, 0.3940125, 3.278137, 5.493484, -9.651306, 
    -6.302612, -4.969269, -4.491669, 6.31015, 16.83359, 6.85495, 8.764832, 
    7.5047, 8.214584, 18.47188, 10.45052, -3.455994, -6.813278, -8.485672, 
    -4.847137, -9.609894, -4.862244, -6.635681, 0.8627625, -0.6471405, 1.00209,
  7.540359, 5.7724, 5.214325, -3.194794, -2.81015, 2.730988, -2.021881, 
    -0.9880066, 5.599731, -0.8197784, 7.810944, 0.4617157, -4.183853, 
    0.1690216, 0.53125, 0.578125, -1.828125, -1.875, -1.973434, 1.045319, 
    2.038284, 5.259384, 2.51355, -0.7934875, 2.726303, 4.265106, 7.390884, 
    5.070053, 3.779953, 2.900513, 4.620834, 3.329681, 1.108597, -3.373184, 
    -5.33905, -4.393494, 7.959381, -1.897919, 2.15625, 6.053116, 0.1669312, 
    -0.2640686, 0.1854248, -1.589844, 3.301315, 1.500778, 6.622406, 4.902863, 
    3.025269, 3.560928, 1.267456, 2.142456, 1.462234, -0.6156158, 1.012772, 
    -0.4536438, 2.733856, 3.482544, 5.054428, 4.463013, 2.909897, 1.692459, 
    4.379425, 2.025528, 5.392975, 6.495575, 2.888275, 6.121094, 3.363541, 
    3.792191, 4.858597, 11.90129, 8.311722, -1.592712, -6.062759, -4.622391, 
    -1.329681, 1.470825, 12.24115, 11.18437, 6.855988, 2.655472, 14.59608, 
    7.111191, 15.13959, 11.24921, -4.245819, -7.014847, -3.805206, -2.52005, 
    -3.560684, 5.208069, 5.314072, 7.586975, 2.352341, 9.322647,
  9.577347, 10.91536, 0.8520813, -10.23723, -3.306503, -2.721359, -3.4375, 
    -2.971085, 0.4708252, -6.254944, -1.683594, 0.3127747, 3.255997, 
    3.106247, -2.054947, 3.083084, 5.158844, 1.230728, 1.3302, 2.649994, 
    2.25235, 3.399216, 0.5614624, -0.971344, 2.012238, 1.192703, -1.320572, 
    -3.746872, 0.1429596, -1.423447, 0.6622314, 5.495834, 3.025253, 2.880737, 
    -0.01329041, -3.546616, -7.42421, -10.96797, -5.810928, -0.1536407, 
    -2.442444, -4.756516, -4.989059, 0.1356812, 2.023697, 5.119537, 5.679428, 
    3.868225, 2.264847, 2.702347, 1.219528, 3.335144, 4.314056, 0.8497314, 
    2.017715, 2.198685, 3.384109, 1.843231, 5.001312, 3.085938, 4.510925, 
    3.468491, 6.616394, 6.381241, 7.336197, 5.2388, 6.907303, 6.881775, 
    7.366928, 7.654175, 8.116135, 5.355728, 6.319016, 0.1398315, -3.337769, 
    -3.257034, 1.335419, 2.816666, -0.4356842, 4.397385, 2.211197, 2.802078, 
    14.00131, 4.349228, -3.083069, 4.540359, 3.020309, -7.182541, -4.595062, 
    -2.742188, 0.8463593, 2.56485, 1.645569, 1.885941, 4.3461, 11.74193,
  4.435684, -0.8002625, -7.406509, -1.435684, -5.046631, -2.8638, -4.423981, 
    -4.111725, -4.17395, -9.145844, -2.259369, 15.41641, 4.53125, 2.786194, 
    2.249481, 4.7388, 3.101822, 3.869278, 3.800262, 2.636978, 3.771866, 
    5.030212, 2.489319, 2.322647, 2.341141, 3.365875, -0.0846405, -7.210938, 
    4.209122, 2.144272, -1.885162, -0.0942688, -0.4898529, 1.746613, 
    3.271622, 1.833603, -17.44922, -28.79739, -9.209106, -2.875793, 
    -0.4020844, -2.71199, -3.680206, -2.392975, 0.6593781, 1.993759, 
    6.382553, 4.284378, 3.4263, 4.834122, 6.083328, 8.806503, 10.02734, 
    7.111206, 6.157028, 6.536469, 4.228653, 2.791672, 2.982025, 1.268494, 
    4.237244, 5.274994, 9.284119, 6.761719, 9.7612, 8.689316, 11.19974, 
    10.93178, 9.322128, 4.795578, 8.887512, 6.389587, 3.302338, 0.1028595, 
    -8.003906, -6.550522, 0.6184845, 0.05183411, -0.9450531, -0.5018158, 
    -0.2408905, 5.251831, -0.646347, 0.05259705, -5.932816, -7.272919, 
    3.879425, 0.2473907, -1.72995, -4.156769, 1.068497, 2.369019, 5.045578, 
    4.147919, 5.01796, 8.150528,
  4.074738, 4.511459, 1.456757, 1.839844, -12.34064, -9.441406, -6.402359, 
    -9.292709, -13.36848, -11.17578, -12.63983, 15.25183, 12.01224, 4.68074, 
    2.738022, -0.4833374, 4.535156, 5.578918, 3.65416, 2.158585, -0.2778625, 
    -3.961456, -3.400269, -3.908066, -3.250259, -0.0161438, -2.004944, 
    1.577087, 1.592712, -3.246353, -4.773438, -8.610947, 5.66745, -7.957291, 
    -7.89505, 3.364319, -2.517975, -16.09089, -10.32655, -6.867447, 
    -7.738281, -3.050781, -4.995575, -9.500519, -10.28412, -9.971878, 
    -12.78073, -18.2263, -20.76225, -18.7198, -22.994, -22.93176, -16.22292, 
    -14.54765, -10.57838, -7.845566, -5.317184, -1.545837, 0.1510468, 
    3.133057, 4.240356, 6.735168, 9.072144, 7.148682, 7.870041, 7.373703, 
    5.671616, 4.215103, 1.875534, 2.078384, 2.809372, 3.233597, -1.356766, 
    -3.219269, -14.95886, -9.103638, 6.681503, 15.85573, -1.022659, 1.9422, 
    4.831512, 3.649231, 1.481781, 5.706238, -1.451828, -1.698944, -1.377609, 
    -3.396103, -9.407028, -9.784622, -4.890625, -4.445572, -2.35495, 
    0.7132721, 3.511719, -1.477081,
  2.396088, -3.287766, -0.1531219, -0.467453, -10.29115, -11.17578, 
    -0.6843719, -0.2268219, 0.9755249, -10.60495, -10.1875, -0.9125061, 
    10.32135, 1.421112, 4.410156, 5.056519, 7.644272, 2.546616, 1.299988, 
    -0.8773651, -2.028641, -3.479156, -4.124222, -7.392441, -5.858063, 
    -3.427353, -6.249237, -8.742706, -9.302094, -7.048706, -0.5830841, 
    -24.78828, -26.04897, -16.95338, -12.7112, -5.803391, -5.114075, 
    -9.414322, -7.684631, -8.9599, -6.573181, -5.045837, -15.56432, 
    -20.72499, -17.84792, -15.02708, -14.1362, -13.04271, -7.957809, 
    -8.938019, -14.09583, -16.87605, -16.40234, -16.33568, -13.16537, 
    -8.980225, -10.52994, -6.486176, -5.098694, -2.893494, 0.7416687, 
    -1.503906, 0.1393127, 3.639069, 2.35495, 1.827362, 1.313538, -2.564316, 
    -1.370575, 0.451828, -6.152084, -6.360687, -11.47917, -13.51746, 
    -21.43437, -14.05702, 5.102859, 0.3132782, -0.9322968, 13.82448, 
    6.087234, 11.1375, 18.08177, 6.240631, 5.175247, 13.1138, 14.08698, 
    12.02501, 3.106766, 4.767181, -2.132278, -0.7025909, 1.279678, 2.490356, 
    1.7677, 1.596359,
  4.022141, -4.588547, 2.067444, 4.5336, -0.6984406, -2.640366, 2.853119, 
    6.11824, 19.12604, 8.887497, -12.43203, -2.773178, 0.9044189, 1.547119, 
    3.955719, 1.870331, 0.9031219, 5.681259, 6.951828, 0.2054749, -3.596878, 
    -9.427078, -12.34686, -9.922928, -5.637238, -2.361176, 1.366135, 
    -12.2328, -3.554947, 3.984116, 3.420044, -2.28125, -9.329956, -6.126556, 
    -0.477356, 0.8486938, 0.3187561, -4.157288, -3.32579, -6.940369, 
    -3.892715, -6.458328, -3.630737, -6.006775, -3.785675, -9.047653, 
    -2.409637, 3.946609, 4.838287, 3.764847, 2.719528, 0.5848999, -1.343231, 
    -0.4466248, -2.132294, -3.507553, -4.795303, -7.241928, -8.322388, 
    -13.5625, -4.105988, -4.277863, -6.515625, 1.377869, -1.819, -4.53801, 
    -10.8461, -2.746353, -2.361984, -5.458603, -9.766663, -7.775513, 
    -13.66145, -15.22266, -12.37917, -3.810158, -13.91536, -8.431763, 
    17.70522, 29.21275, 10.67917, 7.852341, 1.86145, 2.277603, 6.175262, 
    10.9987, 14.01823, 7.343491, 9.711456, 9.6698, -2.460938, -2.173447, 
    1.001831, -5.306519, 5.110687, 10.25677,
  9.065613, 16.96642, 7.748428, 12.55782, 8.966919, 5.758591, 3.202347, 
    6.670319, 16.18333, 25.29765, 7.537247, 0.8999939, -5.169281, -6.611725, 
    -4.487488, -9.168762, -6.074493, -4.232819, -1.697388, -4.532288, 
    -6.674728, -9.294266, -23.04245, -17.77396, -2.855469, 3.242188, 
    0.1893158, 2.538803, 9.318237, 12.55156, 7.486206, 3.597137, 7.216141, 
    3.998962, 7.298431, 8.094269, 5.476303, 3.428375, -1.680481, -1.528656, 
    -0.9380188, 1.53125, 1.938278, 1.376831, 4.646103, -5.738541, -0.8953094, 
    1.050522, -2.801834, -1.287491, -0.3213501, -0.8416595, 0.6828156, 
    3.754166, 3.650009, 1.982819, 3.677597, 3.629944, 2.862762, -4.973709, 
    -3.470306, 4.326294, 12.64375, 12.65025, 14.30104, 11.89844, 13.89375, 
    25.00938, 22.59818, 16.3474, 8.693237, 5.220047, 7.239319, 3.602081, 
    5.877075, 7.324219, 12.50365, 32.2776, 25.01353, 5.751038, 1.092987, 
    4.052856, -2.0737, 2.6073, 1.236984, 5.7388, 5.927078, 0.2770844, 
    1.590363, 4.053116, 7.966919, 4.150269, 8.574997, 17.30495, 20.89011, 
    22.30728,
  9.012756, 8.140106, 0.6557159, -1.471619, -1.508881, -4.076553, 3.031006, 
    7.45314, 14.21771, 23.39558, 20.54817, -1.992432, -2.012482, -6.091675, 
    -5.889832, -6.252838, -10.85156, -9.859375, -11.30026, -12.78725, 
    5.191406, -12.13983, -24.05078, -19.58568, 2.425262, 8.967712, 17.36302, 
    29.79453, 16.82318, 1.863281, 1.401825, 3.431519, 11.37187, 3.40416, 
    5.396103, 4.8302, 2.253647, 1.724731, 3.3349, 0.998703, -4.219009, 
    -7.322403, -3.692978, -5.882553, -3.691666, -1.462234, -3.181259, 
    0.2247314, 0.7494812, -2.183075, -1.522644, -2.454437, 0.1197815, 
    1.649506, 0.5413971, 1.08931, 2.863556, 6.880997, 6.126038, 9.172928, 
    7.769257, 9.537491, 6.835419, 6.648422, 16.45494, 17.49504, 23.06224, 
    33.66484, 31.0453, 24.2578, 17.76796, 10.85626, 21.55367, 19.21823, 
    -6.378387, -4.858063, -3.438812, -2.507538, -2.103363, -8.483856, 
    -7.760696, -3.057556, -6.480728, -2.142456, -2.097656, 1.364059, 
    -4.281509, 1.220047, 1.233597, 7.6922, 6.016937, 5.3414, 14.3414, 
    22.98517, 15.47032, 14.3974,
  6.91745, 0.7518311, -5.2435, -8.548706, -9.397919, -9.390381, -6.85025, 
    -5.7099, -6.97995, -2.6315, -4.066132, -8.8591, -1.125549, -9.520294, 
    -8.275787, -6.668732, 1.465363, -3.353912, -6.559875, -0.734375, 
    7.583328, -13.7776, -12.79375, -10.67317, -1.351822, 15.74637, 25.91302, 
    22.59583, 3.758087, -11.44766, -1.768219, 9.952087, 16.14818, 10.25183, 
    6.433594, 10.03021, 2.611984, 3.630478, 7.631775, 3.260422, -1.481247, 
    -3.880997, -6.055191, -1.483582, -1.315643, -1.642181, -3.340118, 
    -5.381744, -7.740631, -3.393494, -1.960663, -2.730988, 0.6546631, 
    2.670074, 1.128387, 7.743469, 5.523682, 4.385162, 10.1073, 13.54846, 
    13.07059, 14.95337, 18.80963, 16.13361, 21.45676, 25.2854, 23.31146, 
    14.41379, 11.73178, 13.77551, 30.84062, 33.13542, 31.99193, 7.558868, 
    -8.203369, -8.884369, -8.519531, -6.306763, -5.764069, -5.120575, 
    -2.672943, -6.321854, -5.817444, -3.690628, -1.412491, 0.8210907, 
    3.00885, 6.354431, 4.198425, 4.711456, -2.0979, -6.386475, 0.7604065, 
    3.545319, 9.240356, 7.333862,
  -0.9575806, -2.388275, -3.545593, -4.235168, -5.342957, -6.240112, 
    -5.764038, -7.078888, -8.1315, -7.3638, -6.873444, -6.403656, -8.696899, 
    -12.97656, -14.33179, -13.23047, -6.063782, -1.647919, -0.7346191, 
    -5.1138, -9.111725, -4.513016, 1.024994, 3.078384, 9.270325, 17.04531, 
    7.036194, 12.31509, -3.751038, -13.34193, -14.38905, 3.061707, 8.193237, 
    13.47371, 8.951813, 7.787476, 10.37343, 13.50861, 11.83047, 5.685944, 
    3.13205, 1.875, -0.710144, -1.61145, -5.231506, -4.803131, -5.110138, 
    -1.365356, -2.589844, -2.087494, -2.239075, -1.161987, -1.499725, -3.25, 
    -1.256256, -0.9440308, 0.4882813, 4.2724, 8.969269, 12.29898, 11.10989, 
    13.23203, 7.734375, 5.965637, 11.14322, 15.08698, 8.085663, 11.22397, 
    28.23724, 29.46042, 23.65834, 17.43176, 10.94714, -2.571106, -2.873444, 
    -5.974243, -8.608856, -1.61145, 2.672394, -2.0578, -3.360687, -2.651031, 
    2.551056, 2.526581, 0.0249939, 4.3013, 5.2836, 9.292969, 4.892181, 
    2.845306, -3.506531, -2.612762, -2.093994, 3.827881, 7.265381, 2.122406,
  -1.007538, 1.408081, 1.989319, -2.65625, -3.598694, -3.501831, -4.921631, 
    -4.805725, -4.710663, -5.486176, -5.452606, -6.909912, -8.483856, 
    -10.36639, -15.66589, -21.37292, -22.11771, -25.55521, -25.75964, 
    -17.43672, -16.40729, -7.647659, -4.501831, -3.465103, -2.786469, 
    -20.62213, -18.37604, 18.97057, 5.853378, -12.19244, -1.606766, 7.007034, 
    7.185944, 14.26642, 15.43021, 17.10886, 17.94193, 12.10336, 15.55911, 
    7.303101, 5.87735, 6.885406, 3.086212, -1.96225, -6.552856, -3.761719, 
    -2.523438, -2.160431, -2.044006, -2.175781, 1.792206, -1.592957, 
    -10.44452, -13.05597, -10.93123, -6.334625, 1.057022, 1.236725, -0.0625, 
    5.258087, 7.822144, 4.211456, 1.284119, -1.670319, 5.385681, 1.537506, 
    3.179413, 13.49921, 31.21146, 2.419785, -1.672668, -3.902588, -7.159882, 
    -6.114319, -9.256744, -8.041138, -5.056, -6.342194, -7.676819, -6.976318, 
    -6.119537, -5.484375, -3.938538, -2.210175, -0.2263184, 0.8354187, 
    -1.117188, 3.842712, 4.144012, 1.723938, -0.1695251, -1.53775, 0.5932007, 
    2.101044, 2.954163, 2.649994,
  0.9455872, 0.4723816, 0.7822876, -2.69165, -0.8018188, -3.033325, 
    -4.337769, -4.377869, -4.114319, -3.687256, -4.147675, -4.7229, 
    -6.037506, -6.20755, -8.177063, -12.44351, -12.68463, -15.40756, 
    -29.00418, -33.59659, -22.56561, -14.4935, 4.560165, -6.213547, 6.432556, 
    -4.147644, -25.6461, 12.37759, 14.1703, -3.411209, 4.270569, 11.43933, 
    17.86693, 13.23126, 18.38934, 16.99271, 6.606262, 6.570068, 9.238037, 
    3.796631, 2.980988, 4.366394, 7.193207, 1.649994, 0.4070129, 2.075531, 
    2.462738, 5.752075, 3.522675, -1.021881, -1.152863, -0.5971375, 
    -8.443481, -7.858337, -10.11929, -8.878113, -7.334137, -0.4005127, 
    -1.057037, -1.876282, -0.5471497, -6.708344, -6.123444, -6.646362, 
    -15.19479, -3.186707, -1.804688, 1.051025, -1.225525, -17.74036, 
    -12.47525, -8.259888, -8.230743, -5.567444, 2.383057, 0.5491943, 
    -0.5606689, -2.445313, 2.829712, -3.950256, -3.272919, -1.361481, 
    -1.235413, -8.088531, -8.344269, -0.1033936, 2.681763, -1.694519, 
    3.821106, 4.982819, 8.872894, -2.098694, 0.5481873, 0.7255249, 6.110931, 
    4.265381,
  7.036987, 4.590912, 2.546875, 0.1994629, 0.5015564, -0.2549438, -0.619812, 
    -3.47995, -3.092987, -3.144531, -1.509644, -3.464325, -4.780975, 
    -4.932526, -5.008606, -7.761719, -4.8461, -5.168243, 3.905457, -13.90259, 
    -23.22864, -22.41199, -8.579437, -5.55574, 8.446365, 13.88776, 2.197922, 
    23.17395, 21.87395, 5.525787, -5.739578, -6.914063, 4.008591, 9.4375, 
    11.57788, 9.42215, 2.589325, -0.3677063, 2.3349, 0.1041565, 5.903107, 
    1.638306, 2.901062, 2.459381, 0.8979187, 5.98175, 4.510681, 4.007294, 
    3.185669, 3.196106, -0.1057434, -0.745575, -2.164856, -6.598969, 
    -3.861206, -3.852356, -4.404419, -3.253662, -1.574738, 0.6820068, 
    -2.329163, -3.989838, -7.390106, -25.53647, -9.860413, -7.42865, 
    -2.036713, 4.614075, -13.65884, -17.25443, -6.532532, -2.668243, 
    -4.390625, 2.247131, 10.53488, 2.081757, -2.664063, 2.13855, 1.507294, 
    5.075012, 5.472137, 4.925018, -1.961975, -2.7901, -0.497406, -4.495575, 
    -5.411194, 0.3026123, -1.167175, -0.2400818, 2.298431, 6.0354, -12.49323, 
    -2.0112, 0.1864624, 7.561188,
  5.15155, 13.83176, 11.50571, 10.81302, -0.8948059, 0.6270752, 1.515625, 
    -1.569275, -0.3890686, -1.437744, -2.973694, -3.777344, -3.451324, 
    -0.1593628, -4.84375, -7.340881, -6.046082, -4.985931, -1.014069, 
    3.422394, -2.566162, -0.9494934, 2.610413, -4.848694, 1.280212, 9.846359, 
    -3.090118, -7.864319, -5.530472, -5.403641, -3.069275, -10.07918, 
    -14.95729, -14.04454, -6.623962, -0.1695251, 0.9203033, 1.229935, 
    -1.175262, 1.55545, 0.6846313, -2.678131, -6.459641, -6.617447, 
    -8.516678, -8.157288, -6.177094, 0.7640381, 0.05105591, 3.345062, 
    6.753113, 5.671356, -0.8041687, -2.927094, 2.657043, 6.869263, 2.023682, 
    4.884613, 3.726044, 3.765076, 4.916931, -1.066132, -6.883331, -7.319275, 
    -9.990875, -9.924744, -7.411957, 0.7565002, -2.889313, -6.755219, 
    -5.727081, -6.050262, -0.473175, 3.595306, 3.471863, -2.18985, -5.851044, 
    -4.057007, -0.04425049, 2.349487, 6.021881, 2.020569, 5.298462, 10.1008, 
    2.097137, -1.610138, -1.377869, 1.509888, 1.160156, 3.306763, -0.4960938, 
    4.665619, -3.239044, -10.48801, -0.9536438, 0.4570313,
  14.34869, 7.6521, 5.271606, 12.06821, 12.56482, 6.898163, 3.831482, 
    3.586731, 8.375519, 5.453918, 1.054688, 4.425262, 1.894775, -0.3757935, 
    -3.379425, -2.217682, -6.197632, -7.235687, -5.3909, 7.07785, 20.44061, 
    4.751038, -4.194, -1.462494, 0.9778748, -2.701843, 1.58255, 5.5159, 
    -1.219513, -6.802063, -0.9520874, -1.4151, -14.06979, -17.55363, 
    -17.10156, -13.97369, -3.590622, -2.532547, -3.552078, -1.089584, 
    0.4822998, 1.280472, -2.684113, 0.0789032, -3.720581, -8.641144, 
    -9.055725, -7.092194, -11.63124, -8.091156, -3.972397, 2.450256, 
    5.970322, 1.559891, -1.739838, -2.5737, -1.881516, 1.300781, 2.626556, 
    1.330963, 4.150024, -2.199738, 2.353668, -1.401031, -6.700256, -10.88647, 
    -10.54272, -7.927856, -1.694794, -3.967957, -0.2244873, 0.7382813, 
    4.301819, 3.014862, -1.513794, 1.100006, -0.7835999, -3.20105, -2.035431, 
    -1.783081, 1.090363, 4.313293, 7.933319, 3.822144, 2.120575, -10.6026, 
    -11.41223, -7.267944, -7.490875, -0.1611938, 1.866669, 2.024994, 
    3.717468, 3.367462, 3.934631, 7.233063,
  30.70702, 3.293732, 8.790375, 13.78543, 6.246338, 23.59637, 14.3703, 
    8.690369, 7.157562, 4.735687, 5.580475, 10.7901, 10.61823, -2.696106, 
    -4.643494, -6.0802, -7.016663, -8.526581, -7.440613, -4.496887, 
    -1.335938, 4.421875, 2.387482, -0.731781, -2.827087, -3.679688, 
    -1.220551, 5.379669, 2.9664, 6.258331, 4.753662, 1.754669, -3.1492, 
    -9.303131, -12.92709, -15.49844, -9.27916, -6.639313, -3.941925, 
    -1.450516, -3.252853, -4.019531, 1.455719, 1.046616, -0.129425, 
    -5.418747, -5.639587, -0.7596436, -6.367188, -12.83699, -6.719788, 
    -7.016678, 1.875778, 3.011719, -0.2322998, -1.345581, -1.24115, 2.380997, 
    0.04243469, 4.120575, 4.134094, -2.846375, 6.471893, 13.19089, 25.53882, 
    9.567719, -1.1427, -1.730743, -5.405457, -0.5739746, 0.9346313, 2.457031, 
    3.064331, 2.998444, 3.454163, 7.950775, 11.99063, 4.345551, 3.596863, 
    3.399475, -3.132553, 0.518219, -0.3476563, -2.222137, 1.944519, 
    -9.045822, -11.28699, -3.378662, -8.348175, -3.269775, 4.188019, 
    -1.329712, -7.327332, 16.76849, 25.86899, 40.76874,
  33.03697, 23.07005, 39.28801, 29.8414, 8.440613, 7.263535, 8.958344, 3.263, 
    2.045563, 2.437225, 1.081238, 8.498962, 10.93906, 6.806763, -2.368225, 
    -5.250519, -8.436737, -6.948181, -3.986694, -4.492432, -4.325806, 
    -2.172394, 1.057312, -1.896881, -6.023956, 0.9484558, -3.4552, -5.689087, 
    -1.129669, -2.774719, -8.6539, -11.90494, -8.817429, -6.728653, 
    -10.34323, -10.48334, -11.35886, -10.89922, -10.72995, -10.34819, 
    -11.5414, -10.36902, -5.611725, -4.275253, -2.984894, -4.598694, 
    -5.018753, -3.309631, -1.318222, -1.862762, -2.801041, -4.221085, 
    -1.813553, 2.140625, -3.360672, -2.99765, -1.196091, -0.8726654, 
    -0.7307281, -1.035934, -1.297653, -4.143753, 11.03778, 18.05182, 
    28.97919, 32.17993, 13.95392, 12.3909, 11.1008, 2.468231, -2.742432, 
    0.4064941, 5.59375, 7.160675, 8.369781, 8.38385, 4.197144, 9.952087, 
    10.7487, 6.300247, 4.640106, -0.9635468, -9.730728, -13.62604, -5.257294, 
    -9.280731, -13.36615, -5.15625, -9.154938, -13.50259, -1.214584, 
    5.603394, -0.09243774, -1.028625, 12.88202, 30.11954,
  20.70522, 27.06067, 22.66978, 7.567444, -1.739838, -5.016937, -5.443237, 
    3.226563, 4.762482, 2.435425, -5.159119, -7.637756, -5.032806, 1.272888, 
    3.427338, 4.912506, -5.406006, -8.345581, -6.671875, -12.21899, 
    -8.034637, -7.7099, -10.4953, -9.81015, -7.222412, -8.66745, -6.955475, 
    -10.91615, -16.23828, -16.84245, -18.77759, -20.29375, -16.93254, 
    -12.98308, -11.94818, -15.12891, -13.53072, -8.073441, -5.885422, 
    -11.29245, -6.93515, -4.06694, -5.585678, -8.676834, -2.441406, 5.380997, 
    4.505722, 3.389328, 5.506775, 5.005737, 5.336975, 3.669785, 1.364578, 
    -2.320053, -4.124481, -1.755981, -1.983078, -0.3367157, 0.8622284, 
    0.3695374, -4.816925, -3.421097, 11.45157, 17.46353, 23.11041, 23.63933, 
    17.40727, 17.23517, 11.27136, 8.837524, 7.547119, 5.891922, 6.349213, 
    6.990097, 13.48698, 15.55078, 14.10573, 8.221344, 7.9599, 3.75885, 
    0.08984375, 6.161972, -0.2804718, -1.120834, -4.446625, -3.184891, 
    -7.749741, -12.54141, -8.668488, -6.630478, -9.734375, -5.885422, 
    -2.0802, -5.751556, -3.833069, 4.542694,
  7.318497, -5.393478, 1.865372, 13.07552, 11.62474, 14.67474, 5.898178, 
    -2.121628, -3.158859, -5.08255, -1.516403, 0.2992096, -6.368744, 
    -9.103394, -8.772644, -12.23048, -15.34402, -10.29636, -7.856781, 
    -10.45807, -7.629425, -8.932312, -2.922409, -1.471619, -6.052597, 
    -3.784637, -4.582809, -10.61848, -11.59375, -17.05989, -23.10573, 
    -27.9711, -18.8349, -12.64687, -7.642715, -10.07188, -13.71432, 
    -6.509644, -1.260422, -6.24765, -8.069519, -2.998703, 0.3419342, 
    -4.911987, -7.139572, 1.576553, 4.679428, 2.579163, 6.022919, 6.822403, 
    2.311722, 4.234894, 7.052094, 7.849213, 2.225525, -3.517456, -3.769012, 
    -1.947403, -3.469788, -2.984375, -3.057556, 4.091934, 4.213272, 3.000259, 
    3.311707, 0.4947968, 0.8489532, 7.016403, 6.318756, 6.728653, 1.753647, 
    0.1679688, 1.628387, 3.346619, 6.094009, -9.784103, 12.34401, 3.610153, 
    3.598694, 6.8638, 5.871368, -4.78775, -5.186722, -4.506775, -10.13957, 
    -11.84662, -10.90051, -15.04871, -14.50624, -7.400253, -7.549744, 
    -8.448959, -5.284378, -5.614075, 2.693222, 8.316666,
  -3.885406, -7.154678, -10.07603, 4.372665, 11.30469, 6.367706, 1.728394, 
    -0.1609344, -11.82135, -7.71225, -5.710678, -2.950531, -12.43359, 
    -17.93152, -19.61458, -22.70181, -20.12657, -10.22917, -5.300522, 
    -6.061462, -6.234894, -2.672394, -3.244797, -4.4711, -3.56041, -13.38411, 
    -13.869, -14.67812, -10.23932, -7.258606, -15.41615, -16.38776, 
    -7.127335, -0.5984497, -0.1552124, 2.677612, -0.8932343, -6.052078, 
    -0.3538971, -0.5572968, -11.49037, -6.253647, 4.637772, 4.243484, 
    1.308594, 5.311462, 5.169022, 3.169785, 7.009109, 11.14427, 12.24141, 
    5.545319, 4.234116, 12.03723, 9.885422, 3.621613, 1.615875, 2.018219, 
    -2.780991, -3.184372, -3.132553, -0.5836029, 2.166924, -0.0177002, 
    -3.638275, -7.692703, -8.736191, -7.134628, -2.192184, -3.143753, 
    -3.648697, -6.807297, -26.72812, -30.29218, -28.40703, -28.56276, 
    -4.512497, -7.860931, -8.423706, 1.867706, -1.098694, -4.874222, 
    -7.839584, -7.616669, -6.615372, -2.319, -3.333328, -4.987503, -8.113022, 
    -10.3237, -5.020569, -3.701309, -9.672913, -12.46146, -9.060944, -3.675262,
  -14.09949, -10.12135, 1.748688, 15.30573, 10.61458, 3.033844, 4.547134, 
    -0.413269, -2.552078, -4.935928, -5.875519, -2.949478, -6.364578, 
    -7.80365, -2.777863, -0.4028778, -1.548447, 0.7263031, 6.034882, 
    6.924484, 10.33308, 9.727859, 11.81822, 12.17265, 3.603378, 1.720566, 
    -7.31041, -7.668228, -5.834122, -7.331253, -10.52682, -10.9185, 
    -5.024475, -4.279694, -3.141144, -2.730209, 0.4476471, 5.228119, 
    -0.0388031, -3.353134, -4.095322, -1.069275, 4.928391, 4.008072, 
    6.179169, -0.4247437, -0.9567719, -4.536728, -0.3528748, 3.378128, 
    7.326035, 12.66354, 13.85312, 10.94218, 3.852615, 0.9684753, -0.1588593, 
    -1.386978, -5.278381, -3.391403, 4.711472, 4.847397, -1.294792, 
    -9.189316, -12.40234, -12.01353, -7.801041, -5.112503, -1.321625, 
    -9.005478, -11.04115, -16.2724, -22.64166, -31.45079, -34.76979, 
    -30.33775, -11.09036, -8.225769, -25.33281, -15.60052, -7.675781, 
    -12.56041, -15.07214, -8.745056, -0.8653564, 1.326035, 2.720306, 
    -0.154953, 1.872665, -0.9640656, -3.886719, -3.184387, -4.108597, 
    -4.250519, -7.220566, -12.96536,
  -17.21797, -18.12994, -8.429153, -1.848709, -3.545822, -5.2052, -6.902344, 
    -2.489059, -3.294525, -4.013809, -2.924744, -3.589844, -3.228897, 
    -2.304688, -5.197906, -5.475769, -1.757813, 3.136459, 7.734634, 11.825, 
    9.390106, 9.8573, 6.496628, -0.9804688, 1.555481, 5.200516, 5.591415, 
    5.032028, 1.03775, -3.586975, -2.4039, 3.962769, 2.904938, -1.844528, 
    -6.2323, -5.014587, -4.554428, -4.132294, -7.886978, -13.8802, -13.9263, 
    -14.35886, -10.40886, -5.191925, -4.267441, -3.412231, -0.1778717, 
    -2.958588, 0.1031342, 4.276825, 3.285934, 1.167969, 5.226044, 4.784378, 
    2.347916, -1.031509, -3.241135, -1.992706, -0.2424469, -3.806519, 
    -9.0177, -9.673431, -12.21329, -17.88828, -13.95886, -6.078644, 
    -4.156769, -3.689316, -3.842453, -9.035416, -7.194794, -4.878906, 
    -8.555984, -13.11563, -32.97969, -35.75313, -25.61926, -17.44167, 
    -21.44662, -24.0177, -32.82579, -28.72656, -21.54063, -13.44818, 
    -4.647919, 3.11171, 11.99063, 13.06172, 10.3526, 5.088028, -8.330215, 
    -13.4724, -10.5901, -3.378906, -4.105469, -9.445053,
  -1.663284, -2.986984, -8.475006, -13.18698, -16.71771, -12.66745, 
    -7.389847, -7.942184, -11.26797, -13.18854, -12.83047, -13.7224, 
    -12.29089, -14.41277, -18.12474, -17.02995, -10.93906, -3.037766, 
    7.010422, 10.84323, 11.09921, 12.00887, 12.19296, 12.57603, 9.708084, 
    6.257019, -1.013809, 0.2398376, 5.34166, 9.517441, 6.234894, 3.388275, 
    -1.757294, -5.43959, -9.878387, -7.613541, -7.834381, -13.25548, 
    -16.01381, -22.92995, -26.79401, -26.55415, -24.71484, -23.42293, 
    -22.47162, -16.08046, -12.78645, -16.68933, -21.90079, -27.02422, 
    -25.86119, -20.51772, -16.95157, -4.987244, -2.322922, -1.961975, 
    -4.873444, -8.09166, -10.94896, -16.42863, -26.24374, -30.28593, 
    -30.33749, -27.68411, -20.20573, -12.48984, -1.640625, 2.430206, 
    -0.2093811, -5.66745, -2.096619, -7.311203, -17.62839, -32.0526, 
    -31.74011, -37.29688, -24.92317, -24.99454, -32.66251, -44.44115, 
    -37.48465, -23.96277, -18.94035, -11.79898, -0.4739532, 6.253906, 
    9.298431, 6.876297, 0.8242188, -5.344528, -17.71484, -20.87943, 
    -17.70416, -9.86171, -3.203644, -1.117462,
  -9.830475, -8.004684, -6.704697, -8.760162, -13.01146, -14.21616, -14.2948, 
    -16.64844, -19.42188, -20.44687, -17.33359, -14.6651, -13.494, -16.36693, 
    -22.7289, -21.81953, -31.35156, -25.24271, -18.80026, 0.7346344, 
    8.764313, 13.3513, 14.39922, 12.80521, 8.050781, 5.570053, 3.701294, 
    9.196091, 15.825, 15.98358, 14.16771, 10.69583, 5.120834, -2.593216, 
    -6.173187, -7.703644, -6.808075, -7.459366, -6.824738, -7.487244, 
    -13.6414, -17.44141, -17.12344, -13.74089, -12.64401, -17.14168, 
    -19.69089, -21.41458, -21.38152, -18.79662, -13.50287, -10.68776, 
    -11.02423, -13.6711, -15.04478, -14.05547, -13.31796, -11.04636, 
    -13.7487, -18.06537, -23.92267, -27.92265, -27.31902, -14.48724, 
    -9.625259, -6.185684, -2.038025, -3.546875, -7.431503, -12.16223, 
    -17.10338, -21.58151, -25.55391, -32.3013, -31.16223, -28.04036, 
    -16.89896, -32.56354, -34.86354, -35.05963, -30.85312, -23.65497, 
    -20.63904, -18.61145, -16.59296, -17.33255, -15.52759, -11.72238, 
    -11.29401, -14.57187, -21.37944, -27.74687, -24.73906, -19.73463, 
    -13.50208, -13.16953,
  -11.77499, -8.641937, -4.945313, -3.776566, -3.750519, -2.481506, 
    -5.885666, -15.08411, -18.20833, -22.04765, -24.28802, -24.31459, 
    -23.38464, -24.73126, -24.52968, -22.22395, -17.88724, -14.82864, 
    -10.91536, -8.002869, -8.941406, -9.782822, -10.01015, -7.603897, 
    -3.703125, -1.031509, -1.629944, 2.054947, 4.988281, 4.399216, 0.2382813, 
    -8.546097, -10.75183, -10.34323, -11.10651, -11.35001, -9.958862, 
    -10.14088, -11.84584, -15.41016, -18.09973, -19.09114, -19.25494, 
    -18.97656, -18.65962, -18.4388, -19.24869, -19.96536, -18.73907, 
    -17.69896, -15.59557, -16.63959, -17.82214, -19.36797, -20.07864, 
    -19.97943, -20.24428, -20.20911, -19.16302, -20.27031, -22.09479, 
    -25.90364, -30.41745, -38.15157, -42.54453, -36.58385, -38.0625, 
    -38.47682, -37.82396, -39.82109, -41.26042, -34.79922, -28.04793, 
    -19.32318, -11.77577, -20.55208, -21.54663, -26.02084, -18.99792, 
    -20.54947, -21.30652, -21.46017, -18.41821, -17.16617, -15.64688, 
    -15.16223, -18.69818, -23.48462, -25.04974, -26.46301, -27.67993, 
    -35.3578, -43.6875, -43.29845, -30.9151, -17.1935,
  -28.36432, -28.00391, -25.4828, -23.29767, -5.032028, -4.520828, -4.902863, 
    -26.77866, -25.22969, -23.11484, -20.81302, -17.76746, -15.96745, 
    -14.86562, -14.98593, -15.43985, -13.6599, -13.95781, -15.58594, 
    -15.86302, -17.2849, -17.71381, -17.34923, -15.43698, -11.47656, 
    -5.420822, -5.890625, -12.8513, -11.34818, -10.21303, -9.136719, 
    -7.236206, -5.512238, -1.459122, 1.389328, 3.22995, 0.1997375, -3.975784, 
    -9.368744, -13.94557, -17.97162, -22.05782, -23.56302, -23.41928, 
    -21.11198, -18.36745, -15.80469, -13.19687, -11.61067, -12.47969, 
    -14.97995, -18.59818, -21.78568, -24.14244, -27.09245, -29.84921, 
    -31.5177, -29.97527, -27.88594, -23.72917, -20.59869, -19.36276, 
    -19.62839, -21.02786, -24.62553, -28.05469, -30.24582, -28.78542, 
    -25.53699, -19.97371, -14.85651, -1.584381, -7.009644, 1.831772, 
    3.396622, 3.993759, 4.925003, 6.344269, 6.629684, 4.463272, 0.6197815, 
    -3.497406, -5.830994, -7.742188, -9.458588, -12.08905, -15.99817, 
    -19.51248, -21.89948, -24.88541, -26.66406, -29.50574, -43.75259, 
    -42.53645, -35.73595, -30.65625,
  -6.918488, -5.914063, -6.130478, -6.310944, -6.697922, -8.475266, 
    -10.45807, -12.24167, -12.84349, -12.9151, -13.03125, -13.17239, 
    -13.87553, -13.66563, -13.12109, -11.90755, -9.464325, -8.903641, 
    -8.823181, -8.728653, -9.148438, -9.235687, -7.945572, -6.570572, 
    -5.895569, -6.177612, -5.434113, -3.944519, -2.855988, -2.995575, 
    -3.164322, -3.523956, -4.644791, -7.019272, -10.57709, -12.45703, 
    -14.05234, -15.06302, -16.67162, -16.71823, -17.44011, -17.5513, 
    -18.99948, -20.28073, -21.83958, -22.26692, -21.494, -20.92397, 
    -21.02318, -20.43645, -20.81172, -21.22578, -21.92787, -22.52109, 
    -23.39479, -24.15962, -24.31772, -24.27579, -23.73828, -22.62343, 
    -22.39035, -22.30754, -23.29219, -24.34349, -24.43282, -25.07422, 
    -26.9612, -28.00052, -29.96538, -30.45338, -30.50548, -30.13542, 
    -28.99271, -27.57317, -26.39738, -24.91432, -23.20808, -19.72604, 
    -16.94218, -14.61459, -12.58594, -12.11014, -12.06824, -12.7198, 
    -13.52786, -16.18256, -17.72656, -21.24715, -22.68671, -22.99922, 
    -23.05312, -22.08099, -18.70703, -16.50963, -12.87032, -9.153122,
  -25.82838, -25.26588, -25.2224, -24.7289, -24.08827, -23.79713, -24.3336, 
    -24.13881, -24.25677, -23.85025, -23.86511, -23.56042, -22.46536, 
    -21.24272, -19.73463, -18.42004, -17.22266, -15.7224, -14.77266, 
    -14.1086, -13.41484, -12.50104, -12.00444, -11.92447, -11.77344, 
    -11.52579, -11.48724, -12.26797, -12.94818, -13.54402, -14.27943, 
    -14.93333, -15.62057, -16.69531, -18.11511, -19.39427, -20.54271, 
    -21.32813, -21.9724, -22.61406, -23.66512, -24.53854, -25.33516, 
    -25.5237, -25.16536, -25.08958, -24.96068, -24.32942, -23.61354, 
    -22.84192, -22.13907, -21.45078, -20.76381, -20.12839, -19.81198, 
    -19.59636, -19.97058, -20.5573, -20.92526, -20.78645, -21.31328, 
    -22.29349, -22.77786, -23.06848, -22.76875, -22.74113, -22.1013, 
    -21.97005, -22.01692, -22.51563, -22.55182, -22.40651, -21.96588, 
    -22.28569, -22.325, -21.97136, -21.63542, -21.3974, -21.93803, -22.92319, 
    -23.65392, -24.15886, -23.54688, -23.82239, -23.65938, -24.29634, 
    -24.45988, -25.04271, -25.84792, -26.80547, -27.03021, -27.05676, 
    -26.79323, -26.58255, -26.25365, -26.16797,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -0.004687499, -0.006510418, -0.008593753, -0.009374999, -0.009635417, 
    -0.01041667, -0.008854166, -0.005468749, -0.003385417, -0.004947916, 
    -0.006770831, -0.0078125, -0.007031251, -0.005208336, -0.006249998, 
    -0.004166666, -0.003125001, -0.00390625, -0.002604168, -0.002864581, 
    -0.004166666, -0.006250001, -0.0078125, -0.008854168, -0.006510416, 
    -0.006770832, -0.006510416, -0.007552082, -0.004427083, -0.006250001, 
    -0.007552084, -0.006250001, -0.004427083, -0.004427083, -0.002864584, 
    -0.004947916, -0.005208334, -0.005989583, -0.007552082, -0.007552082, 
    -0.007812498, -0.006770834, -0.006510416, -0.007031251, -0.005729165, 
    -0.00390625, -0.002864584, -0.004427083, -0.004166666, -0.005729167, 
    -0.004166668, -0.003125001, -0.003125001, -0.00546875, -0.005208332, 
    -0.01119792, -0.01510417, -0.0171875, -0.015625, -0.0109375, 
    -0.007812502, -0.006510418, -0.006249998, -0.004687499, -0.003906248, 
    -0.0007812511, -0.003385417, -0.00390625, -0.003385417, -0.004427083, 
    -0.003125001, 0, 0.003125001, 0.001822917, 0.0007812493, -0.0002604164, 
    -0.0005208328, 0.001302084, 0.002343751, 0.0007812493, -0.002083333, 
    -0.004166666, -0.00234375, -0.003645832, -0.004427083, -0.003385417, 
    -0.004166666, -0.003385417, -0.003385417, -0.001302084, -0.0002604183, 
    0.001822915, 0.001041666, 0, -0.0002604164, -0.002083335,
  -0.15625, -0.1700521, -0.1880209, -0.2117188, -0.1921875, -0.1768229, 
    -0.1348958, -0.109375, -0.09218752, -0.1, -0.10625, -0.09479165, 
    -0.1023438, -0.09010422, -0.05208337, -0.01458335, -0.006510496, 
    0.01041675, -0.01901042, -0.0135417, -0.01796877, -0.04739583, 
    -0.04947913, -0.0575521, -0.06380212, -0.0703125, -0.06406248, 
    -0.0617187, -0.02031255, -0.02369785, -0.06223965, -0.06796873, 
    -0.09531248, -0.1145834, -0.1200521, -0.1348959, -0.1148437, -0.09218752, 
    -0.0830729, -0.1033853, -0.1622396, -0.2065104, -0.2184896, -0.2476562, 
    -0.2559896, -0.2416667, -0.2416667, -0.2184895, -0.2140626, -0.1994792, 
    -0.1671875, -0.1263021, -0.1179687, -0.1023437, -0.09244788, -0.115625, 
    -0.1085937, -0.05911458, -0.07604164, -0.07265627, -0.07708329, 
    -0.06953126, -0.08072919, -0.1182292, -0.07005209, -0.03177088, 
    -0.02578127, 0.006770849, 0.01718748, 0.01822919, 0.007552087, 
    -0.006250024, 0.009635448, 0.04218751, 0.06015623, 0.03958333, 
    0.006770849, -0.03046876, -0.08177078, -0.1091146, -0.09531254, 
    -0.1377604, -0.1177083, -0.1148437, -0.08020836, -0.04765624, 
    -0.06588542, -0.06718749, -0.1072916, -0.09843749, -0.1242187, 
    -0.1463541, -0.1257813, -0.1111979, -0.1117187, -0.1268228,
  -0.4533854, -0.5523438, -0.573698, -0.6234374, -0.6033854, -0.6161456, 
    -0.5528646, -0.5429688, -0.4679685, -0.4726563, -0.4539065, -0.3617187, 
    -0.2567711, -0.1846356, -0.0562501, 0.01510429, -0.04348946, -0.1799479, 
    -0.1083331, -0.1343751, -0.2286458, -0.3273439, -0.3312497, -0.2940106, 
    -0.2364583, -0.1221356, -0.1401043, -0.1557293, -0.1369791, -0.1330729, 
    -0.0859375, -0.01822948, 0.03645849, -0.03828144, -0.1088543, -0.1125002, 
    -0.1075521, -0.06328106, -0.1158857, -0.2307291, -0.3398438, -0.4513021, 
    -0.50599, -0.4424477, -0.3565106, -0.2835937, -0.3109374, -0.3354163, 
    -0.4190102, -0.4036458, -0.4403646, -0.4377604, -0.4382811, -0.4554689, 
    -0.4380207, -0.5460935, -0.6666665, -0.7054687, -0.6242187, -0.515625, 
    -0.3479166, -0.3773439, -0.3622396, -0.2932293, -0.2533851, -0.1427083, 
    -0.05286455, -0.05911446, -0.09427071, -0.1690104, -0.1614585, 
    -0.2216146, -0.2424479, -0.1570313, -0.2458334, -0.4513023, -0.3697917, 
    -0.4960938, -0.3895833, -0.3010418, -0.3585939, -0.4117188, -0.4546874, 
    -0.5208333, -0.5765626, -0.4828124, -0.4382813, -0.2658854, -0.1770833, 
    -0.2585938, -0.3320315, -0.2460938, -0.1885417, -0.1942711, -0.2234373, 
    -0.309896,
  -0.604948, -0.7138023, -0.9044266, -0.916667, -0.9398441, -0.6372395, 
    -0.3877602, -0.546875, -0.9473963, -0.9666672, -0.7309895, -0.3934898, 
    -0.5072918, -0.5765619, -0.7570314, -0.5473967, -0.3921871, -0.04374981, 
    -0.01744747, -0.06145859, -0.2471352, -0.2380209, -0.160677, -0.1575527, 
    -0.05520821, -0.06692791, -0.2049475, -0.01614571, -0.1744795, 
    -0.004947662, -0.03151035, -0.006250381, -0.1468744, -0.2653646, 
    -0.3552084, -0.2401037, -0.1966152, -0.1802082, -0.3861971, -0.5643234, 
    -0.7028646, -0.7799473, -0.9195318, -0.8929691, -0.9773436, -1.033072, 
    -0.6731768, -0.682292, -0.9187498, -0.9817705, -0.9559898, -0.6747398, 
    -0.6955738, -0.8427076, -1.009376, -1.0625, -1.351042, -1.48151, 
    -1.567449, -1.395052, -1.127864, -0.9169264, -0.8343744, -1.174219, 
    -1.540886, -1.285677, -1.155729, -1.346094, -1.239583, -1.333333, 
    -1.079166, -0.7643232, -0.5315104, -0.03255272, -0.3888025, -0.8479166, 
    -1.158854, -1.617448, -1.547396, -1.120313, -0.8989582, -0.8898439, 
    -0.8770838, -0.9111977, -0.8307295, -0.8924484, -1.059375, -0.7171869, 
    -0.4729166, -0.353385, -0.4179688, -0.2723961, -0.2510414, -0.2893229, 
    -0.4911451, -0.6138029,
  -1.455467, -1.701822, -1.838541, -1.878124, -1.986717, -1.671614, 
    -1.052343, -0.938282, -1.289324, -1.280468, -1.167448, -1.358854, 
    -1.67474, -2.135157, -1.886978, -1.20599, -1.162239, -1.46224, -1.698177, 
    -1.548437, -1.458593, -0.869791, -0.988802, -1.316927, -1.220312, 
    -0.8312492, -0.207552, -0.3468742, -0.2638016, -0.386198, -0.04921913, 
    0.1455727, -0.08671951, -0.3278646, -0.5158854, -0.8161459, -1.039063, 
    -1.599218, -1.601302, -1.664063, -1.917187, -1.904947, -1.777604, 
    -1.501041, -1.558073, -1.426042, -1.847917, -1.68828, -1.702345, 
    -1.167969, -1.264845, -0.958333, -1.029427, -1.040626, -1.253386, 
    -1.024479, -1.012501, -1.487761, -1.019011, -0.8453121, -0.4804688, 
    -0.2585945, -1.011719, -1.986719, -2.722136, -2.641146, -2.082031, 
    -2.049219, -2.680208, -2.816926, -2.61224, -3.31901, -3.096875, 
    -2.860676, -2.796354, -2.620573, -2.343749, -2.586458, -2.349739, 
    -2.341667, -2.378906, -2.839064, -2.456251, -2.234636, -1.66823, 
    -1.633074, -1.594532, -1.577343, -1.19297, -1.257553, -1.358593, 
    -0.6981773, -0.2437496, -0.500782, -1.03828, -1.454687,
  -3.435677, -3.447657, -3.415104, -3.448957, -2.990625, -2.932293, 
    -2.517447, -2.995052, -3.328384, -2.766407, -2.406252, -1.994793, 
    -2.300261, -3.091406, -3.264322, -3.651302, -4.493229, -4.571613, 
    -4.308594, -2.622135, -1.660938, -1.925781, -2.521875, -2.788019, 
    -2.916666, -2.946875, -1.871094, -0.8864574, -0.6911469, -0.3643227, 
    -0.848177, -1.498438, -1.108852, -0.3684902, 0.3156242, 0.3606758, 
    -0.4236984, -0.8783855, -1.315363, -0.7361965, -0.6549473, -1.065365, 
    -2.008333, -2.614584, -1.88776, -1.441927, -1.003645, -1.483072, 
    -1.244011, -0.8210945, -0.7583332, 0.005729675, 0.4598961, 0.5627613, 
    1.35, 1.432032, 1.29974, 0.9359379, 0.2104168, -0.907032, -1.845053, 
    -2.310158, -2.38073, -2.201822, -2.374218, -1.929688, -2.065105, 
    -2.677343, -3.717186, -3.319271, -2.422134, -2.645573, -3.358595, 
    -3.128906, -2.429167, -2.441147, -2.603645, -2.890364, -2.748438, 
    -2.253906, -2.545832, -3.300261, -4.085417, -3.626562, -2.820833, 
    -2.934114, -2.790886, -2.454166, -1.34948, -1.496353, -2.758333, 
    -2.811459, -1.679426, -1.11146, -1.676304, -2.628386,
  -2.678909, -3.420052, -4.796616, -5.272659, -6.014584, -5.576302, 
    -4.332031, -4.343227, -5.320835, -5.769531, -4.359634, -3.042969, 
    -4.068752, -6.113541, -5.982811, -7.365364, -8.355469, -7.61198, 
    -6.092449, -4.327084, -4.167187, -3.541405, -3.427341, -3.21328, 
    -3.439064, -3.169273, -3.589321, -2.427341, -2.942448, -3.168228, 
    -3.046875, -1.552864, -1.298698, -0.8067722, -0.6971359, -0.967186, 
    -0.4963551, -0.2393227, 0.06588745, 0.108593, -0.609375, -1.333595, 
    -2.042969, -1.998436, -0.2479172, 0.311718, 0.8841133, 0.5888004, 
    -0.798439, -0.7497406, -1.54427, -2.155729, -1.677605, -0.8031273, 
    -1.073175, -1.081253, 0, -0.1752625, 0.1059875, 1.466927, 0.3645859, 
    -0.7567711, -1.067707, -0.3994827, -0.3432274, -0.8052101, -0.9385414, 
    -0.0388031, 0.3263016, 0.002603531, -0.6783867, -1.386978, -1.328125, 
    -0.7841148, -1.211718, -1.31901, -0.9973965, -1.332031, -1.09375, 
    0.2752609, 1.064064, 1.496614, -0.9414063, -2.394531, -2.700001, 
    -3.896614, -4.691929, -4.31823, -2.771873, -2.386459, -3.417709, 
    -3.945313, -3.54948, -3.533073, -2.402866, -1.467968,
  -4.338802, -4.364582, -4.489063, -3.534115, -3.235676, -3.25729, -1.872395, 
    -0.5367203, -0.5291672, -3.071354, -2.987499, -1.083595, -1.190102, 
    -1.480206, -1.325001, 0.3148422, 0.3351555, -0.3494797, -1.889061, 
    -3.399738, -4.597397, -3.479691, -1.69453, -1.392189, -1.465626, 
    -0.9570313, -1.729164, -1.04948, -0.800518, -1.117188, -1.927345, 
    -1.788803, -0.8143196, 0.5557289, 1.039063, 0.9148445, 0.1255226, 
    -0.1807289, -0.2520828, -0.02682114, -0.3677063, -0.4510422, -0.8549461, 
    -1.684635, -0.6622391, 0.7523422, 0.2994804, -1.640888, -1.167187, 
    0.4997406, -0.2765656, -0.2005196, 1.494534, 1.267967, -0.6583366, 
    -0.9244804, -1.032551, -1.60833, -0.8476563, 2.108334, 2.603905, 
    1.223961, 0.5999985, 0.7458305, 0.9713554, 2.0112, 1.207554, -0.6999969, 
    -0.01328278, 0.3822937, -0.5325508, -0.8627625, -1.100784, -1.335419, 
    -2.489323, -2.344013, -0.4049454, -1.851822, -2.008335, -0.1697922, 
    1.084373, 2.104427, -0.05182266, -0.2080727, -1.938282, -1.230209, 
    -0.9825516, -1.925781, -2.765625, -2.46172, -2.470573, -3.16172, 
    -3.422657, -4.636719, -4.924999, -4.199478,
  1.264584, 0.216404, -1.211197, -2.025261, -1.269791, 1.481251, 1.049217, 
    0.1885414, -1.038284, -1.396614, -1.331512, -0.4229164, 0.7473946, 
    -1.144531, 0.515625, 0.6026039, 0.8088531, 0.1611977, -1.26276, 
    -1.818489, -0.3718758, 2.328125, 2.375782, 1.38047, 1.869789, 0.3333321, 
    -1.665886, -1.162239, -0.7750015, -0.4023438, 0.1531219, 0.2747383, 
    -0.5471344, -0.282032, -0.8315125, -1.615364, -3.129948, -1.859116, 
    0.985939, 1.079685, -0.6833305, 0.8135414, 1.87656, 0.8763008, 0.5289078, 
    2.159893, 1.587238, -0.2184868, -0.3968735, 0.2091141, -0.2398453, 
    -0.9575539, 0.3481789, -0.8554688, -2.169529, -0.4106789, -0.5101585, 
    -1.402344, 0.8591156, -0.6494827, 0.828907, 2.94323, 2.921616, 0.8330727, 
    0.3794289, -1.458591, 1.853649, 1.459377, -0.8911476, -0.2309875, 
    2.33802, -0.1651039, -0.3723946, 0.4179688, -0.7473984, -2.001041, 
    -2.613541, -1.948959, -0.6445313, 2.037506, 2.646095, 1.453125, 1.469788, 
    0.4572906, -1.394012, -1.37344, 0.7096367, 1.818226, -0.6231766, 
    0.1843758, 0.6348953, 0.9190102, -0.1651039, -2.198177, -1.061718, 
    0.4632835,
  -1.967964, -3.533333, -3.769272, -1.869797, -2.939583, -1.569794, 
    -0.4065094, -2.5513, -2.873436, -1.5625, -1.183075, -0.3093719, -1.32917, 
    -1.425781, -1.420837, -2.947914, -1.364845, -0.09036255, 0.3651047, 
    -0.3226547, 0.549736, 0.06614685, -0.5406265, 0.7809906, 0.6705704, 
    -0.6778641, -0.8544312, 1.496353, 0.8424454, -0.673439, -0.5221329, 
    3.482292, 2.879173, 0.7276077, -0.4476547, -0.9575577, -0.9132843, 
    2.479691, 2.372658, 2.800262, 0.2786484, -1.079948, -0.6278687, 
    0.5249939, -0.0869751, 3.785679, 6.404427, 5.787239, -0.8062515, 
    -2.533073, 0.05208588, 1.477081, -0.01744843, 3.029427, 3.239326, 
    3.698441, -0.9757767, -2.064583, 1.793488, 0.003120422, 1.136978, 
    3.886719, 2.175514, 0.7833328, 1.417709, 0.2835922, 2.018486, 1.476822, 
    -0.4257813, -0.2393188, -0.776825, -0.1598969, 0.8526001, 1.763809, 
    -0.3789063, -2.587242, -0.6385422, 0.2174492, 3.261459, 2.384377, 
    0.1851578, 0.7570343, 0.4499969, -0.548439, -1.582291, -1.098953, 
    -2.131248, -0.3601532, 0.295311, 0.4265594, 1.712242, -0.1304703, 
    -1.192451, -0.07526398, -0.2697906, -1.629944,
  -1.758331, -1.882545, -1.028908, 2.378387, 1.039581, -1.19088, -2.648697, 
    -1.670052, -1.572136, -0.8380203, 2.286713, 3.360161, 2.441666, 
    0.6445313, 1.422401, -0.2554626, 0.04452515, -0.08437347, -0.1372375, 
    1.955208, 0.9604111, -0.433075, -0.9882813, 2.992188, 5.788284, 8.317451, 
    10.68151, 9.348694, 7.161453, 7.247139, 6.385941, 5.243492, 3.884109, 
    4.485413, 4.950516, 1.480209, -0.9338531, 3.552605, 4.763023, 1.074745, 
    2.220055, -2.13932, -3.164322, 1.108849, 2.691666, 1.888023, 1.905991, 
    0.03568268, -1.997398, 0.2148438, 0.3812485, 3.408592, 3.135941, 
    1.465881, 2.381516, 1.290627, 0.09557343, 1.498695, -0.2843781, 
    -2.726303, -0.03723907, -0.3596344, -1.694008, -3.088028, -1.389847, 
    0.326561, 1.041412, -1.30912, -1.978386, 0.9424438, -0.3361969, 
    -0.5601578, 0.401825, 1.860413, -0.7851563, -0.4307251, 1.206512, 
    -0.1070328, -1.609642, -1.007294, -1.53698, 1.852867, 2.701561, 
    -0.2781296, 0.1190109, -0.3666687, -3.260162, -0.9848938, 0.357811, 
    0.5989609, 0.4098892, -0.4124985, 3.417709, 1.921875, -1.296616, -1.487762,
  4.024223, 1.953644, -0.4031296, 2.590622, 1.4375, -1.856773, -2.747131, 
    -2.930984, -6.060677, -3.484375, -1.858856, 0.4348984, 4.129425, 
    4.945831, 1.39167, 2.530991, 4.603905, 3.240891, 1.805725, 1.135674, 
    0.9283829, 4.939842, 5.594788, 7.144005, 6.131775, 6.916672, 10.11198, 
    6.901566, 5.288803, 4.42057, 2.561462, 6.40078, 7.715881, 6.78672, 
    9.478905, 7.710938, 4.59584, 5.457031, 3.980469, 1.000519, 0.6815109, 
    0.3739624, -0.07500458, -1.353127, -0.439064, 2.21302, 1.153122, 
    -0.453125, -1.855469, 2.555733, 2.433853, 1.531769, 3.702087, 1.824478, 
    0.5544281, 2.091408, 2.321609, 3.397133, 0.3848953, -1.733597, 2.634636, 
    2.93959, 1.940102, 2.069008, 1.412239, -0.079422, 0.8320313, -0.342453, 
    0.6408844, 0.1174469, -5.699745, -6.284897, -1.162498, -2.950523, 
    -0.6244812, 2.622917, 7.245049, 7.367966, -0.2432251, -4.59375, 
    -1.872917, 0.249733, -2.542709, -2.662506, -4.708595, -5.116669, 
    -1.264847, -0.9768219, -2.052345, 0.7091141, 4.41745, 3.462494, 3.583855, 
    0.7088547, 3.345573, 1.800781,
  0.7679672, 3.618484, 2.9216, 5.68515, 2.359894, 1.241928, 0.8317719, 
    2.332291, 1.856522, 2.554947, 9.670578, 13.72109, 15.61406, 10.1625, 
    9.839066, 6.172401, 5.3815, 3.092453, 4.970047, 5.803642, 7.227867, 
    9.622406, 11.18282, 4.359634, 5.0224, 6.169273, 6.147141, 4.113274, 
    5.105469, 3.233337, 4.574738, 8.901566, 7.410934, 6.702087, 4.881256, 
    1.266403, 1.046089, 1.663277, -3.334641, -1.499741, 0.3710938, -3.085419, 
    -6.521355, -7.259895, -2.601563, -1.506775, -1.564583, 1.65416, 1.664063, 
    2.660934, 7.822136, 5.104683, 3.052086, 2.616402, 5.890625, 4.515106, 
    0.7315063, -2.593491, -4.632034, -3.988281, -2.165108, -7.04557, 
    -4.445831, 0.2518234, -0.0770874, -0.3197861, -0.002601624, -0.4653625, 
    2.69297, 1.190628, -3.799217, -2.575256, -2.347923, -1.513802, 
    -0.3669281, 0.6671906, 4.153137, 6.46563, -5.047928, -4.497398, 
    -1.885422, 3.039841, 1.239334, -1.747925, -1.71328, -1.817711, 2.764328, 
    3.03672, 0.91745, 4.710678, 1.059372, 1.941666, 1.767189, 3.105995, 
    4.594528, 1.073174,
  3.001038, 2.235413, 4.580215, -2.178909, -3.08255, 1.506516, 3.085159, 
    1.284637, 1.046616, 0.3052063, 5.400269, 8.961716, 6.891937, 5.107819, 
    7.521866, 7.040359, 6.216156, 2.064835, 3.006775, 1.885162, 1.774475, 
    -0.816925, -3.033859, -0.4265747, -1.633331, -1.6698, 2.230469, 1.234375, 
    0.7489624, 2.091675, 9.741394, 13.49662, 4.156769, 7.871094, 1.413284, 
    -10.89063, -6.454422, -3.638535, -9.415359, -8.703659, -8.481247, 
    -7.821884, -5.931244, 0.3434906, 2.299744, -1.016663, 1.975266, 5.488022, 
    4.675781, 3.746613, 7.659637, 1.81459, 1.771881, -2.471878, 0.5078125, 
    1.390366, -0.7606812, 1.788544, -3.475525, -2.912247, -4.421356, 
    -1.606766, -2.41172, 0.3216171, -0.3023453, 1.084633, -0.9598923, 
    -4.666145, -3.50885, -5.826302, -1.164581, -3.45105, -7.619019, 2.820831, 
    4.401306, 3.438538, 3.5336, 2.165878, -0.8796844, 1.391663, 1.735153, 
    6.72422, 5.738014, -0.04922485, 3.98204, 4.839066, 5.678116, 4.133865, 
    3.919266, 2.072906, 1.946625, -0.4007874, 3.838806, 4.157028, 3.304688, 
    2.441925,
  1.710159, 2.065369, -0.1453094, -2.716156, -1.909119, 1.77475, 3.272659, 
    1.514328, 3.516922, 1.357819, 6.497391, 8.262756, 5.291138, 5.184631, 
    5.286987, 6.5737, 1.781509, -2.549728, 0.7651062, 2.785934, 1.423965, 
    3.323441, 1.474228, -1.974487, -5.240616, -2.114578, 4.117706, 4.430725, 
    7.581253, 6.528137, 14.52213, 9.344788, 2.797394, -3.154419, -2.817184, 
    -5.46405, -10.89453, -11.42863, -12.05026, -14.73906, -17.34714, 
    -8.38855, 2.585678, 3.894531, 4.280472, 5.201035, 6.634384, 5.710678, 
    0.84375, 3.276566, -1.974747, -0.3588562, -1.618744, -0.6388092, 
    -0.2018127, -1.811981, 2.20755, -2.947906, -8.444794, -7.392456, 
    -10.67084, -6.538284, -8.102081, -7.0224, -5.313293, -7.197128, -11.6685, 
    -10.98569, -6.039581, -5.244537, -2.31015, 0.7117157, 0.5049438, 
    2.637756, 2.503387, 0.3403625, -4.756241, -4.342972, -4.587769, 2.412231, 
    4.352615, 12.33775, 10.19635, 11.46094, 0.4268188, 2.599213, 3.275253, 
    1.176041, 0.2486877, -2.165359, -1.216675, -0.5351563, 0.2830658, 
    1.358856, -1.172653, 3.144272,
  1.201035, -0.1929626, -6.791672, -2.373169, -0.9515686, -3.396362, 
    -2.248444, 3.149994, 5.057556, 3.699219, 2.807297, 4.987503, 5.738022, 
    5.830994, 8.361191, 6.413528, 2.077606, 5.756241, 3.48671, 2.227341, 
    2.769791, 5.01329, -2.030472, 6.061462, 5.095581, 5.7164, -0.5817719, 
    -1.478394, 2.545303, 10.36693, 4.563797, -1.958069, -8.321884, -17.51588, 
    -10.89011, -9.067184, -15.99115, -17.49869, -15.28384, -16.48985, 
    -13.02916, -5.209122, 0.2677002, -2.611725, 0.6135406, 4.067444, 
    3.799225, 1.561447, -4.604431, -3.9711, -0.3971252, 3.834381, -0.2901154, 
    -0.7338562, -1.74765, -6.741409, -8.170578, -10.84738, -12.11928, 
    -10.9151, -12.39246, -8.297394, -9.209366, -11.16484, -4.151566, 
    -5.471085, -6.901825, -4.527084, 2.168228, -0.6002655, -1.454681, 
    -0.2861938, -0.0234375, 0.3950653, 3.3685, -0.77005, -7.624481, 
    -5.905991, -7.496872, 0.6062469, 13.87526, 19.71329, 10.02162, 17.05157, 
    14.36328, 2.241928, -2.014313, -7.440094, -1.011719, -5.038025, 
    -3.408859, -5.377609, -1.088547, 0.1440125, -2.125778, -0.5401001,
  -0.3197937, 0.1598969, -2.105469, -1.96199, -4.753647, -4.431519, 1.945313, 
    3.427353, 6.014847, 12.08855, 6.251038, 5.38385, 16.40077, 12.49297, 
    3.802856, 2.860947, 3.378906, 5.963013, 4.626831, 7.71875, 2.067703, 
    -1.710159, 0.6799469, 2.107544, 4.929169, 2.10495, 1.227081, 3.981781, 
    3.502609, 7.137238, -3.882553, -13.4828, -18.1422, -16.07552, -18.8026, 
    -18.3427, -21.64297, -17.52995, -12.99402, -8.638794, -0.7843781, 
    0.002609253, -2.910934, -4.45755, -1.021866, 4.146606, 3.349472, 
    2.245316, 2.140625, -0.06822205, 0.2307281, 1.733337, 5.345306, 1.012512, 
    -3.184891, -8.973434, -13.79713, -9.339584, -3.393478, -7.401825, 
    -9.647659, -4.8862, -3.116409, -1.867447, -4.9888, -0.01223755, 1.040359, 
    -0.9658813, -3.261185, -0.3486938, 2.610413, 0.1359406, 0.9351654, 
    2.009369, 1.786987, -12.50807, -7.161713, -8.410416, -3.329956, 12.25287, 
    17.58621, 13.39427, 5.139847, 9.815369, 23.46172, 6.822922, -3.679413, 
    -9.8797, -7.606247, -6.914841, -4.367188, -1.258331, -3.389069, 
    -4.975006, -4.147385, -2.843231,
  1.300781, -0.1596375, -4.202866, -4.545288, -6.507278, -6.059128, 
    -2.477859, -1.90155, 8.06041, 11.44427, 10.00261, -0.6697845, 3.381256, 
    4.265625, 6.355988, 3.5065, -0.4208374, 4.189056, 2.128647, -2.876312, 
    -10.23412, -7.159378, -2.879425, -1.899994, -0.5645752, 2.384384, 
    0.5846252, 0.453125, 8.86171, 9.783585, -2.759369, -9.913803, -9.542191, 
    -10.45313, -11.65157, -14.78673, -7.289322, -7.199997, -1.359375, 
    6.098694, 5.627075, -0.7260437, -1.168228, 2.783081, 1.62291, 1.753387, 
    5.526566, 4.046356, 4.110168, 6.996353, 9.154419, 6.942978, 5.14035, 
    3.897919, 0.2437592, 2.301559, 1.566147, 2.063797, 4.208847, -2.334381, 
    -0.453125, -1.471863, 7.415115, -1.74765, 0.003646851, 4.098694, 
    3.577347, 3.171875, 4.576828, 7.898178, 1.02449, 1.307297, 1.745056, 
    -0.2966156, 0.7145691, -7.656509, -8.0979, -6.934097, 12.1203, 23.65025, 
    8.707031, 5.926559, 7.157288, 3.633072, 30.19766, 7.063797, -4.162506, 
    -12.8862, -12.92291, -7.686981, -6.070313, -6.335938, -3.188538, 
    -2.084641, 2.910934, -0.9505157,
  7.322922, 5.901031, 1.984634, -3.54895, -3.902863, -2.17865, -1.447388, 
    -0.6338501, 4.891144, 11.82994, 12.37994, -2.569275, 1.853134, 0.2744904, 
    -0.3937531, 1.975525, -4.054169, 0.1609344, -4.932556, -4.738022, 
    -0.7624969, 0.9059906, 2.827332, 5.649734, 4.114319, 1.344528, 3.720047, 
    2.828903, 9.371613, 11.5289, 3.346878, -3.429169, -5.615356, -6.311462, 
    -6.619507, -7.845322, -2.266144, -4.598419, 0.9460907, 6.239594, 
    2.385666, 2.6763, 4.263016, 1.801834, 1.931763, 7.651306, 7.246872, 
    8.071884, 9.371353, 9.932816, 12.47552, 11.73073, 8.896606, 8.188538, 
    5.914322, 6.17395, 6.908859, 7.563538, 3.58046, 2.719788, 7.027603, 
    1.702072, 2.867981, -1.545837, 7.263535, 2.539322, 4.557037, 6.042191, 
    6.540375, 4.377609, 3.219788, 5.182556, 1.290619, -0.7531281, -7.941681, 
    -8.209915, -1.392975, 9.412231, 27.17293, 11.23672, 4.441147, 0.07421875, 
    5.846359, 0.6593933, 18.47447, 12.8875, -4.1073, -5.580719, -10.54375, 
    -6.121613, -8.934891, -4.687241, -2.591156, 1.076813, 7.807022, 7.274734,
  7.755981, 7.307816, 3.489594, -4.345047, -5.332031, -3.405212, -3.586975, 
    -2.758087, -1.541931, 8.745834, 10.61926, 5.939056, 5.984375, 4.043503, 
    2.799484, -0.079422, 1.776306, 2.235413, -0.813797, -2.002853, 4.114319, 
    4.315887, 3.000778, 3.427353, 4.639069, 2.550522, 5.986969, -0.5072937, 
    0.2744751, -0.6557312, 3.656769, 2.280212, -0.2398376, -1.552856, 
    -4.3685, -6.470306, -10.3474, -6.642181, -2.754944, 5.45105, 8.509369, 
    3.735413, 1.965363, 4.071869, 6.382294, 12.17889, 9.581512, 8.431519, 
    8.703644, 9.702347, 9.860413, 6.855209, 3.168228, 4.530472, 3.556503, 
    6.6698, 6.653641, 6.181519, 6.708069, 6.856766, 10.37761, 5.846878, 
    2.815369, 0.2695313, 3.003647, 2.710938, 8.346619, 3.715103, 8.365097, 
    4.595566, 4.989075, 3.815628, 3.383072, -1.432037, -14.66954, -9.761978, 
    20.75339, 15.48932, 0.9278564, 1.208862, 1.972137, -0.4210815, 1.0224, 
    0.1726379, -0.1262817, 3.502869, 3.387756, -8.363022, -1.823425, 
    -2.477341, -0.9752655, 0.1481781, -1.748962, 10.68855, 11.50209, 16.35262,
  7.439316, 3.405197, 2.570053, -1.864059, -4.401825, -4.453644, -3.268219, 
    -4.526825, -4.49765, 1.396362, 15.59818, 12.60364, -0.2585907, 4.101563, 
    4.20755, 5.215363, 3.144257, 2.872665, 4.160934, 6.140625, 6.181778, 
    9.049469, 4.258331, 5.452866, 2.084381, -2.6875, -1.059906, -7.773438, 
    -1.636978, 6.774734, -0.5515747, 6.47319, 4.398956, 1.83725, 2.960403, 
    0.8432312, -16.60104, -10.83359, 0.1611938, 4.103119, 8.282288, 8.770844, 
    8.322922, 11.34297, 8.076569, 10.66069, 14.63152, 13.52316, 14.48125, 
    12.21875, 10.56276, 6.101563, 2.148956, -0.1958466, -0.3903656, 
    -0.07577515, 2.745316, 6.221878, 6.527084, 7.957809, 9.211716, 8.132034, 
    9.976303, 7.210678, 10.24661, 6.41745, 4.085419, 5.621872, 5.74324, 
    4.974472, 6.815369, 7.401306, 2.697647, 4.306259, -10.03568, -8.292465, 
    0.9484253, 3.110153, 3.809631, -1.879425, -0.4046936, 4.517975, 2.025269, 
    3.720551, 0.3442688, -2.186462, 6.843231, 4.138809, 1.887756, -0.552597, 
    0.96875, -4.046356, 5.787491, 7.602615, 10.96146, 17.05522,
  -0.2874908, 4.04895, -1.725006, -6.460678, -10.38957, -3.157028, -2.845062, 
    0.1112061, -9.047134, -7.374741, -3.293747, 13.94948, 12.27344, 5.612762, 
    4.372665, 5.399216, 7.30574, 5.650803, 8.140625, 6.158844, 0.9002686, 
    -1.566406, -1.5578, -0.5255127, 0.9864502, -3.229156, -4.397919, 
    -0.6588593, -4.536209, -5.724487, -13.90862, -10.42552, 10.11328, 
    -1.316666, -3.328918, -2.646088, -8.827866, 5.782043, 3.374741, 
    -1.939575, 3.271362, 6.724228, 5.62265, 1.392441, -7.760666, -9.934128, 
    -15.37604, -15.11537, -15.0724, -13.45651, -12.61197, -10.24167, 
    -4.709381, -4.562775, 0.6236877, 1.89325, 3.904968, 5.924744, 7.897919, 
    8.1828, 5.266418, 4.4552, 4.643494, 7.065613, 6.9758, 5.210419, 6.6922, 
    8.023712, 6.385681, 6.092712, 3.4086, 2.430206, 0.754425, -0.6997375, 
    -5.538803, -0.9622498, 0.6140594, 12.00391, -7.220047, -10.03491, 
    -7.517456, 3.683334, 13.81952, 13.01901, 4.121613, 3.048981, 5.155975, 
    7.313797, -2.341141, -6.117706, -7.469009, -7.592712, -9.273697, 
    -9.510681, -0.4317627, 1.538803,
  -1.039581, -1.389847, -6.092712, -5.698181, -10.62994, -1.271088, 9.967972, 
    11.33698, 6.890625, 2.815887, -3.806519, 7.332031, 13.00053, 2.605194, 
    2.905212, 6.279938, 4.005219, 3.056519, 3.6138, 2.029449, -2.084106, 
    -3.643494, -4.924225, -5.777588, -5.907837, -3.146881, -4.171631, 
    -10.89194, -9.686981, -6.633331, -13.29843, -16.40573, -2.236984, 
    -11.44688, -9.834641, -7.539841, -7.786713, -4.136719, 1.929947, 
    1.859634, 2.357559, 2.611969, -5.128387, -12.05363, -22.925, -27.08385, 
    -31.49635, -32.60103, -28.56616, -25.8867, -24.50078, -21.30389, 
    -15.53723, -12.48047, -6.917969, -3.282562, -0.7333374, 1.057007, 
    1.432281, 1.552612, -0.3005066, 3.123718, 1.099487, 6.78775, 3.167694, 
    1.748169, -0.9140625, 1.327087, 1.242432, -2.091156, -1.692459, 
    -7.689056, -11.14037, -20.50703, -18.08046, -1.666931, -1.233063, 
    -3.677872, -7.789841, -15.2737, 2.199478, 4.634384, 24.10886, 8.485657, 
    14.62111, 19.29401, 19.6974, 3.916931, -6.409378, -7.04895, -10.92995, 
    -8.972137, -8.658081, -10.80417, -6.724472, -6.626831,
  8.164063, 0.8822937, 1.595825, -7.110931, -4.90834, 7.341141, 14.69141, 
    11.5974, 12.98645, 9.904434, 5.135933, 19.49219, 5.196625, 2.575256, 
    2.170563, -1.559113, 2.68515, 2.097137, -1.8078, -2.222122, -7.778381, 
    -8.754425, -6.355988, -13.83907, -9.188782, -4.214325, -1.683075, 
    -9.483078, -8.751312, -9.839325, -13.84323, -11.28229, -12.48932, 
    -7.973709, -5.154678, -2.264847, -4.14505, -1.524216, 6.630463, 7.442444, 
    7.84375, 1.558853, -15.40051, -22.02995, -21.82161, -14.66693, -6.454956, 
    -10.63568, -6.233337, -7.016144, -3.458069, -3.522919, -5.477081, 
    -9.389572, -5.916656, -2.478912, -9.093216, -0.9989624, 5.201035, 
    4.490616, 5.139069, 1.423172, -2.998703, -1.459625, -6.514587, -4.994522, 
    -16.05963, -9.569016, -5.84166, -11.15833, -6.673447, -8.792191, 
    -16.05441, -22.07553, -13.37318, 6.155724, -3.074219, -7.282303, 
    17.00782, 12.98204, 7.993744, 7.4646, 5.863281, 7.351318, 18.29271, 
    12.39272, 12.80754, 0.8846436, -7.178635, -3.226044, 1.720566, 8.072388, 
    8.073425, 3.338028, -3.200516, 2.570572,
  6.767441, 9.955475, 10.05313, 4.671875, 7.773178, 13.8409, 18.16119, 
    9.736465, 17.00835, 17.09584, 15.31485, 11.47916, -4.307556, -5.300781, 
    -4.837738, -12.46484, -10.27527, -5.495575, -5.46666, -8.661987, 
    -6.199738, -8.751816, -16.79871, -15.71432, -2.674225, -3.116928, 
    -6.496872, -8.660416, -5.74324, -6.414581, -11.56328, -10.14168, 
    -10.17448, 1.970047, 1.764587, 5.365891, 8.173691, 6.761459, 10.63905, 
    2.46875, -2.389328, -1.073441, -14.44218, -18.87968, -13.64218, 
    -8.607544, -2.808853, -5.865616, -3.644531, -0.3924408, 5.484375, 
    5.206772, 3.014587, 4.985672, 7.372925, 10.52422, 12.14896, 16.81641, 
    21.02605, 22.46016, 16.19063, 12.0289, 13.76379, 17.75885, 11.31017, 
    19.26588, 17.17552, 13.55937, 15.64764, 24.20078, 14.75833, 9.374222, 
    23.29193, 12.83438, 8.796356, 14.66353, -0.1067657, 15.49089, 14.58438, 
    5.988007, 1.103638, 0.4070129, -0.984375, 2.310181, 0.5021057, -2.482056, 
    2.206512, 1.974213, -0.09191895, 7.625259, 10.17526, 13.31042, 15.69948, 
    9.694534, 11.88646, 3.8974,
  6.802597, 1.131516, -8.839325, -9.79454, -9.282028, -2.4599, 9.193237, 
    20.49895, 11.46327, 10.14297, 17.05493, 7.459381, 0.3286438, -4.901031, 
    -6.757813, -6.401581, -12.85443, -7.078644, -0.2406311, 0.7921906, 
    9.677864, -3.420044, -12.61719, -10.67917, 2.204163, 4.728912, 0.7398376, 
    1.896103, -9.635674, -12.01276, -12.60391, -10.92319, -7.030991, 
    -3.446365, 2.931763, 10.55521, 11.01953, 6.992447, 4.840118, 3.029419, 
    -4.147141, -3.833847, -8.084106, -10.74557, -3.134109, -3.727859, 
    -8.879425, -6, -6.824738, -5.77681, -6.457291, -7.638031, -4.24559, 
    -0.8195343, -0.07240295, -4.720566, -2.910675, -2.2211, 3.250778, 
    4.069016, 6.530457, 12.57552, 13.61954, 12.04688, 11.07683, 15.41902, 
    21.34818, 22.69324, 20.37422, 15.71797, 12.22499, 18.38174, 40.88229, 
    28.95442, 4.146851, -1.051056, -5.496094, -6.988281, -1.957825, 
    -4.417206, 2.208862, -3.06665, 1.114349, -5.875275, -5.391693, -2.894012, 
    -4.314056, -0.8236847, -0.610672, -0.03747559, 4.488037, -2.722916, 
    5.813278, 13.47786, 4.770569, 5.860413,
  -5.536957, -5.777863, -10.0094, -11.51666, -12.04477, -9.078125, -5.314056, 
    -0.02578735, -2.141418, 1.252594, -0.5075684, -3.880463, -4.899231, 
    -8.3302, -10.10547, -7.660156, -0.9335938, -3.873932, -6.101807, 
    7.236969, 8.357292, -2.657028, -0.9523468, -3.900787, 9.1875, 9.140884, 
    6.651306, 5.921875, -8.115891, -26.64479, -12.50833, -2.973175, 2.682281, 
    2.116409, 0.8083344, 10.07005, 5.821365, -1.636459, -2.7724, -5.094788, 
    -2.972916, 1.204422, 0.2549591, -6.038803, -4.997391, 0.0328064, 
    2.460144, -0.09609985, -3.949234, -3.860413, -4.538544, -2.801575, 
    1.933594, 2.150269, 0.7122498, 1.345032, 4.297394, 9.846863, 10.57968, 
    5.01825, 8.259903, 11.84296, 16.45651, 10.00104, 10.49582, 9.767944, 
    10.88617, 5.6091, 9.765625, 15.08751, 28.86171, 44.96173, 44.83098, 
    7.142456, -2.152863, -3.455719, -4.436462, -6.191162, -4.716156, 
    -7.017181, -3.128906, -5.158081, -2.885406, -4.610931, 0.0953064, 
    -2.307297, -2.547653, 3.473434, 3.502869, 7.71875, 0.4671936, -3.145844, 
    6.833069, 3.743744, 0.7291565, -5.040619,
  -3.489349, -2.970306, -5.984894, -5.085938, -5.696106, -5.524475, 
    -3.980988, -5.393494, -4.663818, -4.14505, -5.353912, -6.681274, 
    -8.033051, -11.14166, -10.60104, -8.650787, -6.5177, 1.051544, 2.451324, 
    -2.808594, -4.655197, -7.019272, 4.012756, -0.2054749, 2.935684, 
    13.21588, 7.052605, 9.22448, 2.527863, -6.985413, -8.982544, -11.96432, 
    -3.876831, 3.621613, 5.052353, 6.961975, 7.697388, 3.588806, -6.045822, 
    -10.82213, -3.391663, -0.5304718, -1.339584, 2.309113, -1.941925, 
    0.01405334, -1.17865, 4.70311, 9.226807, 5.174225, -0.0796814, 3.785156, 
    -0.4468689, -3.579163, -4.270309, 0.7463684, 2.897659, 4.593491, 
    9.372665, 8.134369, 11.70261, 11.84088, 9.146088, 9.302094, 8.839294, 
    3.133606, 7.092712, 8.575775, 31.50885, 30.59557, 33.58516, 23.6781, 
    15.27762, -0.9682312, 0.6216125, -4.013031, -0.2252808, 0.8250122, 
    0.2088318, -3.743744, -3.378113, -3.638, -3.039307, -1.101044, 0.1424408, 
    -2.486969, 1.413269, 1.667969, 1.033844, 3.905212, 1.90625, -0.4716187, 
    2.510132, -0.6749878, -3.232269, -3.639832,
  -0.8942871, 6.438538, 0.193512, -2.583862, -2.6297, -3.097137, -3.484375, 
    -3.782562, -4.63205, -5.10025, -5.011993, -5.958344, -6.6987, -9.186707, 
    -13.14038, -13.16431, -14.72867, -22.96378, -24.09583, -23.08125, 
    -14.12787, -13.81328, -11.34634, 0.3924408, 5.891922, -3.789581, 
    -3.080734, 13.36667, 17.04323, 6.191666, 5.944794, 2.614838, 0.8148346, 
    1.092453, 2.78595, 4.073425, 3.181503, 1.581253, -3.422394, 0.7361908, 
    4.603638, 1.96405, 3.246613, 10.86717, 5.214066, 0.8018188, 3.494537, 
    4.3526, 9.655731, 8.302887, 7.993744, 9.505997, 4.351288, -7.402603, 
    -8.920059, -1.465622, -0.4377594, -1.542175, 5.065094, -2.154434, 
    3.391907, 2.884888, -3.27475, -4.257538, 1.869781, -10.70364, 9.950012, 
    15.87943, 25.59322, 1.639328, 9.064575, 0.8346558, -1.97995, -0.4744873, 
    -2.622406, -5.583588, 0.3656311, -3.072906, 0.02578735, -2.296356, 
    -0.3567505, -3.019531, -3.870819, -0.1601563, -1.355469, -4.721619, 
    1.147903, 1.443237, 3.378906, 4.828125, 2.545319, 0.5617065, 1.5466, 
    1.857544, 0.7880249, -1.058319,
  0.8903809, -0.2765503, 0.2098999, -2.842987, -0.5559998, -2.142426, 
    -2.861206, -2.998962, -3.224487, -4.454437, -4.916656, -7.145294, 
    -6.857025, -5.905975, -6.993744, -10.28906, -11.49713, -11.10416, 
    -21.72867, -27.71954, -22.27527, -17.36588, 3.09166, 1.670059, 2.497398, 
    0.5926971, -13.9474, 0.4151001, 17.23828, 10.94426, 12.82085, 14.88672, 
    22.24271, 8.858063, 3.878403, 1.661713, -0.7911377, 1.217438, 1.960144, 
    0.003662109, 0.8465881, 0.0619812, 4.864838, 7.2435, -1.4599, -1.854675, 
    -1.529694, 0.9666443, 4.453644, 7.159637, 5.916656, 10.23126, 9.751831, 
    -2.759399, -6.676819, -6.178131, -0.1411591, 2.782303, 0.1604156, 
    0.4023438, -4.20105, -4.451828, -4.496857, -10.41721, -10.96301, 
    1.285156, 4.084625, 9.546082, 2.632263, -6.406525, -6.49295, -11.53412, 
    -6.329163, -3.654694, 7.217438, 7.215118, 4.427612, 1.519806, 2.76825, 
    3.188049, 2.184631, 0.007049561, -5.146606, -3.159637, -3.043732, 
    -6.22316, -5.291946, -1.282303, 1.913025, 2.255707, 8.198151, -8.702866, 
    -1.658051, 0.8664246, 3.291656, -1.172394,
  3.851044, 6.424469, 6.570313, 1.588287, 0.7179565, 0.7406311, -0.7640686, 
    -2.406769, -3.682037, -2.559906, -4.85965, -4.895813, -4.851807, 
    -5.102081, -7.833862, -9.74115, -6.297119, -5.114563, -2.139038, 
    -9.565887, -14.91901, -19.65729, -14.32031, -17.52734, -8.635422, 
    -4.237244, -10.22421, 2.878906, 30.39922, 18.55937, 0.5049591, 3.065353, 
    3.218216, 2.286438, 1.566925, -1.111176, -3.007538, 1.331238, -4.281769, 
    -1.1716, -1.973175, -4.221893, 0.04348755, -2.093231, -5.27005, -7.1987, 
    -1.682831, -0.6940002, -0.4976501, 1.232574, 4.273193, -1.405731, 
    -4.540375, 6.751038, 6.680725, 0.7007751, -0.5320282, 1.372925, 
    -4.851303, 0.6145782, -3.603638, -6.029144, -12.78751, -24.84113, 
    -4.061188, -0.7153625, -0.83255, 2.661713, -6.175781, -7.266418, -9.9664, 
    -7.769531, -4.605713, -4.321869, 3.685135, -0.8562622, -1.103119, 
    1.117706, 2.879425, 1.528656, 5.004669, 2.236725, 2.824738, 1.142456, 
    0.9765625, -2.129425, -2.752075, 0.9778748, 0.5330811, 2.633331, 0.4375, 
    1.435425, -19.31355, -3.215881, 2.430481, 7.323181,
  5.733856, 13.03906, 16.64844, 10.03699, 0.8401184, -0.8919067, 1.66275, 
    -0.950531, -2.177582, -3.033356, -4.173706, -4.595825, -4.572906, 
    -5.266144, -7.355194, -7.788544, -6.862244, -5.10025, 1.911987, 5.08075, 
    -2.65155, -11.32501, -9.615097, -9.442947, -0.3257751, 5.118225, 
    9.047409, 18.10678, 32.2612, 20.13698, 7.232544, 2.052353, -0.8283844, 
    -10.89818, -5.985413, -9.210938, 1.126312, 6.292969, -8.688278, 
    -9.655457, -10.23647, -5.520325, -2.873947, -0.634903, 1.436203, 
    -3.576553, -1.523178, 1.135422, 3.529434, 2.005203, -2.0289, -5.317184, 
    -4.516144, 2.959625, 4.427612, 5.318481, 4.77005, 3.942963, 4.289856, 
    1.041931, -0.5377502, -3.262756, -10.18124, -7.285156, -7.754944, 
    -3.817169, 1.875244, 0.5664063, 1.089844, -6.583588, -7.5177, -5.224731, 
    -5.175018, -4.098969, -4.296112, -8.431778, -9.036987, -4.132538, 
    -2.203125, 2.103394, -0.7807312, -3.5383, 3.262238, 1.9888, -0.2781372, 
    0.7471313, -4.279144, -1.915863, 0.7416687, 4.633575, -1.148438, 
    0.4825439, -9.198456, -17.54453, -1.926849, 1.463287,
  7.85675, 5.090637, 1.909363, -1.123199, 3.566925, 7.020325, 6.217712, 
    1.78125, 4.804413, 4.893738, -0.2914124, -2.405731, 0.349762, 0.120575, 
    -3.875519, -6.500793, -5.199463, -6.62265, -5.928131, 1.929413, 6.332794, 
    -2.765381, -5.63205, -1.843231, -0.7268066, -0.9570313, 8.449997, 
    20.16197, 18.58855, 17.29297, 18.9948, 12.00885, 3.421616, -3.820572, 
    -10.34479, -9.853134, -6.986191, -2.009888, -7.971085, -6.896103, 
    -8.006516, -8.602859, -6.106781, 0.3507843, 3.433334, 5.746094, 1.129425, 
    1.510162, 5.823441, 3.699997, -1.583847, -0.1158905, 4.529694, 6.30365, 
    3.592453, -0.9028625, 2.192978, 4.315628, 6.702087, 2.027863, 1.498962, 
    -0.701828, -5.526825, -5.457825, -7.248444, -3.760956, -3.690369, 
    -1.936737, 2.608337, -4.171082, -6.147369, -8.922913, -8.414581, 
    -6.757019, -4.397125, -6.757294, -6.597656, -5.905212, -0.2283936, 
    3.632813, 0.3666687, 3.979431, 2.084106, -2.921875, -3.178391, -6.529434, 
    -2.138275, -5.914337, -5.40625, 1.848694, -0.2463379, -3.702332, 
    -0.2330933, -1.693481, -2.347656, -1.329681,
  15.3573, 5.090088, 0.694519, 4.3284, 1.822906, 19.86746, 25.64429, 
    5.628113, 5.293213, 5.211456, 7.703918, 13.89063, 4.965637, -5.512482, 
    -6.471375, -7.125, -6.625519, -5.169525, -4.562225, -3.869781, 1.037506, 
    3.029419, 0.8026123, -2.7453, -3.307312, -6.399994, -3.057556, 2.34375, 
    5.427856, 10.5789, 9.402863, 9.944534, 6.963287, 7.707809, 3.009903, 
    -3.810165, -4.022659, 0.5747375, -1.865097, -5.133331, -11.21614, 
    -14.02422, -8.722137, -10.11771, -9.697144, -1.3638, 0.0473938, 
    -1.014587, 4.091141, 1.9375, -0.02474976, 3.001312, 3.031769, -1.370316, 
    -4.721359, -5.722916, 2.802078, 0.9294281, 0.02449036, 4.155212, 
    5.151566, -6.97084, -0.8031311, 2.776031, 6.014069, -3.712494, -6.857544, 
    -4.372681, -8.876053, -12.04401, -3.380737, -3.9646, -4.505478, 
    -2.094528, 3.166931, 6.778381, 5.996872, 2.463287, 3.919022, 5.891159, 
    0.1158905, 6.15625, 7.417709, 1.835159, 4.29245, -11.59323, -17.12187, 
    -13.06094, -14.40625, -2.793503, -1.804169, -8.559113, -7.361725, 
    5.123962, 5.748444, 9.651825,
  30.11485, 24.88385, 30.77057, 12.75, 2.125259, 9.018234, 4.466141, 
    -1.239319, 5.098938, 6.1297, 6.101044, 7.786957, 8.056244, 2.248962, 
    -3.283081, -3.706512, -4.147125, -6.487244, -3.544006, -2.137238, 
    -0.7807312, 0.7783813, 1.947906, 5.782288, 0.04815674, 4.633057, 
    9.291412, 2.521622, -0.1065216, 1.349487, 0.5940094, 0.5114594, 2.419266, 
    1.228394, -2.637497, -8.373428, -3.661194, -10.96223, -9.687241, 
    -8.919525, -14.07187, -11.21875, -9.133072, -10.93282, -9.809372, 
    -6.219528, -1.571884, -1.707031, -0.02005005, 1.585938, 1.1875, 
    -1.647141, -4.802078, -1.67865, 3.344009, -3.784378, -3.661987, 
    -3.291397, -5.718491, 0.9960938, -1.334366, -7.964325, 0.4593658, 
    6.594269, 16.74843, 6.713013, -5.134644, -6.671356, -8.374481, -4.944275, 
    -2.686722, -1.258865, 2.302597, 1.770844, 1.772919, -3.152863, 2.308594, 
    9.210159, 10.62552, 11.66797, 7.771606, 1.219528, -3.000259, -5.583847, 
    2.131516, -0.2294312, -4.894531, -2.129166, -5.874741, -7.193497, 
    1.993759, 4.564056, -1.378128, -0.06562805, 7.173447, 19.6823,
  18.85338, 21.50104, 15.94844, 0.8528595, -7.284363, -5.416138, -4.154953, 
    -4.827606, -1.580215, -2.43985, -2.88829, -0.9752655, 1.496613, 
    -2.452606, -7.936188, -5.734894, -3.527084, -6.212494, -1.453888, 
    1.646088, -0.8856812, 0.440094, 4.413818, 7.595581, 9.269012, 9.279953, 
    6.248169, -2.922134, -3.224213, -1.846603, -4.837234, -5.092453, 
    -4.134628, -6.932816, -8.491653, -12.02812, -11.20105, -9.943741, 
    -9.770569, -9.640366, -4.044022, -0.1177063, -5.418228, -10.12057, 
    -6.913544, -4.926559, -1.346359, 0.2177124, -0.5223999, -2.444, 
    0.4729309, 0.2932281, -4.424225, -6.951813, -2.896881, -0.9291687, 
    0.9554749, 3.101822, -1.76535, -4.524475, -3.4888, 5.3349, 15.09792, 
    21.81615, 20.71223, 12.75156, 5.886978, 6.68074, 3.870575, 3.977081, 
    3.257553, 3.420822, 4.753387, 3.694794, 2.769012, 5.430466, 8.029434, 
    3.27005, 5.963287, 10.37578, 6.522659, 4.386993, 2.33905, 2.568222, 
    2.89296, 1.313293, -1.435944, -5.599991, -8.9039, -3.724747, -3.233582, 
    -4.047394, -0.3716125, -0.8549347, 0.5802002, 9.630203,
  9.129425, -0.0526123, 1.483078, 2.965103, 1.866409, 2.985947, -2.004684, 
    -14.03438, -18.09792, -19.24739, -17.6815, -13.05782, -5.318481, 
    -9.496353, -12.8349, -13.79166, -10.33073, -6.403915, -5.810425, 
    -7.717972, -1.507553, 4.222656, 2.548172, 3.161972, 3.595322, -1.4263, 
    -4.270065, -6.021362, 0.5187531, 3.651306, -1.326309, -6.404694, 
    -4.685669, -6.154953, -11.18958, -9.763535, -7.472397, -4.132034, 
    -9.878372, -8.626297, -3.029175, -2.18985, -1.030991, -6.1362, -8.589066, 
    -12.21225, -10.73724, -2.916672, -0.2039032, -0.3184814, 0.1458435, 
    3.154953, 2.444794, -0.2752533, -1.633072, -2.773697, -0.8328247, 
    2.746094, 1.989334, -2.558075, -0.822403, 5.806259, 1.536201, 3.191406, 
    1.752342, 5.402603, 10.64348, 10.77161, 9.852081, 10.88698, 11.12708, 
    8.907043, 5.103378, -0.7166595, -3.486725, -13.52501, -9.239059, 
    -4.373947, -1.049744, -0.691925, -2.657547, -5.986191, -1.5914, 
    0.7945251, -8.450012, -7.639832, -0.6877594, -2.84819, -6.744003, 
    -2.919525, -1.218491, -5.526031, -7.669266, -5.2276, -0.524231, 6.792709,
  -8.415619, -6.377594, -4.053391, 1.136719, 0.1190033, -1.25235, -5.49556, 
    -6.756256, -14.25286, -11.55885, -17.43906, -22.07266, -24.61458, 
    -23.7224, -18.94218, -16.075, -14.2151, -11.25494, -7.072144, -6.584381, 
    -5.5625, -4.849213, -7.752869, -6.372147, 0.3085938, 2.051559, -1.46666, 
    -6.6539, -4.334381, -1.684387, 0.1283875, -0.8796844, -3.794785, 
    -4.976303, -8.293503, -5.471085, 0.1242218, -0.2989502, -6.436722, 
    -7.265366, -8.766159, -9.384644, -6.340103, -4.240364, -4.379166, 
    -1.422913, 1.092178, 3.851303, 4.862244, 4.670319, 3.312241, -3.317963, 
    -2.853912, 3.050781, 6.898956, -0.6747284, -3.3974, -1.422134, 2.354172, 
    1.864334, 1.199219, 2.107033, 4.596359, 1.834892, -4.123688, -5.703644, 
    -2.110672, 2.625534, -1.066925, -3.233856, -6.46875, -4.411453, 
    -11.59375, -15.39246, -8.416138, -4.845566, -2.873962, -8.549484, 
    -12.63776, -12.32786, -5.259888, -3.452606, -1.521362, -4.841934, 
    -8.482285, -5.257034, -1.223434, 1.652344, -2.423172, -2.785934, 
    -2.690887, -4.788544, -8.948166, -9.940628, -4.945053, -4.429428,
  -9.603912, -7.743484, -1.052605, -0.5945282, -3.616409, -8.971359, 
    -8.032806, -7.021881, -8.63932, -7.468491, -10.86953, -13.90547, 
    -11.43959, -10.32944, -6.626297, -4.017975, -3.930481, -3.626572, 
    -3.319778, 0.3817596, 5.623703, 3.101303, 3.897659, 1.739334, 2.797668, 
    -0.795578, 1.373184, -1.183594, -2.125, -1.464325, 1.137772, 4.51796, 
    3.257553, -0.3599091, -6.191925, -6.877869, -9.45079, -4.818748, 
    -3.677864, -4.926048, -3.502861, 0.4286499, 0.1877594, -0.6846313, 
    4.969009, 9.007813, 2.661461, -8.139328, -7.672394, -2.022125, 2.543228, 
    5.207291, 5.380211, 7.509369, 6.476822, 1.749214, -4.97422, -4.851303, 
    -2.84375, -0.6348953, -0.08776093, 6.205727, 6.341408, -3.300003, 
    -9.913284, -10.67526, -7.835159, -5.821869, -4.038284, -2.745056, 
    -6.982803, -8.653397, -8.8573, -7.625259, -10.70677, -14.83932, 
    -14.28724, -11.13229, -11.03671, -9.184372, -7.738541, -11.99739, 
    -13.06902, -7.332291, -5.541397, -12.29218, -17.52421, -12.76485, 
    -5.077087, 0.1911469, 1.460159, -2.26796, -7.191925, -7.464844, 
    -5.119278, -6.178894,
  -17.68776, -19.65, -10.75574, -3.760162, -1.5737, -1.111198, -4.908333, 
    0.1388016, -1.434113, -5.004425, -3.612244, -8.170052, -12.20365, 
    -13.0539, -12.99193, -6.177345, -1.553902, -0.1380157, -2.116669, 
    -1.806511, -5.14505, -5.344788, -10.36771, -14.13879, -13.01875, 
    -11.6763, -10.19167, -4.512505, 0.1773453, -0.4809952, -1.093491, 
    -1.161209, -4.853653, -6.627869, -7.680466, -7.878654, -7.353127, 
    -2.556511, -5.997917, -7.092712, -2.91198, 1.87812, 1.197655, -1.449478, 
    -0.03307343, 2.404427, 4.271614, 0.775528, -6.649223, -4.103386, 
    -0.07682037, -1.299477, 0.1984329, 0.3351517, 2.208069, 4.673958, 
    3.367973, 3.495049, 4.316406, -0.1151047, -3.344009, 0.654686, 5.427864, 
    4.712234, -2.470055, -10.31615, -13.85182, -12.72292, -11.06719, 
    -11.84192, -9.097916, -8.913017, -4.340363, -2.656509, -12.47735, 
    -11.04219, -12.2112, -10.06068, -8.241669, -10.08568, -14.61015, 
    -16.60651, -15.60078, -11.3466, -10.28384, -10.13646, -12.95703, 
    -13.89037, -11.08047, -8.633331, -8.0112, -3.120316, -2.361465, 
    -0.4395905, -2.263809, -9.35833,
  -3.691147, -4.2724, -4.015106, -5.820831, -7.655991, -2.942451, -1.775787, 
    -4.153908, -2.217445, -0.006767273, -0.4145889, -5.745056, -10.48776, 
    -12.58932, -11.24088, -10.10911, -7.303123, -6.734375, -7.045578, 
    -6.855988, -3.461197, -2.819794, -2.615372, -6.155212, -7.553909, 
    -2.99427, -4.990364, -6.771095, -4.767189, 0.8643188, 4.836197, 7.269531, 
    5.146873, -0.2911453, -5.734375, -5.521614, -4.529427, -4.504433, 
    -6.595833, -9.313019, -12.07343, -14.93281, -15.90234, -14.89948, 
    -13.93463, -12.25833, -8.59687, -5.790886, -5.609375, -13.41068, 
    -6.126823, -7.067451, -9.961723, -4.386978, -3.27005, -3.29557, 
    -3.140106, -2.747658, -3.831512, -6.055725, -8.521873, -9.613541, 
    -8.377342, -5.859634, -7.408852, -10.80052, -9.988541, -6.501305, 
    -2.995834, -3.542694, -0.8507843, 0.673172, -0.0783844, -2.851563, 
    -5.670319, -15.59792, -11.07813, -10.40365, -11.43047, -15.46616, 
    -12.70442, -11.51927, -12.6987, -12.44479, -9.973694, -9.827866, 
    -9.137756, -9.312759, -11.78307, -13.17162, -11.54844, -10.92656, 
    -10.17838, -4.308075, -2.43541, -2.120056,
  -4.271355, -1.678383, -0.3289032, -1.146614, -4.671097, -7.084373, 
    -11.80183, -16.18464, -15.29766, -11.35313, -7.720055, -5.359375, 
    -5.541672, -6.523697, -8.24192, -9.708595, -20.80547, -19.39088, 
    -19.03958, -13.44505, -12.67162, -12.26563, -13.10755, -12.2651, 
    -9.938805, -5.753387, -1.004166, 1.527344, 3.625, 7.077339, 7.529167, 
    4.475525, 1.190102, -0.54245, -0.6671906, -4.216927, -3.862503, 
    -3.450783, -4.49427, -8.957558, -13.89922, -12.74114, -10.35209, 
    -8.871613, -9.150253, -11.1151, -12.02525, -12.96537, -14.35313, 
    -14.63698, -14.34635, -15.57135, -16.17317, -14.99375, -13.89896, 
    -13.48438, -16.00365, -18.3401, -18.28645, -16.12187, -12.88359, 
    -11.18098, -10.99974, -6.32708, -6.219269, -5.134895, -2.211723, 
    -2.196358, -3.795052, -6.612762, -9.196617, -12.42057, -13.91146, 
    -11.23985, -9.039581, -9.964584, -8.69323, -18.55964, -15.80859, 
    -11.51668, -7.923447, -5.352859, -5.296341, -4.189331, -4.227081, 
    -6.678909, -9.275269, -6.950531, -5.150513, -5.371094, -7.492981, 
    -7.572647, -3.319527, -3.396095, -4.752609, -5.393227,
  -7.799225, -8.404686, -8.183853, -7.556511, -4.900261, -3.067192, 
    -3.257294, -5.812241, -6.372917, -7.283333, -8.442184, -10.09322, 
    -10.19245, -11.42136, -12.43177, -12.71146, -11.95625, -11.43229, 
    -10.23932, -10.32995, -11.03125, -12.15234, -12.53958, -12.14063, 
    -10.39948, -4.742714, -1.851036, 1.539063, 3.564064, 3.014587, 
    -0.4463577, -9.960678, -11.6125, -11.18932, -10.74454, -8.7901, 
    -6.743492, -7.036194, -7.296097, -8.595055, -12.17838, -12.82604, 
    -11.66693, -10.52579, -9.220573, -8.316147, -8.069794, -9.586456, 
    -12.64063, -15.29765, -16.10963, -15.10313, -13.55677, -12.07369, 
    -10.47709, -9.098694, -9.219528, -10.41458, -13.0711, -14.63516, 
    -16.17474, -17.26979, -19.98776, -22.38359, -26.36875, -17.03073, 
    -17.73074, -17.31068, -17.28672, -17.10078, -17.93021, -15.21875, 
    -12.32917, -8.369011, -7.290108, -18.88541, -19.83438, -14.93359, 
    -10.72084, -11.17319, -10.13152, -8.507034, -6.357803, -2.501312, 
    0.9460907, -1.738022, -6.573441, -8.205215, -8.001312, -7.169006, 
    -5.7388, -9.946869, -16.12526, -11.70755, -7.501564, -7.112244,
  -12.2513, -14.23073, -14.5862, -16.21041, -11.4776, -11.15443, -9.848961, 
    -18.36302, -19.075, -18.619, -16.88281, -15.08749, -15.03464, -13.9888, 
    -12.6763, -12.60755, -12.1375, -11.71953, -12.9474, -14.19297, -14.29948, 
    -14.30286, -11.92422, -9.141663, -5.814064, 1.167969, 3.734894, 
    -4.433334, -4.057297, -6.488281, -8.797913, -9.827087, -10.43281, 
    -10.35078, -9.748436, -9.655472, -9.143753, -8.964584, -8.808853, 
    -9.460159, -9.72995, -10.33828, -10.88932, -11.05885, -11.66198, 
    -11.0276, -10.2474, -9.953644, -10.20573, -10.9586, -12.24974, -13.9185, 
    -13.48854, -12.4862, -12.01719, -12.37292, -12.96015, -12.56015, 
    -11.44609, -10.55729, -9.62838, -10.33776, -11.56172, -13.21667, 
    -14.82474, -15.11458, -15.08803, -13.73099, -12.19896, -9.983589, 
    -7.875259, -0.6424408, -3.209373, -0.2028656, -1.498962, -2.095566, 
    -2.83046, -2.774734, -2.916656, -3.876053, -3.414581, -3.375778, 
    -2.814056, -3.110687, -4.839844, -8.066147, -10.51563, -11.30521, 
    -11.31198, -10.55208, -11.20599, -13.34088, -20.52969, -19.02422, 
    -14.35703, -12.77917,
  -11.3526, -10.96016, -11.18906, -11.3763, -11.8263, -11.67657, -10.91744, 
    -9.850266, -8.760933, -7.670578, -7.633598, -7.989586, -8.42057, 
    -8.019012, -7.66198, -6.784897, -5.991142, -5.669533, -5.52578, 
    -5.822136, -5.884377, -5.587761, -5.290627, -5.334892, -5.100777, 
    -4.679947, -4.021347, -3.796349, -4.524223, -5.761986, -6.936455, 
    -8.365097, -9.841667, -10.93463, -11.66589, -11.96953, -12.12734, 
    -11.87526, -11.34088, -10.47447, -9.019791, -7.570053, -6.783852, 
    -6.805725, -6.764587, -7.38073, -7.924477, -8.560936, -9.911201, 
    -11.87605, -13.57317, -14.81224, -15.79219, -16.32057, -16.62031, 
    -16.13854, -15.39427, -14.52161, -14.24088, -13.75885, -13.46068, 
    -14.07265, -14.50105, -15.25521, -16.00417, -17.2875, -18.30469, 
    -18.48203, -18.67084, -18.98021, -19.33541, -19.80807, -19.5375, 
    -17.70808, -16.09557, -14.79011, -14.20052, -12.45103, -10.89792, 
    -10.1388, -9.538284, -9.273705, -9.369019, -9.738281, -10.53073, 
    -12.01459, -14.34557, -15.56509, -16.1763, -16.8336, -16.66171, -16.6625, 
    -15.90652, -14.89662, -13.45625, -12.28099,
  -15.13047, -15.5461, -16.11459, -16.52631, -16.81536, -17.12969, -17.22292, 
    -17.12474, -17.01276, -16.90417, -16.62813, -16.19505, -15.61849, 
    -14.83828, -14.03698, -13.20495, -12.17057, -11.37917, -10.76719, 
    -10.30756, -10.07005, -9.730209, -9.200523, -8.89193, -8.596359, 
    -8.252602, -7.9263, -7.595573, -7.387238, -7.234634, -7.163277, 
    -6.964058, -6.615364, -6.244537, -5.9888, -5.732292, -5.348961, 
    -5.059372, -4.601303, -4.348175, -4.370049, -4.547913, -4.780464, 
    -4.914589, -4.954163, -5.067444, -5.299736, -5.759369, -6.124481, 
    -6.453903, -6.560677, -6.381775, -6.345573, -6.434113, -6.329163, 
    -6.092453, -5.563805, -5.216927, -4.680725, -4.312759, -3.950256, 
    -3.727867, -3.453125, -3.167709, -2.754951, -2.639587, -2.642967, 
    -2.547653, -2.54792, -2.509636, -2.647919, -2.651306, -2.640106, 
    -2.438797, -2.179428, -2.222656, -2.331772, -2.373955, -2.445572, 
    -2.568748, -2.829948, -3.571617, -4.064583, -4.767967, -5.522133, 
    -6.239067, -6.822136, -7.631508, -8.741669, -9.498962, -10.37161, 
    -11.35963, -12.30911, -13.15417, -13.85365, -14.61015,
  -0.02099609, -0.0108397, -0.01266265, -0.01682949, -0.02203774, 
    -0.02672529, -0.03505874, -0.0577147, -0.07594395, -0.1157877, 
    -0.1486003, -0.1691732, -0.1926105, -0.227246, -0.242871, -0.2454753, 
    -0.257715, -0.264746, -0.2788086, -0.2834961, -0.2696941, -0.2657878, 
    -0.2728188, -0.2866211, -0.2887044, -0.2933919, -0.3012044, -0.3025064, 
    -0.2996418, -0.2933919, -0.2931316, -0.2980795, -0.2996418, -0.3014648, 
    -0.3084962, -0.321517, -0.3272462, -0.334017, -0.3433919, -0.3584962, 
    -0.3707356, -0.3816731, -0.3884439, -0.3905275, -0.3874023, -0.382194, 
    -0.3749025, -0.3691733, -0.3579752, -0.3600588, -0.3558915, -0.3532872, 
    -0.3431306, -0.3444326, -0.3394847, -0.3303702, -0.3233387, -0.3282869, 
    -0.341568, -0.3613596, -0.3660471, -0.3790681, -0.3954742, -0.402245, 
    -0.4142249, -0.4173496, -0.4191725, -0.4230788, -0.4202142, -0.4155269, 
    -0.4058914, -0.3983395, -0.3845372, -0.3616207, -0.3470373, -0.3376622, 
    -0.3379226, -0.3314123, -0.3178706, -0.2985997, -0.2780268, -0.2566726, 
    -0.2295897, -0.2124023, -0.1915689, -0.1920898, -0.1842773, -0.1884439, 
    -0.17959, -0.1754231, -0.1538086, -0.1342773, -0.1207356, -0.1014647, 
    -0.07724595, -0.04052734,
  0.325881, 0.2545271, 0.1753597, 0.1019249, 0.06728935, 0.03759956, 
    -0.01969147, -0.06213951, -0.1170874, -0.1556311, -0.220211, -0.3077126, 
    -0.3722954, -0.4439096, -0.4652643, -0.5259409, -0.5821896, -0.6387005, 
    -0.65693, -0.6587524, -0.7017212, -0.755888, -0.823597, -0.8803673, 
    -0.922555, -0.9639606, -1.00146, -1.021253, -1.005888, -0.9571896, 
    -0.9150019, -0.872035, -0.7910452, -0.7163057, -0.7069311, -0.7488565, 
    -0.8209915, -0.8488569, -0.8454733, -0.8449526, -0.9079742, -0.9441729, 
    -0.9631824, -0.9808884, -0.9259415, -0.8866205, -0.8014641, -0.7332344, 
    -0.5957355, -0.53584, -0.5332365, -0.5446949, -0.5449538, -0.4650059, 
    -0.3652668, -0.3262038, -0.3314137, -0.35537, -0.3600588, -0.2506847, 
    -0.1834965, -0.1808915, -0.2280269, -0.3642244, -0.4767251, -0.6090164, 
    -0.7571945, -0.8793302, -0.9202151, -0.8587556, -0.718132, -0.7043295, 
    -0.6814132, -0.6665697, -0.6608405, -0.5918298, -0.5803709, -0.5470381, 
    -0.5314131, -0.5530276, -0.5486007, -0.4329758, -0.2618809, -0.1217766, 
    0.04645252, 0.2394209, 0.4133792, 0.5727539, 0.6365561, 0.6373367, 
    0.6636391, 0.6344728, 0.5581703, 0.5136404, 0.4795256, 0.3990564,
  -0.1525078, -0.1314144, -0.1926136, -0.3436546, -0.4751644, -0.5626659, 
    -0.6170921, -0.7816753, -0.8512096, -0.9907932, -1.082458, -1.185844, 
    -1.259541, -1.331417, -1.361624, -1.396259, -1.372562, -1.257198, 
    -1.100166, -1.00824, -0.9308968, -0.9124069, -0.9605827, -1.049906, 
    -1.15173, -1.266573, -1.290272, -1.323605, -1.346783, -1.322042, 
    -1.307198, -1.335321, -1.393396, -1.49626, -1.583759, -1.554853, 
    -1.573866, -1.522301, -1.411886, -1.405115, -1.43376, -1.51918, 
    -1.664228, -1.827511, -1.909283, -1.811626, -1.616312, -1.451727, 
    -1.392612, -1.106415, -1.025946, -1.084278, -1.245996, -1.343131, 
    -1.576466, -1.65329, -1.615269, -1.413446, -1.455635, -1.323082, 
    -1.224123, -1.102251, -1.154593, -1.326206, -1.687661, -1.967608, 
    -2.231931, -2.310838, -2.19313, -1.834795, -1.182714, -0.7230759, 
    -0.7280254, -0.5941715, -0.4696941, -0.2394867, -0.1241207, -0.08323574, 
    -0.3741236, -0.6462584, -0.9095402, -0.9491234, -0.6686535, -0.3733406, 
    -0.1100597, 0.05817127, 0.1115561, 0.1875973, 0.4386387, 0.5667648, 
    0.5917625, 0.5055637, 0.1987896, -0.04756737, -0.2139683, -0.2556362,
  -1.360313, -1.416306, -1.426464, -1.379848, -1.393654, -1.364742, 
    -1.487659, -1.518391, -1.41188, -1.31839, -1.451725, -1.671257, 
    -1.762138, -1.834274, -1.780369, -1.804329, -1.892612, -1.768913, 
    -1.727245, -1.57959, -1.309799, -1.150421, -1.044952, -0.9853134, 
    -1.096519, -1.31292, -1.633755, -1.756672, -1.616833, -1.515266, 
    -1.518654, -1.461357, -1.601204, -1.699379, -1.654064, -1.473858, 
    -1.310314, -1.199116, -1.362663, -1.373341, -1.250938, -1.31292, 
    -1.178806, -1.005627, -1.118389, -1.60667, -1.990261, -1.91787, 
    -1.805367, -2.025681, -2.245995, -2.205891, -1.951723, -2.096514, 
    -2.619432, -2.882713, -2.775948, -2.738449, -3.043137, -2.729855, 
    -2.122564, -1.965271, -2.048864, -2.324905, -2.708241, -3.204334, 
    -3.660843, -3.466574, -3.08923, -2.894438, -2.775427, -2.791313, -2.3335, 
    -2.211624, -2.154072, -1.844177, -1.587667, -1.846785, -1.718397, 
    -1.717875, -2.074905, -2.198084, -2.220739, -2.144436, -2.086102, 
    -2.097822, -2.032454, -1.858234, -1.491827, -1.268133, -1.355894, 
    -1.604588, -1.859013, -1.782711, -1.556927, -1.426205,
  -1.737408, -1.956944, -1.650955, -1.667099, -1.756683, -2.21814, -2.657467, 
    -3.131687, -3.548092, -3.491318, -3.252777, -2.807461, -2.716316, 
    -2.590275, -2.283245, -1.899128, -2.011627, -2.432465, -2.233246, 
    -1.900692, -1.89262, -1.854858, -2.503815, -2.574909, -2.426212, 
    -2.369442, -2.372307, -2.174648, -2.076477, -2.169701, -2.322826, 
    -1.99939, -2.168137, -2.589233, -2.884285, -2.826733, -2.588451, 
    -1.96085, -1.26762, -1.212669, -1.297829, -1.166058, -1.10434, -1.091579, 
    -1.078819, -0.2374077, 0.3383713, -0.07907104, -0.3118858, -1.026466, 
    -2.042618, -2.987667, -3.607197, -2.880634, -2.700161, -3.238701, 
    -3.540264, -4.087399, -4.496254, -4.650158, -4.204586, -3.970474, 
    -3.681412, -4.073082, -4.102768, -3.550423, -2.911362, -2.677505, 
    -1.824123, -0.6991158, -0.5866184, -2.146519, -3.038181, -3.128029, 
    -2.538181, -2.206413, -1.428543, -1.214222, -1.244949, -1.761875, 
    -2.356934, -2.700684, -3.222557, -3.083237, -3.285839, -2.953289, 
    -2.885056, -3.089481, -3.275684, -2.998333, -3.201462, -3.185055, 
    -2.916832, -2.638443, -2.200165, -1.595222,
  -1.560593, -1.068161, -0.02412415, -0.620491, -0.6040802, -1.448349, 
    -3.486893, -4.643665, -5.790279, -5.245228, -3.816578, -3.761883, 
    -4.462936, -4.51606, -4.718407, -4.415543, -3.798615, -3.42543, 
    -2.630127, -3.088982, -3.129868, -2.753304, -2.536636, -2.277, -2.647575, 
    -3.421532, -3.31945, -2.8507, -3.235596, -4.201996, -4.605644, -3.735073, 
    -2.023876, -2.087154, -2.892365, -3.316841, -3.21553, -2.718662, 
    -1.649391, -1.28429, -1.779083, -1.926208, -2.325951, -1.081161, 
    -0.003040314, -0.03168488, -1.522568, -1.953033, -2.59444, -3.200172, 
    -3.953297, -3.771008, -3.731419, -4.266319, -4.358501, -4.276733, 
    -4.449913, -5.063454, -6.262413, -6.44809, -6.349915, -5.144447, 
    -4.251999, -3.155384, -2.438713, -1.465275, -0.7582436, -0.5509529, 
    -1.4184, -1.602512, -2.211887, -2.340534, -1.783764, -1.599915, 
    -2.235847, -3.232979, -2.451988, -0.6915779, 0.6430664, 0.1271782, 
    -0.3988686, -0.5980835, -0.8605804, -0.07725525, -0.5543404, -1.974911, 
    -4.2822, -6.124908, -5.872307, -4.918137, -4.906677, -4.962677, 
    -5.204861, -4.548866, -2.296009, -1.341583,
  -7.571007, -6.263191, -4.929588, -4.706169, -4.264244, -4.132477, 
    -2.491066, -2.829346, -3.132217, -4.146011, -4.934296, -4.821014, 
    -6.66346, -7.346016, -6.075699, -5.198616, -4.747574, -5.896538, 
    -7.849136, -8.085075, -5.840019, -3.822311, -2.999657, -3.068665, 
    -2.810593, -2.798615, -2.978043, -2.679085, -3.078568, -2.260071, 
    -2.016327, -1.518669, -0.9868927, -2.313454, -3.017097, -3.711891, 
    -3.948601, -3.528824, -3.33559, -3.504082, -5.218666, -6.159554, 
    -6.344707, -4.917107, -3.170746, -4.706425, -6.492626, -6.98872, 
    -6.913986, -4.89653, -2.635075, -1.894707, -1.952263, -2.466843, 
    -3.602524, -4.440285, -4.943924, -4.426727, -3.800964, -4.793144, 
    -5.153557, -4.606171, -4.097572, -3.90799, -6.23299, -5.804611, 
    -4.612411, -3.802513, -4.669701, -5.303043, -6.622311, -7.202, -6.041843, 
    -6.1908, -5.811111, -6.058514, -5.965023, -5.209808, -3.67543, -1.868935, 
    -2.992104, -4.676476, -4.904079, -3.68351, -3.198097, -3.50877, 
    -6.554867, -6.423359, -5.676735, -5.633507, -6.169701, -7.197048, 
    -8.385853, -8.126213, -6.872314, -6.767105,
  -4.238968, -2.611885, -1.936104, -2.357452, -4.463959, -5.619171, 
    -4.939751, -4.958244, -3.928299, -6.113441, -7.038971, -5.268402, 
    -4.929077, -6.172577, -7.515541, -8.631432, -8.827515, -8.576469, 
    -6.919693, -5.552254, -5.168137, -6.915794, -7.504333, -6.402763, 
    -4.930115, -2.921005, -2.510582, -3.987923, -4.049393, -2.832726, 
    -0.3707504, -2.387421, -2.797836, -4.029335, -4.835594, -6.162933, 
    -5.983253, -3.122841, -5.401482, -6.620232, -8.060593, -9.308762, 
    -9.84288, -10.22934, -8.926472, -7.570232, -5.713455, -2.405388, 
    -0.5801392, 1.358673, 2.000351, 1.345657, 1.174828, 1.770126, 1.615448, 
    0.1758575, -1.090546, -2.469193, -3.084557, -2.160072, -2.93898, 
    -5.474136, -6.723358, -5.224136, -7.807213, -9.093147, -7.764244, 
    -6.061623, -7.022831, -6.835335, -5.938972, -7.268135, -9.423862, 
    -10.50303, -8.454338, -8.727768, -8.452515, -7.607727, -7.841846, 
    -8.36866, -9.117104, -11.27805, -8.060852, -5.394188, -5.07074, 
    -5.467369, -6.076744, -3.80851, -5.128548, -7.754082, -9.714241, 
    -8.840019, -7.301735, -6.330376, -6.706947, -6.399399,
  -6.641327, -9.126991, -8.824654, -9.875702, -12.2481, -12.8546, -11.37154, 
    -10.02232, -11.23168, -12.88896, -10.38401, -10.14365, -10.29964, 
    -12.48532, -13.95382, -14.44262, -17.21086, -17.43012, -16.3197, 
    -13.63091, -13.94367, -13.02856, -10.47388, -6.261116, -3.604866, 
    -3.613457, -4.117622, -5.207207, -5.610062, -4.483238, -2.490028, 
    0.06283569, 0.7224731, 0.6597137, -0.9967957, -3.023613, -5.648094, 
    -5.919968, -5.890282, -5.71476, -5.462158, -2.978569, -3.447838, 
    -3.188202, -2.702003, -2.226479, -0.5652847, 1.15139, -0.3298645, 
    -1.334816, -2.025703, -2.416061, -1.424919, -0.475441, -1.150696, 
    -0.5428925, -3.131157, -3.321533, -2.630653, -1.324135, -2.251205, 
    -2.779861, -0.7090302, -1.310066, -2.348091, -3.468666, -2.732994, 
    -0.2616425, -1.56424, -2.050179, -2.015541, -2.520493, -3.708511, 
    -3.34211, -2.090546, -1.887413, -3.38221, -2.287674, -2.192368, 
    -2.592621, -2.392883, -2.838722, -1.684555, -5.744965, -8.287659, 
    -10.37074, -9.827255, -6.600174, -6.181427, -7.188461, -6.809036, 
    -6.0783, -8.697044, -9.394974, -9.596535, -6.752266,
  -10.71658, -13.00929, -11.533, -8.581421, -6.594711, -7.390282, -7.1231, 
    -6.106171, -6.134293, -4.732475, -5.324135, -5.518929, -5.96814, 
    -4.481155, -4.456421, -5.50148, -4.212677, -2.504868, -4.687416, 
    -10.5494, -14.70331, -12.57752, -7.304611, -5.782471, -3.47023, 
    -1.508255, -2.094963, -2.560326, -1.669441, -0.7837601, -1.615273, 
    -1.169441, -0.01371002, -1.294434, -2.760056, -3.276733, -2.342102, 
    -1.533241, 1.545403, -0.004859924, -0.3280334, -2.425957, -3.91684, 
    -5.904861, -0.05433655, 2.770142, 2.548782, 0.1980057, 0.8097305, 
    0.8365479, -1.810593, -1.016579, 0.2584229, -1.519196, -0.1967773, 
    0.6972198, 0.9662323, 3.151398, 3.206863, 2.763893, 1.766235, 1.687065, 
    -1.876472, -2.224648, 3.944366, 3.881592, -0.773613, -2.082207, 
    -0.1996536, 0.973526, -1.410591, -3.632988, -5.576485, -3.973099, 
    -1.884285, -2.700432, -5.869705, -8.459297, -3.578049, -0.6618958, 
    1.129242, 0.9313431, 0.6990585, -3.400948, -6.571793, -5.551743, 
    -6.423874, -8.360596, -10.17831, -11.46815, -14.11632, -14.98898, 
    -13.70747, -12.83898, -10.03403, -9.504601,
  -3.72596, -3.595482, -2.181419, -1.772575, -2.971008, -1.852783, 0.3677979, 
    2.389938, -0.7512207, -3.231949, -2.536102, -0.961113, 2.319099, 
    2.086029, -3.015015, -3.027252, -3.757202, -1.826729, -1.599129, 
    -1.39444, -0.2993927, -1.527779, -3.746521, -1.810333, 1.396957, 
    2.992271, 3.23394, 2.776909, 0.3985214, 0.7456512, -0.4267426, -0.322319, 
    1.378212, 1.248009, -1.499397, -1.142357, -2.231689, -1.310593, 
    -0.2796021, 2.025352, -0.5017471, -2.042107, -0.05304718, -3.006424, 
    -1.252525, 2.350868, 2.498795, 0.5206604, -0.3131866, 1.164146, 
    0.4024353, 3.932899, 2.723785, 0.7076416, 2.25634, 0.487854, -1.296524, 
    -0.6496506, 3.030815, 0.1873322, -2.194443, 3.007118, 0.07873535, 
    -1.780899, 4.956078, 5.312325, 0.5589447, -2.777, 1.676384, 0.9951401, 
    -1.176476, -2.104599, -1.7994, 1.852173, 2.249046, -3.281944, -8.996796, 
    -4.909554, 0.0612793, 0.1732635, 3.963104, 3.600868, 3.515976, 3.823265, 
    -0.9246445, 0.2933197, 2.991493, 2.034988, 2.132645, 0.8745728, 
    -5.205894, -5.051216, 0.269104, 2.524307, -1.583771, -3.890549,
  1.411804, 1.007385, -1.757469, -1.508499, 0.5539856, 2.422478, 2.185242, 
    0.6813354, -2.656952, -1.602264, -0.743927, -0.8501892, -0.7311554, 
    -1.388725, -0.5715332, -1.112671, -3.859283, -5.048355, -1.199638, 
    -2.040802, -0.762146, -0.8678741, -5.381157, -0.7595367, 3.593582, 
    0.5277023, 3.780304, 6.39151, 1.940201, 1.814163, 1.535774, 1.037079, 
    6.312065, 6.192024, 2.203476, 2.681854, 4.009727, 3.946442, 2.516762, 
    4.758163, 2.062057, -4.328308, -1.087158, -0.2470551, 2.201645, 3.157646, 
    2.956589, 5.72171, 4.381851, 0.2443542, 1.046707, 6.270653, 6.559464, 
    1.310501, -0.492363, -0.9105911, -5.368668, 1.32692, 2.163643, -1.139755, 
    -1.350418, 1.552696, 2.260773, 3.842285, 2.731071, 1.15242, 0.6649399, 
    -1.138199, -1.893936, 0.6868057, 0.6972198, 2.056084, -1.287422, 
    -0.9046021, -1.389229, -5.968407, -3.243408, 4.807892, 3.020912, 
    3.101929, 6.415741, 2.658188, 2.094894, 1.689682, 3.511795, 3.092789, 
    2.991486, 1.836807, -1.066071, -1.92543, -2.30043, 0.5956421, 4.696953, 
    3.717804, 1.490715, 0.3266602,
  3.317291, 2.222214, -1.58194, -1.659012, 2.080048, 1.93187, -1.296249, 
    -6.118637, -5.364471, -2.057968, -0.8485718, -3.481155, -0.269165, 
    3.290741, 1.832657, -2.636612, -0.9181213, -2.149384, 2.141769, 1.889175, 
    -1.067337, 1.187088, 0.14151, -0.2436371, 7.385788, 5.736267, 8.601929, 
    10.22015, 6.743576, 11.44463, 13.11493, 9.452179, 7.663116, 8.614685, 
    9.092819, 4.723007, 5.227982, 6.422501, 3.899063, 2.377945, 2.664963, 
    3.476685, 0.6839752, -2.880081, 2.874603, 1.091232, 2.128212, 5.54361, 
    4.587875, 6.339951, 4.440994, 5.127457, 2.563919, 1.135529, 1.233185, 
    -0.2339935, 0.5490723, 3.983673, -1.461868, -4.634521, -3.32959, 
    -3.562653, -4.442871, 1.367538, 4.052719, 1.925354, 1.302948, -1.205872, 
    -0.3865967, 4.033142, 2.264145, -0.1670837, 0.1493073, 1.15477, 1.225372, 
    0.6087036, 4.615959, 3.271698, -0.2655487, 0.1277161, -0.5839996, 
    -1.401459, 1.007126, 2.069901, -0.503006, -1.722549, -3.255356, 
    -1.892334, -2.930359, -4.076202, -5.876465, -2.334534, 2.327164, 
    1.043076, 4.930832, 4.491745,
  4.983963, 1.2173, 3.134995, 6.317032, 4.072235, 1.55481, 0.01417542, 
    -6.405365, -6.942337, -3.335831, 1.483704, 5.826401, 1.602463, 3.942825, 
    1.069382, 0.5199127, 6.415466, 3.000626, 2.080582, 3.692307, 2.561813, 
    7.136566, 8.334488, 11.07928, 6.876678, 5.725632, 7.357666, 11.32381, 
    11.17953, 8.353241, 8.937607, 5.42276, 6.417023, 10.48318, 11.99648, 
    6.767303, 1.272247, 0.3274384, 4.129791, 2.925858, -0.3704529, 
    -0.6613464, -2.043625, -1.712906, -0.1413116, 2.180847, 5.687363, 
    9.031586, 0.5227509, 1.822769, 3.631363, -1.332443, 0.7011566, 2.983459, 
    4.200897, 0.4131317, 3.057922, 2.599594, -2.783218, -0.9767151, 4.124069, 
    4.2285, 1.494385, -0.01914978, -0.7329559, -2.550156, 0.1675568, -3.5952, 
    -2.089462, 1.07225, -2.443893, -0.4444122, 0.1618347, -0.4595184, 
    1.069122, 1.942032, 5.3246, 5.659981, 1.124832, -3.630096, -4.151947, 
    -4.453537, -6.112137, -5.052246, -5.215775, -5.717087, -7.290253, 
    -8.611084, -5.9702, -2.834518, -1.361084, 1.030319, 2.267563, 2.187607, 
    3.423294, 6.67981,
  4.59021, 7.462616, 9.70195, 4.489456, 1.050156, 3.782974, 2.582962, 
    1.029861, 1.831161, 6.661591, 10.12381, 9.197769, 6.788925, 7.598282, 
    3.342819, 2.601425, 10.21391, 9.937881, 8.688126, 11.77225, 14.83032, 
    10.09023, 9.616257, 7.654816, 3.132156, 1.350388, 3.491791, 3.862106, 
    2.622528, 1.05246, 5.900635, 12.83397, 10.39413, 1.948318, -2.037354, 
    -4.763138, -3.840485, -2.135818, -5.05069, -4.439987, -11.05975, -13.241, 
    -11.67433, -9.694382, -5.712112, -1.803787, 2.986832, 3.616776, 
    0.1495819, 0.5555725, 7.194107, 4.075882, 2.01236, 1.011826, 2.82225, 
    5.930588, 0.4209442, -4.238449, -5.829071, 1.670166, 2.489166, 
    -0.3931122, -0.682724, 1.163925, -0.465271, -1.923843, -1.979065, 
    -3.137634, -2.594177, -5.205872, -6.895203, -7.526718, -5.71994, 
    -0.2149963, 3.806107, 1.807159, 4.190781, 5.583191, -9.475128, -10.1301, 
    -6.236343, -4.304077, -6.079025, -2.1754, 0.901413, -5.256927, -7.338959, 
    -3.714218, -3.837402, 0.2506409, 2.724579, 4.641006, 6.258438, 6.493347, 
    7.661301, 5.744385,
  3.623611, 5.416306, 6.692871, 1.92778, 3.319443, 8.26944, 7.131149, 
    9.756424, 6.687637, 3.572296, 5.279327, 8.523605, 2.801727, -0.422226, 
    1.098312, 2.285812, 5.4702, 6.018906, 8.60405, 8.217606, 5.827499, 
    0.01577759, 1.444443, 2.192093, -1.365204, -2.764679, -5.871964, 
    -6.758942, -4.288132, 2.42334, 13.98245, 16.70457, -1.275101, -10.7803, 
    -11.42952, -17.16858, -12.56259, -7.145416, -13.14436, -17.30663, 
    -25.0798, -22.92796, -15.99648, -11.27901, -7.472244, -0.6902313, 
    -0.7290344, 2.930069, 3.427979, 5.477997, 1.282669, -0.2339935, 
    -2.531647, -3.462891, 1.302475, -0.6977997, 0.3576965, -0.5852966, 
    -4.372543, -0.8537903, -2.170715, -3.434006, -2.098846, 1.40976, 
    0.4894409, -2.492065, -4.6017, -7.097015, -4.980057, -3.655884, 
    -3.920181, -5.967041, -2.345703, -2.504028, -1.12587, -2.307129, 
    -1.140457, -2.964157, -9.226135, -6.807663, -7.451706, -0.8433838, 
    -5.579315, -8.9785, 0.4170837, -0.6626434, -4.509766, -4.539459, 
    0.2931061, 3.96315, -0.03633118, 0.973587, 2.257172, 7.255875, 4.873581, 
    1.913681,
  3.32515, 1.825424, 0.5123901, -0.9532318, 0.7563782, 3.475922, 1.830872, 
    5.096008, 7.094681, 4.044434, 0.1637115, 3.175415, 4.872803, 8.21579, 
    10.63713, 6.074646, 9.787659, 6.456421, 3.09314, 3.075684, 1.636093, 
    4.442871, 1.08168, -3.310532, -6.158432, -7.956375, -4.863892, -5.82196, 
    0.465271, 5.012665, 7.911087, -1.312378, -12.85298, -15.63501, -16.33528, 
    -19.42615, -12.01132, -11.53032, -16.66782, -16.76471, -23.74022, 
    -22.49854, -2.80011, -5.627701, -3.164932, 1.133759, 0.1040649, 7.462662, 
    -2.324051, -5.455307, -8.669388, -0.1751251, 0.1962585, 1.215744, 
    0.8816528, -5.828766, 1.258469, -2.729034, -7.354294, -4.973831, 
    -4.713928, -4.013931, -7.849854, -4.111053, -5.847244, -7.923019, 
    -6.32016, -8.972244, -4.763107, -5.136826, -8.131607, -6.036835, 
    -0.205307, -3.181351, -3.423523, -4.247238, -6.804535, -8.324066, 
    -10.5397, -3.419891, -0.503006, 5.891785, 0.3311005, 8.494125, 10.73454, 
    0.9636993, -2.079788, -0.9323883, -0.644104, -3.688644, -4.817291, 
    -4.726669, -0.1177979, 1.749115, -4.852448, -1.956604,
  -0.2271729, -0.3938446, 0.2433929, -1.497253, -4.168365, -3.955078, 
    -4.701935, 1.865784, 0.387146, 8.21814, 2.080627, 1.060547, 4.110306, 
    9.054321, 8.423859, 9.018661, 6.256927, 0.591568, 2.608749, 3.997025, 
    4.124634, 7.032196, -0.4206696, -1.225876, -2.359222, 0.7970276, 
    -0.6912384, -0.1404572, 2.051987, 4.172287, -3.13504, -7.490997, 
    -14.07019, -9.357666, -14.61002, -20.19856, -15.98502, -20.25819, 
    -20.9902, -23.16417, -26.31911, -11.36729, 1.619949, -1.861557, 
    -1.831604, -0.0526886, -0.1719666, -0.4292603, 1.094177, 1.522034, 
    -3.673538, -2.826401, -1.783691, -4.757416, -6.463654, -7.067825, 
    -5.906631, -12.04646, -11.71991, -12.41522, -11.20636, -10.64177, 
    -9.31572, -6.687592, -7.936035, -4.200104, -1.221451, -1.175354, 
    -0.0001068115, -5.191772, -3.794098, 0.8631897, -3.416779, -5.981857, 
    -0.420166, -3.702209, -5.784515, -8.323822, -13.28293, -1.499313, 
    10.07698, 13.74052, 6.629852, 18.10432, 13.02751, -1.028732, -3.499313, 
    -4.391495, -6.342819, -8.137863, -4.259216, -3.742798, -2.364426, 
    -3.94931, -3.634201, -6.540466,
  3.458496, 2.850403, -4.657913, -4.052704, -4.417023, -3.525391, 1.470428, 
    1.500397, 4.908966, 11.32565, 2.13501, -4.265747, 13.2012, 18.58975, 
    0.6431274, 1.606934, -0.1602631, 1.834534, -0.8162537, -0.5995789, 
    -0.8107758, 0.3668365, -3.397751, 3.346252, 4.03064, 0.6918335, 5.916824, 
    9.209549, 4.833481, -2.153259, -9.117798, -9.325104, -10.49335, 
    -19.82227, -25.93527, -22.42538, -20.45093, -18.1488, -19.13762, 
    -20.14203, -6.570419, 2.968643, 1.593918, -3.417023, -0.1769104, 
    4.623337, 2.767868, 5.385056, 3.332199, 1.777496, 1.416306, -3.148788, 
    -1.892807, -1.351395, -1.572235, -3.482132, -6.686813, -6.868591, 
    -5.840454, -6.095413, -8.791763, -10.63916, -9.167282, -3.867294, 
    -0.7243195, 2.366318, -2.428482, -0.9469757, -2.015717, -0.7922821, 
    1.525696, 0.1600647, 1.76944, 1.128265, -0.7597656, -13.27666, -7.139679, 
    -10.4061, -12.19492, 14.04703, 12.49834, 12.02596, 6.975403, 14.06058, 
    27.72047, 11.76215, -7.968582, -11.12563, -11.81026, -12.48163, 
    -10.89751, -5.480072, 1.728806, -1.28241, 2.478546, 2.901978,
  3.00563, 2.863922, 0.03451538, -5.012909, -2.217834, 1.85144, -2.181091, 
    -3.224823, -0.4829712, 7.918365, 2.017578, -7.485809, -2.637619, 
    1.692062, -2.309998, -2.4673, -2.136032, -2.769882, -0.5701447, 1.054337, 
    1.40303, -2.072754, -2.009735, 0.8066711, -2.179001, 3.15538, 3.546265, 
    7.776474, 2.213684, -2.579559, -7.237335, -6.30896, -7.790741, -11.38602, 
    -16.2056, -17.60663, -12.61392, -10.98813, -7.330078, -2.761566, 
    1.944183, 2.977249, 0.2806091, 7.029587, 5.555099, 8.430374, 7.928284, 
    10.65146, 8.342865, 8.149643, 6.101196, 6.586624, 5.342621, 7.349915, 
    4.200684, 0.1907959, 2.274124, -1.900101, 0.7915649, 0.8613586, 
    0.3931274, -0.4318695, -0.4506226, 3.971771, 2.317078, 6.663696, 
    0.8639679, 1.886612, -1.515457, 2.605377, 1.732193, 0.3603058, 2.617584, 
    -1.57489, 0.5366211, -4.938629, -8.238892, -8.752228, 1.364197, 18.20276, 
    4.614471, 4.786072, 2.412109, 8.068359, 23.35329, 7.178772, -14.28917, 
    -13.63603, -13.32433, -10.81755, -0.3292694, -0.4581757, 5.7314, 
    7.013702, 6.089996, 1.533234,
  5.681381, 6.913925, -10.95975, -6.511078, 2.234497, 4.351166, -3.271484, 
    -2.726166, 2.908997, 4.65976, 12.3811, -8.500671, -8.046478, -3.01004, 
    1.807968, 0.9436035, -1.000153, -0.3904877, -1.274857, 0.1816711, 
    0.4446869, 3.207718, 5.322037, 3.279327, 5.115524, 5.640793, 4.173599, 
    2.968658, -1.098846, -6.356384, -5.275085, -6.995667, -7.319153, 
    -7.219391, -9.496735, -11.52802, -7.723572, -8.126709, -7.459503, 
    5.072296, 0.2553406, 4.660583, 0.1881866, 5.893356, 3.68425, 6.194946, 
    9.069946, 7.332962, 8.496506, 9.57695, 7.236084, 6.543091, 6.943634, 
    5.748291, 4.557159, 4.030853, 1.981628, 4.608978, 4.242554, 1.657684, 
    4.360565, 1.095474, 3.352509, 1.477509, 0.04417419, 2.368393, 3.451462, 
    4.402496, 4.572052, 7.593399, 4.979065, 3.814224, 5.034241, 0.4529724, 
    0.04391479, -4.696991, -8.752182, -0.9738464, 21.20511, 6.101166, 
    -0.4959717, 0.7139587, -0.7808838, 0.888916, 8.890228, 3.203537, 
    -10.04515, -12.55428, -6.976669, -2.954788, 4.364746, 8.402496, 7.564758, 
    11.05641, 6.884796, 7.774597,
  3.24469, 5.954559, 2.491821, -10.30923, -0.2425537, -1.60379, -7.040222, 
    -8.266785, -2.562897, 11.43008, 9.647003, -1.235535, -1.698578, 8.097778, 
    0.7055969, 5.799866, 1.600922, 2.346741, -5.289169, -2.457428, 
    -0.5852966, 3.193604, -0.6967163, 6.058502, -4.086823, -0.5808411, 
    1.924896, -2.18631, 4.176666, -2.250397, -4.152222, -5.498291, -5.251648, 
    -7.230042, -9.359222, -9.093842, -10.4118, -17.96573, -21.547, -4.873016, 
    0.2532959, -8.635513, -3.553772, 1.107712, 6.625168, 9.046249, 8.118652, 
    7.272293, 1.201202, 4.117599, 6.398605, 6.666824, 5.222549, 2.547806, 
    0.3155212, 3.154297, 3.877228, 3.790771, 6.314209, 7.662628, 5.452728, 
    1.861588, -0.02093506, 0.637146, 5.944946, 4.285065, 7.597031, 7.225433, 
    8.256943, 10.64287, 7.401733, 5.513443, 2.295959, 6.425659, -4.176941, 
    -4.499603, 11.1707, 10.44232, 0.7623901, 4.466278, -0.4962158, -1.079041, 
    -2.114471, -0.8008728, -0.3279419, 5.611053, -0.117569, -9.427185, 
    6.275162, 6.297043, 6.952499, 10.68687, 10.45381, 11.71344, 3.791824, 
    6.321228,
  5.713181, 3.651154, 4.294693, 4.051941, 2.038147, 1.709778, 1.937927, 
    -6.47847, -7.039703, 2.35611, 20.19313, 8.398315, -0.1967468, 2.441772, 
    3.565002, 6.494415, 1.523834, 5.31131, 5.32254, 7.442581, 8.620712, 
    7.476715, 6.915253, 5.85849, 0.7212219, -2.761841, -5.634003, -5.783691, 
    -0.5480194, 4.349884, -1.157959, 1.647278, -0.05221558, -0.5040283, 
    0.8769531, -4.933472, -11.57536, -26.40485, -19.53712, -14.08345, 
    -11.12979, -6.628754, -1.771454, 8.716049, 15.03792, 22.42906, 17.04782, 
    19.87646, 12.5999, 7.298859, 5.109543, 1.295471, 0.04910278, -2.120148, 
    1.220978, 1.13501, 2.627502, 3.538666, 4.678284, 7.401947, 4.066528, 
    5.479828, 8.638916, 6.333481, 6.485565, 10.28714, 8.751999, 10.84001, 
    12.17177, 9.689224, 9.349106, 11.20433, 7.331635, 8.659515, -5.960007, 
    -1.281097, 4.095459, 11.89334, 11.83844, -7.331345, -7.397522, 2.903259, 
    0.488678, -0.4712219, 3.441071, -0.7797852, 6.00769, -0.732132, 7.10144, 
    4.810059, 4.619949, 7.869431, 10.18871, 5.160034, 7.87204, 9.687637,
  1.744415, 9.05484, -2.468628, -7.10379, -0.5415039, 8.556152, 5.459778, 
    -0.7457275, -10.88345, -10.13994, 2.506683, 8.95929, 4.822784, 3.411316, 
    2.216003, 3.220428, 3.337891, 3.475922, 8.96756, 9.34259, 9.261841, 
    6.086304, 2.607697, 0.1699219, 5.649597, 0.9769287, 1.118866, 12.86891, 
    -1.948792, -5.015747, -12.85065, -20.21468, -6.830048, -7.97641, 
    -7.70871, -1.507126, 0.8308411, 9.321716, -9.143066, -16.41106, 
    -9.520157, 3.403809, 0.1801147, -0.3998413, -6.530045, -12.17903, 
    -13.43057, -17.01938, -17.27017, -16.36523, -10.66443, -1.842316, 
    1.785797, 5.680359, 6.833191, 6.767548, 6.537872, 4.589935, 5.354553, 
    7.894409, 4.258972, 2.748291, 6.164459, 8.086853, 6.492035, 10.5405, 
    7.63501, 11.56967, 7.812103, 7.01474, 0.09622192, 0.696228, -1.424622, 
    -6.209503, -5.174057, 6.830612, 4.41655, 12.37282, -0.4730072, -23.46262, 
    -14.25923, -1.713928, 9.161865, 7.326172, 0.9022217, 0.2189331, 
    -2.443604, -1.959778, -5.724335, -3.942841, -3.587097, -3.410553, 
    0.8584595, 1.583984, 2.036316, 3.280334,
  -5.599625, -1.172485, -2.850357, -0.3113556, 7.683762, 11.29051, 13.50017, 
    11.02852, 6.424072, -0.569931, 1.275421, 4.322784, 6.816803, -2.166534, 
    -3.637634, -1.893372, 0.9805908, 3.119904, 11.59961, 7.299866, 4.772552, 
    -0.1644287, 0.4245911, 1.719666, 1.891785, 2.255859, 5.580841, 22.40871, 
    0.4512177, -12.22852, -18.33293, -11.39729, -2.0327, -14.06963, 
    -13.21886, -3.962845, -8.416504, -5.192551, -5.319122, -3.953751, 
    -0.4256439, 4.287918, -5.515472, -14.77144, -20.85741, -26.79987, 
    -31.65898, -33.67822, -29.77667, -22.8345, -18.6785, -11.84464, 
    -8.781097, -4.711792, -2.322998, -0.5462036, 0.7618713, 3.358765, 
    2.720459, 1.837677, 1.531952, 2.279022, 0.8243103, 5.439972, 2.658997, 
    1.891541, 0.9165344, 4.147522, -0.07904053, 0.03973389, -10.90532, 
    -16.93581, -22.36598, -24.59854, -14.72073, 4.732384, 7.528809, 
    -0.2628632, 0.2761993, -12.07121, -4.648285, -4.084747, 14.84152, 
    -0.5386963, -0.368103, 0.4902649, 0.07043457, -5.579788, -8.291016, 
    -5.421509, -7.398834, -5.968628, -5.583191, -5.199615, -1.374359, 
    -7.807144,
  -3.393112, -5.15271, -3.143906, 10.04202, 11.96838, 7.162399, 12.1447, 
    16.92464, 20.88501, 15.90198, -0.7267532, 13.7137, 5.032959, -3.753265, 
    -5.347015, -6.193878, -4.493103, -6.130341, -1.854019, -4.210526, 
    -3.969894, -8.21962, -7.419388, -2.255844, 0.02069092, 1.895966, 6.07724, 
    -3.028275, -7.485519, -8.077454, -5.73082, -0.6946411, -10.1501, 
    -11.63786, -10.62457, -11.78473, -8.597488, -2.063385, 2.810333, 8.07724, 
    11.39365, 15.03973, 9.567078, -3.113892, 0.3699493, 7.797821, 1.881668, 
    -0.4167633, 0.9014587, 0.9478149, -0.2211914, -4.678223, -10.46806, 
    -6.288116, -4.698029, -6.550354, -5.804794, -2.014938, -1.962097, 
    -0.1938782, 0.7608337, -3.752991, -9.065216, -7.980057, -7.250366, 
    -5.100357, -9.956604, -0.9021759, 2.385834, 0.5342865, -7.629532, 
    -19.8027, -34.98135, -27.66161, -11.05069, -6.634277, 0.4756317, 
    -8.011292, 22.68005, 10.03116, -0.4550781, -1.801453, 4.295441, 
    -5.362625, 4.121002, -3.257904, 4.341568, 10.6059, 6.413712, -0.7625885, 
    -2.763641, -6.217285, -3.640213, -2.054825, -2.145721, -7.434784,
  7.422531, 13.27641, 17.44881, 22.00459, 11.47205, 7.437408, 6.073074, 
    9.277252, 19.76709, 28.93344, 36.88162, 1.712891, 1.150391, -5.344147, 
    -6.337097, -8.580872, -10.5405, -11.23265, -12.41286, -16.4462, 
    -8.833954, -6.832947, -9.94046, -7.948273, -6.381363, -1.084213, 
    -1.019882, -2.867813, -22.84491, -20.94231, -9.057144, -5.935776, 
    -8.874573, -0.9355621, -8.513641, -9.162857, -6.102432, -0.7472382, 
    3.367081, 3.940536, 11.5986, 12.46996, 6.486893, 3.46553, 8.573608, 
    13.05147, 7.481415, 2.315277, 2.201981, 13.09288, 16.20901, 12.2939, 
    8.757202, 7.645477, 11.06787, 7.861099, -0.9995728, -0.7688446, 1.973343, 
    8.747559, 18.82411, 4.178284, 1.77803, -4.198547, 0.1230927, 1.829071, 
    0.0254364, 8.908234, 16.09599, 16.66577, 16.71526, 9.64624, 3.058472, 
    9.915482, 12.90608, 24.24332, 12.3275, 24.45172, 16.46005, 10.71082, 
    -3.439697, -3.342041, -2.840759, -0.2032776, 1.039749, -2.643097, 
    0.07720947, 3.437378, 7.248032, -1.142044, 2.095734, -5.35791, 3.05719, 
    19.96053, 16.33865, 15.00558,
  -1.898788, 0.6319427, 1.149384, 3.375641, 3.66394, 6.727997, 6.841034, 
    14.06863, 7.751434, 21.07671, 6.077484, -3.765472, 0.7004089, -4.984467, 
    -4.890503, -0.103241, -8.016266, -7.067581, -8.105835, -6.673782, 
    3.902939, -4.270203, -6.890717, -0.1714935, -1.835541, -6.405579, 
    -8.134506, 1.955826, -12.89939, -16.29234, -11.73422, -8.512344, 
    -7.982376, -3.557922, -16.06833, -11.05403, -8.711288, -6.981598, 
    -1.993851, 0.7243805, -0.3264008, 2.970474, 4.744965, 3.348602, 4.665253, 
    3.491318, -6.321716, -9.009735, -3.074844, 4.433746, 7.032181, 4.481644, 
    -2.356613, -0.7243347, 0.8563843, 0.6058655, -1.563934, 0.9696808, 
    -3.334213, 4.018341, -0.219101, -3.664185, -8.912354, -9.501938, 
    -9.744644, -3.801147, -0.05531311, 12.67099, 9.049637, 11.33923, 15.8405, 
    23.50432, 37.16913, 31.13162, 14.41866, 16.56369, 3.787903, -2.778778, 
    0.973053, -0.3694153, 5.969406, -0.3701782, 0.2876282, 0.9733429, 
    -6.410553, -2.082947, 1.864212, -0.6662598, 1.942871, 0.7824402, 
    2.563446, -4.189957, 3.168396, 13.85121, 4.009018, -0.4402161,
  -0.8438721, -2.242035, 0.7366028, -0.7996216, -1.404297, -1.990997, 
    -2.181641, -0.553772, -1.232941, -0.3824158, -2.208984, -5.018616, 
    -5.956635, -8.196472, -7.875336, -7.205292, -1.317322, -3.30249, 
    -3.247757, -5.006363, -5.051483, -7.064743, -2.751923, 5.153549, 
    -6.649582, -16.65923, -12.13475, -21.3665, -22.47198, -20.33813, 
    -16.37068, -8.130325, -1.318619, -2.265228, -7.902725, -6.570435, 
    -6.991501, -10.53447, -4.187607, -5.998795, -1.781616, 9.109802, 
    10.97958, 3.387924, 1.390259, 3.184799, 2.840271, 4.950424, 6.424911, 
    4.659271, -3.158447, -3.871994, -6.237076, -2.388657, 7.41864, 
    -0.1800537, -2.211548, 0.8785553, -0.2045135, 1.71788, 2.387146, 
    0.1631622, 0.5715027, -0.7800446, -4.613892, 1.280334, 2.515274, 
    -1.765717, 1.970718, 14.9913, 13.95612, 32.13969, 39.62172, 9.330627, 
    6.406937, 5.973846, -0.7175903, -1.272247, 3.225677, 0.04959106, 
    -0.9998474, -0.8972321, -2.183426, -6.467819, -3.514679, -2.429779, 
    -1.914154, 6.80014, 5.421524, 6.394928, 1.493103, 3.903015, 3.349335, 
    1.303253, -1.922791, -1.815735,
  -1.037903, -2.310822, -1.486603, -3.05246, -2.568878, -4.097504, -3.676483, 
    -4.108459, -3.755066, -3.095184, -3.581635, -6.455078, -6.256134, 
    -7.84494, -9.769165, -12.94281, -13.60117, 1.72644, -2.589966, -8.450119, 
    -6.780075, 7.197769, 2.987335, 6.726685, -6.475876, -9.460815, -6.076721, 
    -1.457428, -9.401688, -10.44437, -8.627441, -6.212341, -10.30818, 
    -4.599335, -8.157669, -4.735504, 0.2079773, 1.809799, 2.501465, 5.776993, 
    7.522034, 11.98401, 10.00771, 3.257462, 1.043381, 1.444687, 7.51239, 
    7.882721, 12.80669, 9.424652, 2.688187, 3.454834, 3.875168, -1.29776, 
    -0.6516724, -4.206604, 1.38974, -0.1045227, 2.206665, 2.181152, 4.717087, 
    9.266571, 12.14128, 9.768631, 9.439453, 9.241821, 3.53688, -3.901154, 
    8.445724, -14.046, -1.837601, 28.20042, 28.22803, 3.392334, 5.685059, 
    7.517349, 6.659012, 5.714218, 3.524643, 1.345215, 0.2707367, -3.017548, 
    -3.219376, -5.286285, -0.5076447, -1.393845, 0.141571, 4.938431, 
    0.8569031, 6.652191, 0.03448486, 1.365509, 2.801208, 1.310059, -1.998016, 
    -1.759216,
  1.970764, 0.8894653, 1.618103, -2.088409, -2.404572, -3.129303, -3.320709, 
    -4.181396, -5.052734, -4.606903, -5.059235, -6.946747, -6.178802, 
    -5.772522, -9.414734, -11.85687, -14.13843, -11.71732, -16.32327, 
    -14.6837, -14.51808, -9.345413, -7.915985, -6.315994, -6.446503, 
    -4.043854, 5.352768, 9.503738, 3.845169, -0.06703186, -10.35739, 
    -5.802444, -11.70712, -11.14098, -1.575104, 1.615524, 7.531418, 8.485062, 
    3.410843, 7.129852, 7.660583, 5.486618, 6.646255, 2.56813, 8.695999, 
    7.143646, 9.841309, 10.36371, 10.17386, 16.32826, 8.597824, 5.601212, 
    1.319687, 3.097824, 2.28949, 2.997299, -1.720932, -2.77536, -0.8144226, 
    -1.044617, 5.292099, 4.134277, 2.781158, -1.954834, -1.136322, 4.052216, 
    8.632172, 5.04129, 12.55275, -5.939453, -5.126923, 0.8087158, 4.885315, 
    1.12178, -1.207123, 2.476212, 5.576736, 6.470734, 3.734543, 5.941055, 
    1.595993, -1.444885, -3.726151, -1.592285, -8.517029, -2.830566, 
    3.891312, 3.381668, 6.847031, 10.26837, 7.638153, 1.535034, 0.3415527, 
    2.402527, 0.5535278, -0.137085,
  1.935577, 2.64621, 5.154816, 1.837402, 1.685272, -2.070679, -3.096191, 
    -3.352448, -3.387085, -3.981659, -5.357178, -5.723572, -5.952728, 
    -4.754028, -5.369659, -7.508423, -7.608704, -9.456085, -15.13086, 
    -9.991501, -11.24596, -10.10063, -0.2769318, -2.496246, -4.245209, 
    -0.03013611, 1.152191, 9.644882, 8.490982, 2.080093, -12.60452, 
    -13.36574, -4.082413, -4.207397, -4.225098, -2.287079, -0.8396912, 
    5.329849, 4.864212, 10.99469, 8.039215, 4.991043, 7.310318, 9.029846, 
    9.979843, 6.655899, 5.890533, 7.190002, 5.096008, 5.335846, 6.475677, 
    3.747818, 1.539734, -2.329529, -0.5988007, 0.7577209, 2.261887, 
    -2.207901, -0.6977539, 3.019684, 0.2509308, -4.717285, -6.986832, 
    -11.12827, -13.63631, -0.9376221, -0.1092224, 2.311081, 6.812119, 
    -1.194122, -4.38942, -8.777176, -6.296188, -4.100357, -0.1446533, 
    -2.309738, 0.04000854, -1.208176, -1.432129, -0.7701416, -0.4644165, 
    5.983231, 5.567612, -0.9334412, -4.419373, -3.220413, -5.170929, 
    2.079849, 5.726715, 4.417618, 9.16214, -1.086304, 0.09725952, -1.037354, 
    -0.2027283, 2.015472,
  5.367584, 7.359253, 3.96759, 1.254303, 5.111328, 0.6576843, 0.2933655, 
    -1.22644, -3.017059, -2.818878, -3.625366, -3.891785, -4.33606, 
    -3.912354, -4.309204, -5.205597, -5.36026, -5.967804, -3.098572, 
    -4.382172, -7.982422, -16.6936, -16.98741, -16.85976, -16.27617, 
    -17.01839, -4.48819, 5.339684, 11.49332, 8.425629, -6.113373, -10.92822, 
    -9.106873, -8.473801, -2.783173, 1.823074, 2.422302, 5.592606, 7.353806, 
    9.367355, 8.487396, 4.252762, 5.646255, 0.3290558, 4.735306, 6.108246, 
    5.009796, 1.84288, 2.938965, 3.398071, 3.222824, 1.705109, -0.611557, 
    2.851456, 0.8340149, -0.9131165, 0.003555298, 1.056946, -0.3907166, 
    -1.35817, -2.432648, -4.07431, -9.41391, -17.00114, -5.332428, -3.395721, 
    -6.548035, -1.239426, -2.304016, -6.415482, -5.56781, -3.289688, 
    -2.576401, -3.400879, -1.693085, 3.060837, 0.5251617, 1.862411, 
    0.2147522, 2.283508, 2.273849, 1.58194, 3.89444, 5.33194, 3.418915, 
    0.467865, -0.8987885, -0.5631256, -1.385254, -0.1797791, 9.906158, 
    9.893646, -4.608948, 0.3808594, 1.78476, 1.594421,
  8.493896, 12.63507, 15.50304, 9.002762, 1.029327, 0.1900024, 4.892853, 
    0.4129028, 0.5397034, 2.019135, -1.508728, -2.627472, -3.973816, 
    -2.122528, 0.9540405, -0.7891846, -3.196991, -2.05246, -1.150909, 
    -0.511322, -0.7472534, 3.381668, 3.74678, -3.934998, -5.975357, 
    -5.819107, 0.1430969, 1.559219, 5.278503, 4.396988, 1.000122, -4.850632, 
    -10.05713, -8.173004, -7.840988, -4.552963, -4.211868, -2.644165, 
    -0.2175903, 2.853256, 5.001968, 0.8165741, 1.930099, 0.03688049, 
    0.7949524, 6.338974, 7.465271, 1.549377, -2.976395, 1.912399, 4.068924, 
    3.742874, 2.856415, 3.645737, 3.022034, 3.027771, 2.006943, 1.613434, 
    0.7754211, -0.0758667, -0.3920288, -2.448013, -9.565491, -8.214447, 
    -7.545959, -6.778259, -3.243622, -0.3438568, 0.07984924, -1.617279, 
    -5.191757, -3.853745, -2.832397, -3.653732, -3.963135, -0.3644257, 
    3.574112, 4.716309, 1.449112, 0.2254181, 2.783234, -0.9464417, 3.04834, 
    6.227768, 0.4827271, 1.612396, -0.5139008, -2.334991, -3.700104, 
    -4.005829, -2.796448, 6.381683, 5.341309, 0.436615, 7.123566, 6.184784,
  12.87933, 4.174393, 2.425949, 3.178818, 4.835052, 4.898865, 10.39653, 
    7.279846, 7.201965, 9.462112, 4.558197, 3.029053, -0.2579193, -5.256363, 
    2.23114, 3.161575, 2.519928, -0.7972717, -2.012909, 3.439209, 4.432724, 
    2.515259, 1.692078, -2.183456, 0.3400116, -3.435776, -5.898788, 
    -0.06416321, -1.583435, -5.801422, -2.544418, 2.182953, -3.71991, 
    -3.808701, -6.538147, -7.798279, -2.140213, -3.544937, -3.996506, 
    0.8014069, 0.8865814, -0.8519897, -3.882446, -2.35405, -8.837906, 
    -11.341, -4.698059, -2.138687, -5.600937, -1.971512, 1.321732, 2.487869, 
    4.869904, -0.09988403, 1.710007, -0.3748627, 1.23764, 4.863937, 5.499863, 
    1.966553, -1.044907, -2.481079, -7.120163, -7.294388, -5.651138, 
    -2.618835, 1.067093, 1.566833, 4.468384, -6.315979, -1.80426, -0.2581787, 
    -2.596985, -1.695419, 0.7832031, 3.927734, 5.959793, 3.297546, -1.643326, 
    -1.874069, -0.07824707, 5.443115, 3.022797, 0.08686829, 3.455612, 
    3.769684, 2.246521, -0.5230408, -3.080582, -2.979263, -2.419373, 
    4.012131, 3.5439, 5.049118, 8.700424, 12.43402,
  20.21886, -4.001938, 3.567352, 10.42435, 2.640015, 10.26208, 13.94334, 
    7.224915, 5.254852, 4.418121, 7.634277, 14.36394, 13.37878, 7.136353, 
    2.026993, 2.888977, 3.550674, 2.713699, 2.609543, 2.835587, 4.587921, 
    9.063705, 4.437408, -0.6667633, -3.25296, -3.248276, -3.732651, 
    -4.748016, -2.153488, -2.832642, 1.362366, 1.482941, 4.400635, 2.758438, 
    4.484756, 4.316513, 4.658234, 7.468094, 4.661804, 1.549072, 3.049042, 
    -0.5772247, -2.207962, 1.135269, -1.185028, -4.729309, -2.513168, 
    -3.48114, -3.975677, -5.051437, -3.261856, 1.136826, 2.2845, 2.53241, 
    3.289673, 1.5905, -1.553284, 0.07537842, -0.5991211, -0.8644562, 
    2.574081, -2.154816, -4.680817, -2.614944, -3.107391, 3.469437, 4.736618, 
    4.259277, 0.3613586, -7.614182, -8.685532, -4.67511, -2.390488, -5.57901, 
    -3.603241, 2.190216, 3.455307, 1.898575, 0.7014618, 1.119934, 2.319138, 
    4.252716, 2.392822, 1.530853, 0.5693817, -2.161346, -1.234512, -1.246231, 
    -2.519684, 0.8553314, -2.042862, -1.595963, -0.08241272, 7.679321, 
    14.98396, 20.80638,
  9.350601, 2.328766, 11.65245, 10.94045, 5.295685, 5.653503, 11.82042, 
    8.969376, 4.410278, 4.064178, 0.03033447, 3.274857, 7.492813, 6.443619, 
    2.271759, 2.172531, 1.167603, 0.4501648, 4.637146, 2.000412, 2.865265, 
    5.888702, 8.807175, 4.804337, 2.600693, 5.030899, 8.863144, 5.067078, 
    5.000153, 1.326706, -0.711319, 3.725662, 7.849335, 7.508713, 9.30217, 
    3.601669, 3.286835, 3.229279, 2.685013, 6.541504, 4.456619, 5.156097, 
    5.785522, 1.048553, 0.3948975, 2.327454, 2.443329, -1.0327, -0.3959656, 
    -2.123062, -3.894928, -2.693375, -5.825668, -6.825165, -1.460815, 
    1.358414, -0.001449585, 2.412354, 0.227951, 1.586578, 2.489944, 
    -0.7561493, -1.91394, -2.560318, -4.577225, -8.003799, -3.002487, 
    2.36261, -0.2105713, 1.742844, 1.104294, 1.413132, 0.9787598, 0.167038, 
    -1.167847, -1.78479, 2.539429, -0.5449371, -3.049881, 5.278748, 
    0.06832886, -3.113953, -6.78244, -7.242615, -4.593903, -4.748062, 
    -3.382965, -6.2155, -7.868637, -5.557709, -3.600937, -2.828537, 1.818848, 
    0.5623627, 3.993347, 13.5647,
  10.37482, 7.514153, 3.161537, 0.9823761, -2.012939, 0.5529556, 3.157639, 
    6.775085, 5.419113, 3.453995, 3.3871, 3.597, 4.687347, 5.026398, 
    2.716766, 1.960022, 0.736557, 1.111038, 1.26442, 0.07562256, -0.5490875, 
    -1.735291, 1.883209, 3.744644, 7.16832, 12.13368, 7.916245, -2.805359, 
    -2.933212, -0.155365, -1.118896, 0.134491, 7.883926, 6.420944, 3.553482, 
    0.3842163, 3.986557, 4.290466, -0.1347809, -4.870453, -2.450424, 
    -1.047287, -3.107712, -2.573608, -3.163177, -4.340546, -3.63768, 
    0.331604, 1.556595, 1.138626, 1.947205, 2.807373, 2.013626, -1.112946, 
    0.6953888, 4.118042, 5.258163, 2.398262, 0.00112915, -1.715271, 
    0.3396606, -0.6616364, 0.1203995, -0.6108475, -0.4189301, -2.630386, 
    -2.280365, 1.060532, 3.362854, 6.093842, 3.686584, -0.05670166, 5.413651, 
    5.180832, 2.118835, 2.644882, -0.1751709, -5.231682, -1.923607, 2.840454, 
    -1.195724, -2.292358, -3.203308, -5.907722, -9.221283, -4.276459, 
    -1.498093, -9.277771, -9.606941, -5.779083, -9.494949, -10.48271, 
    -0.840271, -1.294159, -2.334274, 3.247772,
  4.300095, 0.7300262, -0.7025146, -4.031433, -0.4751816, 1.054001, 3.120132, 
    6.890976, 7.83889, 0.9292526, -0.06007385, 1.030807, 2.113632, 1.103989, 
    1.087051, -0.3061676, 0.1326447, 0.3672638, 1.414658, 4.167801, 3.509216, 
    2.348282, 6.280289, 6.736809, 4.062576, 2.161789, -0.06788635, 
    -0.3762207, -1.28611, -2.743141, -1.645737, -0.6142349, -1.756943, 
    -3.484558, -5.105385, -6.507996, -2.507729, -4.295212, -3.846512, 
    -6.128296, -6.630127, -6.109818, -4.43116, -3.521271, -6.61866, 
    -2.427765, 0.1154633, -2.47908, 0.6555557, 1.739937, 1.554253, 
    -0.6009521, 0.348793, -1.505119, 0.8477402, 1.503998, 0.6487885, 
    -2.28038, -0.9850693, -1.488968, -5.993141, -5.483253, -4.250954, 
    -6.263718, -1.651474, 3.495659, 3.338882, 4.477692, 3.371185, 0.8394165, 
    2.39592, 0.04122925, 0.7253494, -2.954597, -9.523613, -7.96711, 
    -5.976204, -8.06266, -3.520226, 0.9826431, -0.113205, -2.697571, 
    -1.428566, -2.671524, -6.26268, -4.092888, -1.055641, -7.538452, 
    -5.23793, -2.205383, -4.692886, -7.991318, -6.173607, -7.448868, 
    -5.709801, -3.159546,
  -1.776741, -1.640282, -2.147827, 1.588623, 5.113884, 3.031601, 1.345924, 
    1.078735, -0.8184052, -4.67205, -6.986618, -12.06214, -12.51501, 
    -10.94834, -8.518402, -5.508492, -1.742363, -2.037407, -0.452774, 
    -3.236374, -1.389496, 1.769623, 3.339409, 1.475609, -2.39315, -2.917358, 
    -2.162941, -5.713982, -7.794716, -7.916321, -7.069443, -6.619705, 
    -4.994171, -7.780373, -7.624138, -6.359543, -5.878571, -8.06398, 
    -8.953041, -9.204079, -9.532471, -10.14028, -7.128288, -7.428802, 
    -7.673103, -7.351486, -1.581421, 1.709457, -1.376213, -3.28299, 1.248009, 
    3.138634, -1.012672, -1.009285, 0.2474747, 0.8573837, 0.4347229, 
    0.6219635, 2.307381, 0.3789902, -2.180382, -4.203556, -4.412411, 
    -0.07829285, 1.626389, 2.050087, 3.599571, 3.706085, 2.494102, 0.7951431, 
    -4.151474, -3.794189, -6.79966, -7.956421, -7.369965, -9.068138, 
    -11.29392, -11.95044, -4.524658, -4.153557, -6.023613, -5.742882, 
    -2.474129, -3.616325, -6.556953, -7.962677, -5.710854, -5.476471, 
    -6.81736, -8.759033, -6.985596, -4.277512, -4.122047, -7.928032, 
    -5.815536, -1.693398,
  -3.295219, -2.803284, -0.9590302, 1.552959, 3.167797, -0.4608459, 
    0.6956558, 0.1784668, -0.5389786, -3.71085, -5.084538, -9.14027, 
    -10.25746, -11.30694, -8.103821, -7.380898, -6.56163, -6.917892, 
    -5.813461, -3.039246, -0.3796082, 1.170654, 1.357117, -0.6866379, 
    -4.696014, -5.34523, -1.673355, -3.251221, -4.90773, -5.228302, 
    -4.255386, -4.197037, -2.697823, -5.654335, -8.738205, -8.912422, 
    -8.274139, -4.399658, -2.75174, -5.068405, -5.859818, -5.71685, 
    -5.401222, -4.562424, -4.695488, -2.497581, 1.438103, 4.530815, 5.248528, 
    4.237579, 2.195656, 0.170929, -1.925697, -4.470226, -4.064762, -3.351738, 
    -1.779076, -1.762405, -2.304852, -4.048344, -5.313446, -7.026215, 
    -5.859818, -4.396011, -6.285583, -6.612152, -2.363205, 0.6784744, 
    0.4709091, -3.967888, -8.067627, -7.352249, -4.874916, -2.991577, 
    -2.590279, -5.545998, -6.179855, -4.595497, -0.932724, -1.203812, 
    -4.58741, -4.395477, -5.743652, -5.444176, -7.665802, -5.77803, 
    -4.357979, -0.9525146, -1.757729, -5.886887, -7.411888, -5.397575, 
    -2.536888, -3.82283, -5.966331, -5.837677,
  -4.511368, -4.795753, -2.907471, -1.681683, 1.068062, 1.950874, 1.725861, 
    1.489414, -1.512409, -3.664497, -5.568661, -7.540016, -9.175949, -7.8447, 
    -8.521519, -10.15903, -10.37074, -9.249386, -7.542103, -6.772835, 
    -7.259289, -8.155647, -7.59679, -5.659286, -5.498875, -5.153561, 
    -6.568928, -8.788719, -9.264233, -9.865276, -8.147316, -7.032722, 
    -5.634552, -5.225437, -5.102001, -4.529335, -6.901474, -7.026997, 
    -6.202259, -5.960594, -6.026733, -4.169708, -3.475697, -7.335323, 
    -10.09809, -10.36997, -7.823875, -4.860332, -3.924393, -4.938969, 
    -5.05069, -3.369705, -4.353565, -3.740795, -4.067612, -1.499645, 
    1.233166, 2.562851, 1.160767, -0.9556389, 0.3579025, -0.2910652, 
    -0.6871567, -1.283249, -0.6309052, 1.15556, 2.516228, 2.86858, 0.1724854, 
    -3.796013, -5.462677, -5.040798, -5.353558, -6.094448, -7.297836, 
    -6.837936, -3.605125, -3.425182, -4.725697, -4.898617, -3.754341, 
    -3.391052, -0.2426224, 3.601654, 3.254776, 3.743843, 3.008942, 1.444092, 
    0.01987457, -2.021011, -4.434811, -3.904068, -3.355118, -2.634552, 
    -3.350441, -4.687149,
  -1.224129, 0.2209206, -0.2548599, 0.6011314, 0.720665, -0.4535522, 
    -0.6571922, -1.159275, -1.580105, -2.646519, -1.623341, -2.379337, 
    -2.647831, -2.550442, -4.035061, -7.175686, -6.168919, -6.227509, 
    -6.249386, -7.604855, -8.885841, -7.592876, -5.819439, -3.972301, 
    -4.070221, -6.771515, -9.423603, -9.808498, -6.185322, -4.330898, 
    -5.478298, -7.82621, -8.918396, -7.98558, -5.21241, -2.849133, 
    -0.05928421, -0.5884514, -1.657982, -3.221264, -3.234547, -5.567619, 
    -6.568134, -8.455631, -9.045219, -8.036892, -6.50798, -4.977772, 
    -4.701469, -6.262672, -4.483768, -4.499138, -4.261375, -3.082714, 
    -2.986885, -0.8465157, 0.04880142, 0.2993164, -0.6577187, -0.4246445, 
    0.535511, -0.1324577, 0.5654526, -0.9790802, -4.02179, -5.736107, 
    -6.209801, -5.857719, -5.455372, -5.48064, -3.610584, -3.906418, 
    -3.919174, -3.4231, -7.827774, -10.18716, -8.324909, -7.469959, 
    -8.144699, -6.657722, -3.287933, -2.216309, -2.805389, -1.224899, 
    -0.7259598, 0.5112839, 1.642006, 1.960495, 0.5826263, -2.426735, 
    -4.445229, -5.480896, -7.435844, -6.426472, -4.062153, -3.129341,
  -0.7509422, -0.9842758, -0.9933929, -1.084274, -0.9894829, -0.6233406, 
    -1.238445, -1.406681, -1.886364, -2.232716, -2.073082, -3.041054, 
    -3.789742, -3.953548, -3.753288, -2.752764, -3.720474, -3.472557, 
    -5.113449, -4.96891, -4.391567, -4.525421, -4.834015, -4.464226, 
    -3.623856, -3.285835, -3.72073, -4.184532, -3.766823, -1.844948, 
    -1.39547, -2.793388, -4.973602, -6.567871, -6.39782, -6.610325, 
    -4.185326, -2.169697, -0.6111031, -0.640522, -3.366055, -4.170223, 
    -5.868137, -7.005634, -9.069958, -10.62621, -11.31241, -11.43558, 
    -10.87621, -9.37178, -8.35017, -7.005116, -7.047562, -8.258503, 
    -8.650684, -7.44001, -7.558495, -8.391312, -8.247307, -8.67569, 
    -9.548088, -9.291313, -8.316315, -6.080635, -7.200684, -7.835064, 
    -7.622303, -5.926468, -4.110062, -1.582199, -1.594955, -2.741829, 
    -2.859543, -5.764748, -7.364223, -6.596779, -4.179852, -5.56892, 
    -3.075951, -2.523613, -2.628304, -2.598091, -2.452263, -1.980644, 
    -2.009811, -2.480133, -2.474922, -2.017105, -0.9210129, -0.8288269, 
    -3.375175, -2.110332, -0.4407921, 0.3589554, 0.9782295, 0.4456711,
  -1.494431, -1.384274, -0.9467735, -0.2926064, 0.335516, 0.8073883, 1.01572, 
    0.6222305, 0.2053051, -0.6121407, -1.341568, -2.101982, -2.470997, 
    -2.739223, -3.409016, -4.244953, -4.462925, -5.039486, -5.477505, 
    -5.761358, -5.225679, -4.886879, -4.057192, -3.366564, -2.920992, 
    -2.654594, -3.363447, -4.457199, -4.790531, -4.981417, -5.01475, 
    -7.042351, -6.64053, -5.89209, -5.361881, -5.40094, -5.321251, -5.713177, 
    -5.687138, -6.082191, -5.851198, -4.992603, -4.178547, -3.930107, 
    -4.479847, -4.607716, -5.290527, -6.51162, -7.471256, -8.100426, 
    -7.515526, -6.785057, -5.400681, -4.335835, -3.336878, -3.173855, 
    -3.434013, -4.463703, -5.734016, -6.357452, -7.548862, -8.283234, 
    -8.530109, -8.266308, -9.041573, -5.346516, -5.537663, -5.395473, 
    -4.912401, -4.189745, -4.152504, -3.919958, -4.486099, -4.124119, 
    -3.624115, -6.325424, -6.32074, -4.505379, -1.927776, -1.388451, 
    -2.080383, -3.219177, -4.294708, -3.894188, -1.140537, 1.282379, 
    1.584457, 0.3953934, -0.0642395, 0.4391441, -0.2707443, -2.965271, 
    -5.838448, -4.255108, -2.032192, -1.3874,
  -0.9014683, -0.6842804, -0.2486019, -0.1881886, 1.725616, 1.37952, 
    0.9935837, -2.423862, -3.220217, -3.15303, -2.822302, -2.826208, 
    -3.766054, -4.160585, -3.875689, -3.128033, -2.362406, -2.244436, 
    -2.792355, -3.472822, -3.452253, -3.534023, -3.394438, -3.168135, 
    -3.188448, -1.505636, -1.960583, -4.43923, -4.162928, -3.576471, 
    -2.730377, -2.218399, -2.059544, -1.878292, -1.634802, -1.764229, 
    -2.372822, -2.948082, -3.679853, -4.34053, -5.112667, -5.473083, 
    -4.969177, -4.35277, -3.726208, -3.58975, -3.381678, -3.027771, 
    -2.848606, -2.963448, -2.844437, -3.007719, -2.562666, -2.062403, 
    -1.912922, -1.559015, -0.8436508, -0.2540665, -0.4996395, -0.9108391, 
    -1.434019, -1.23402, -1.211363, -1.372564, -1.595999, -2.099125, 
    -2.595478, -2.771257, -2.772816, -2.168911, -1.51318, 0.7800465, 
    0.8222389, 0.750885, 0.2980156, -0.3176079, -0.8850555, -1.924118, 
    -3.080368, -3.825417, -4.641567, -4.584015, -4.015003, -3.154846, 
    -1.906151, -0.9868813, 0.2675438, 0.6928024, 0.9219742, 1.156086, 
    0.9550514, 0.6175499, -1.782452, -1.957458, -1.7085, -1.569435,
  -1.323601, -1.202507, -1.071517, -0.9819336, -0.988184, -1.212142, 
    -1.150163, -1.026204, -0.9816723, -0.9071941, -0.7663078, -0.5897465, 
    -0.3402681, 0.1336908, 0.3792648, 0.3263988, 0.02379417, -0.2311535, 
    -0.3728199, -0.5480843, -0.9780331, -1.385063, -1.778551, -2.087666, 
    -2.538967, -2.87933, -2.923342, -2.672039, -2.431933, -2.284798, 
    -2.189222, -1.965785, -1.704847, -1.597555, -1.374901, -1.084538, 
    -0.8624029, -0.8376617, -0.8626652, -0.782196, -0.5202198, -0.2462616, 
    0.1258736, 0.5467091, 0.8388996, 0.8902016, 0.8758783, 0.6771812, 
    0.3490572, 0.1149435, 0.04619408, -0.1801081, -0.5144835, -0.7082338, 
    -0.8181314, -0.7933931, -0.7142248, -0.5702143, -0.4975586, -0.5736017, 
    -0.5376644, -0.4545898, -0.3595371, -0.3160496, -0.5178719, -0.8337593, 
    -1.074644, -1.155895, -1.253813, -1.348347, -1.104073, -1.012669, 
    -0.9790745, -1.033762, -1.134542, -1.103292, -1.406157, -1.678293, 
    -2.129072, -2.455635, -2.505896, -2.781416, -2.600161, -2.247036, 
    -1.943649, -1.423597, -1.159012, -1.048079, -1.011099, -1.121519, 
    -1.32152, -1.537405, -1.685846, -1.846783, -1.734541, -1.513185,
  -0.486618, -0.5902634, -0.7900028, -0.9972944, -1.107711, -1.090004, 
    -1.108754, -1.093128, -1.094952, -1.055629, -1.068129, -1.088703, 
    -1.113443, -1.045735, -1.008756, -1.009015, -1.056671, -1.054587, 
    -1.050159, -0.9993782, -0.9709949, -0.9551096, -0.9650059, -0.9691725, 
    -0.9329748, -0.936101, -0.9217777, -0.8910494, -0.8551111, -0.7603188, 
    -0.6332359, -0.4295893, -0.2040691, 0.0214529, 0.3047867, 0.554265, 
    0.8326511, 1.054006, 1.234213, 1.43239, 1.599319, 1.745413, 1.837598, 
    1.938379, 2.039941, 2.139421, 2.17666, 2.183431, 2.164942, 2.063378, 
    1.909213, 1.798535, 1.628744, 1.495672, 1.391246, 1.267027, 1.106868, 
    0.9498367, 0.8050451, 0.6206713, 0.4094744, 0.2623386, 0.1118174, 
    0.01077557, -0.07776642, -0.1249027, -0.1819305, -0.2196913, -0.2147436, 
    -0.2475576, -0.3105783, -0.3074532, -0.2853174, -0.2735996, -0.2553682, 
    -0.2587528, -0.2691698, -0.2334948, -0.1866198, -0.1501617, -0.05458832, 
    0.02223492, 0.1347351, 0.2422867, 0.3081713, 0.3313484, 0.3678064, 
    0.3792648, 0.3055677, 0.257391, 0.1805677, 0.1019211, -0.02438068, 
    -0.1777649, -0.2785454, -0.3553677,
  -4.77813, -4.710419, -4.623955, -4.565361, -4.554169, -4.520317, -4.572136, 
    -4.683594, -4.765625, -4.898956, -4.930473, -5.175522, -5.380989, 
    -5.544525, -5.660934, -5.704689, -5.647659, -5.630997, -5.517967, 
    -5.447403, -5.307297, -5.195572, -5.151306, -5.039581, -4.89817, 
    -4.748436, -4.532806, -4.287498, -4.106247, -3.890884, -3.67083, 
    -3.442184, -3.243225, -3.053383, -2.859116, -2.697395, -2.531509, 
    -2.419533, -2.334892, -2.228905, -2.135414, -2.052864, -2.030212, 
    -2.120575, -2.271355, -2.448441, -2.646347, -2.868225, -3.117973, 
    -3.364845, -3.704948, -4.038544, -4.375778, -4.65052, -4.896088, 
    -5.043755, -5.158592, -5.283073, -5.320839, -5.293747, -5.355995, 
    -5.473434, -5.584373, -5.597397, -5.519272, -5.435936, -5.284378, 
    -5.188545, -5.089325, -4.980209, -4.955467, -4.801048, -4.601303, 
    -4.508072, -4.253906, -3.977341, -3.710159, -3.490891, -3.322655, 
    -3.245834, -3.241409, -3.197136, -3.151566, -3.1586, -3.341408, 
    -3.555984, -3.760414, -3.946609, -4.050781, -4.134109, -4.262497, 
    -4.404686, -4.552597, -4.7099, -4.808861, -4.812241,
  -4.484894, -3.756775, -3.302345, -2.79818, -2.444267, -2.333595, -2.486458, 
    -2.666664, -2.861458, -2.980217, -3.134125, -3.21302, -3.353378, 
    -3.57135, -3.872925, -4.084625, -4.265884, -4.477341, -4.697395, 
    -4.723183, -4.713799, -4.71328, -4.777084, -4.662239, -4.502342, 
    -4.346092, -4.243752, -3.984375, -3.725784, -3.479431, -3.386459, 
    -3.603394, -4.046097, -4.417435, -4.815628, -5.295319, -5.788017, 
    -6.257553, -6.533592, -6.618752, -6.549736, -6.507027, -6.422142, 
    -5.995049, -5.346092, -4.333595, -3.482285, -3.386452, -3.793228, 
    -3.978905, -4.264061, -4.738548, -5.034637, -5.044533, -5.209633, 
    -5.898438, -6.348961, -6.230988, -6.453651, -6.577866, -6.61615, 
    -6.341667, -5.998184, -6.086456, -6.207298, -6.390366, -6.410942, 
    -6.598434, -6.633072, -6.176819, -5.700783, -5.398178, -5.18438, 
    -4.770836, -4.289581, -3.466408, -2.860672, -2.1875, -1.830208, 
    -1.708069, -1.680206, -1.560944, -1.960678, -2.515099, -3.086983, 
    -3.256508, -3.398956, -3.720573, -4.304169, -4.82682, -5.455994, 
    -5.822922, -6.037498, -6.144005, -5.642975, -5.059631,
  -1.630203, -1.438278, -1.868225, -2.564835, -3.375534, -3.998962, 
    -4.549744, -4.590363, -4.789063, -5.0336, -5.161987, -5.140625, 
    -5.086456, -5.117447, -5.103378, -4.960938, -4.667969, -4.504944, 
    -4.471344, -4.140106, -3.782028, -3.661987, -3.670822, -4.03125, 
    -4.33255, -4.78125, -5.435944, -5.717194, -5.734909, -5.749207, 
    -5.639053, -5.459381, -5.527084, -6.003906, -6.404953, -6.545044, 
    -6.867706, -6.874481, -6.928391, -7.113022, -7.195313, -6.891937, 
    -6.417976, -6.073692, -5.360161, -4.547394, -4.542442, -5.192444, 
    -5.657288, -5.650787, -5.96328, -5.797661, -5.590881, -5.464844, 
    -5.481514, -5.209373, -4.910416, -3.973434, -3.203125, -2.99688, 
    -3.082809, -3.03125, -3.629173, -4.912758, -6.250526, -7.423958, 
    -7.805725, -8.165108, -8.142967, -7.283852, -5.558594, -3.657806, 
    -1.590889, -0.04244995, 0.4143219, 0.4895782, 0.4760437, -0.1434937, 
    -0.3937531, 0.2304688, 1.253128, 0.8882828, 0.2208328, -0.3093719, 
    -0.6843719, -1.362244, -2.045837, -3.211716, -4.094009, -4.663803, 
    -4.739067, -4.358589, -3.667969, -2.80677, -2.114578, -1.914841,
  -2.411713, -3.240631, -4.381256, -5.128128, -5.401306, -6.108597, 
    -6.672134, -6.944534, -6.969543, -6.889587, -6.945572, -6.54895, 
    -5.981247, -5.786194, -6.428375, -7.354431, -7.787231, -7.446091, 
    -6.832031, -5.838287, -4.9375, -4.496353, -4.283585, -4.639847, 
    -5.080734, -6.157028, -7.079697, -7.228134, -7.587509, -8.445313, 
    -8.824738, -8.457291, -8.181244, -8.302078, -8.487488, -8.952606, 
    -9.607803, -9.603119, -9.10495, -9.011459, -9.438293, -9.752075, 
    -10.34375, -10.73386, -10.84349, -11.66355, -11.2151, -11.78645, 
    -12.45599, -12.06509, -11.00521, -9.073959, -6.704956, -5.148705, 
    -5.125778, -5.037758, -4.50547, -3.802864, -5.309639, -6.626823, 
    -8.570839, -9.953384, -11.53463, -12.26459, -12.83099, -12.67109, 
    -11.93047, -10.89583, -10.09636, -10.07734, -8.971352, -6.27552, 
    -3.813805, -2.723961, -1.297661, 0.4210968, 2.21875, 2.204948, 2.547142, 
    2.916924, 1.682289, 1.923958, 2.117706, 2.526825, 2.799217, 1.20182, 
    -1.107811, -1.846611, -1.49662, 0.4848938, 1.946877, 2.329948, 1.942444, 
    0.5695343, -0.6075439, -1.509109,
  -1.819275, -3.360428, -4.300003, -5.272919, -6.465363, -8.120575, 
    -9.285156, -9.847397, -10.15808, -10.08827, -9.657028, -9.472916, 
    -9.257294, -8.958847, -8.229691, -7.476303, -7.423172, -7.449219, 
    -7.381241, -7.839844, -8.556, -8.432816, -7.217712, -6.543228, -7.328903, 
    -7.956772, -7.58255, -6.993759, -6.976822, -7.604416, -9.078384, 
    -9.704681, -10.23647, -10.24193, -9.849472, -9.386719, -9.10051, 
    -8.853134, -8.984634, -9.846359, -10.24271, -9.903122, -9.715881, 
    -9.401047, -9.327591, -8.549484, -8.242706, -9.294525, -8.948959, 
    -7.449997, -5.260666, -4.579178, -4.332031, -4.789063, -6.515625, 
    -8.034889, -9.376045, -9.289833, -8.587502, -6.998177, -6.918755, 
    -8.607033, -11.73568, -13.71303, -13.50625, -12.26484, -10.19219, 
    -10.22604, -9.848694, -10.33907, -9.742966, -10.61718, -9.601295, 
    -8.765099, -7.781258, -8.104424, -7.530464, -5.199478, -3.680466, 
    -1.34037, -1.608856, -1.077347, -1.826042, -1.755203, -2.234894, 
    -3.637756, -3.724739, -3.559113, -1.880989, 1.641159, 2.548965, 3.700264, 
    3.051559, 1.706497, 1.471603, 0.3364563,
  -4.422394, -4.991928, -4.844803, -5.31041, -4.924225, -4.9375, -5.943497, 
    -6.613541, -7.239853, -7.69426, -8.197662, -9.362244, -9.58699, 
    -8.702866, -8.521622, -8.531769, -6.846878, -5.346085, -6.01355, 
    -6.642181, -6.887238, -6.353653, -5.107819, -4.858597, -6.131775, 
    -7.668747, -8.253372, -7.589584, -8.071609, -8.505981, -9.780472, 
    -11.01666, -10.22475, -8.969528, -8.423447, -7.576569, -6.389313, 
    -6.15834, -5.796875, -4.797394, -4.264587, -4.633072, -4.45546, 
    -4.346359, -2.857803, -2.666656, -2.419281, -0.7880249, 0.3364716, 
    -0.2791595, -0.3999939, -0.6210938, -0.6703186, -1.015884, -2.191406, 
    -5.592972, -8.695053, -11.05833, -11.68645, -11.95625, -11.1125, 
    -11.29869, -12.85469, -12.37187, -10.4474, -8.123962, -8.2789, -10.33411, 
    -12.60573, -13.89687, -14.86537, -14.32162, -11.04271, -8.884109, 
    -8.686981, -9.777863, -10.06172, -7.075775, -3.097397, -3.630989, 
    -5.527084, -6.262238, -6.785156, -7.359116, -7.012756, -6.364319, 
    -6.33255, -7.285416, -5.13855, -3.492188, -2.401566, -3.364838, 
    -4.884384, -4.683853, -3.980988, -3.456253,
  -7.766922, -9.513275, -8.308853, -6.739853, -6.277084, -9.28334, -10.49323, 
    -9.354431, -9.043762, -9.396606, -8.619003, -6.986191, -6.244019, 
    -6.827347, -10.30026, -10.13489, -8.027863, -6.640366, -8.074997, 
    -10.69193, -9.604691, -9.025513, -7.927338, -6.592972, -5.717972, 
    -5.2388, -5.403381, -6.548691, -6.989334, -7.514587, -7.21875, -9.166931, 
    -10.26614, -11.11145, -11.36067, -10.34167, -9.152344, -9.403137, 
    -5.178391, -2.97084, -5.128387, -7.3461, -6.463287, -7.333847, -6.764587, 
    -6.675262, -8.769791, -7.149994, -0.1184845, 5.045837, 3.971619, 
    0.5809937, -0.8734283, 0.6101532, -0.4130249, -2.319534, -1.739578, 
    -1.26796, -4.664322, -8.769791, -11.33749, -12.43567, -11.22527, 
    -9.630219, -7.599228, -6.670319, -10.58646, -13.00261, -12.34088, 
    -13.21198, -13.85182, -17.57265, -19.26953, -18.06094, -16.44479, 
    -15.38698, -13.51772, -13.23776, -13.97839, -12.75365, -12.18491, 
    -12.75157, -9.5961, -6.765106, -5.382553, -6.638794, -11.44037, 
    -13.37709, -10.94583, -10.74062, -10, -9.563278, -9.071106, -7.067703, 
    -6.188538, -6.498947,
  -10.01797, -9.781509, -6.442719, -7.775009, -10.25755, -13.57916, 
    -11.92943, -7.890106, -8.661972, -9.795303, -8.640625, -6.0513, 
    -7.779175, -8.030472, -9.170044, -7.77005, -5.327087, -6.166931, 
    -9.479691, -9.340622, -6.731003, -7.679688, -10.00078, -8.664063, 
    -4.382294, -2.079163, -1.147141, -3.861984, -3.114059, -0.7796783, 
    0.1546936, 2.892456, -2.173965, -5.668488, -6.097137, -10.12968, 
    -11.44246, -13.41589, -12.57527, -12.74583, -11.33411, -9.550262, 
    -11.80521, -12.21303, -12.08541, -10.14687, -9.91954, -9.085403, 
    -4.188797, 0.3835983, 2.734116, 1.754684, 2.501053, 1.574219, 1.848953, 
    2.416138, 1.135162, 0.7294312, 2.457809, -0.3367157, -4.322144, 
    -5.542709, -11.26068, -15.03412, -17.63333, -20.25807, -18.91147, 
    -15.44557, -14.79974, -14.86067, -14.5625, -12.83307, -14.97239, 
    -11.04063, -8.686203, -10.90938, -14.27838, -16.40781, -16.78542, 
    -16.03386, -18.84245, -21.8078, -22.27812, -18.67604, -13.86797, 
    -12.55885, -10.92265, -9.539063, -7.445313, -7.654175, -9.247391, 
    -10.68021, -9.716141, -8.598694, -8.6539, -8.6362,
  -13.53386, -16.07005, -15.97293, -16.31224, -18.91954, -21.73438, 
    -20.29999, -20.70338, -23.26668, -23.18491, -19.73463, -20.39479, 
    -20.91562, -19.75417, -25.52657, -29.64818, -30.09479, -26.57942, 
    -27.89635, -29.81848, -28.38776, -26.17265, -21.8526, -20.02969, 
    -16.66121, -10.55235, -8.016922, -5.3685, -4.925781, -4.498962, 
    -3.550522, -2.471344, 0.3252716, 0.1007843, -2.630478, -5.140625, 
    -7.856247, -8.517197, -10.04141, -11.02475, -9.083847, -5.200531, 
    -0.8158875, -2.470581, -3.308334, -2.103394, -0.006515503, -3.777084, 
    -5.0737, -4.363815, -4.478378, -5.233337, -7.96225, -6.579422, -3.664063, 
    -2.133331, -1.059891, 0.02500916, 0.1664124, -3.639069, -4.438019, 
    -0.9031219, -0.4026031, -0.4570313, -3.5625, -5.533325, -2.949738, 
    -2.479172, -6.103912, -8.594025, -8.774216, -5.135666, -3.983856, 
    -5.965881, -5.529694, -8.611984, -10.63776, -8.840881, -3.742447, 
    -2.75235, -2.183334, -5.612503, -7.186203, -11.23465, -15.78854, 
    -18.33488, -23.30287, -26.98308, -25.28333, -21.1703, -17.42162, 
    -14.86926, -15.64323, -15.53099, -11.62735, -9.792969,
  -16.88515, -13.02057, -13.14583, -10.26198, -2.008865, -4.274994, 
    -9.527603, -8.823959, -10.01225, -4.715881, -1.839844, -3.578644, 
    -5.854172, -4.382553, -1.371353, -2.359894, -4.425781, 0.2705688, 
    2.336716, -3.435684, -8.135147, -8.282288, -6.154953, -4.566666, -1.1586, 
    -2.757278, -4.883347, -2.255722, -0.8244781, -2.415878, -1.691406, 
    -1.291412, 0.6184845, -2.205475, -7.085403, -7.441666, -1.215363, 
    -1.0289, -5.025787, -3.730469, -3.683334, -7.094528, -2.858078, 
    -2.494522, -0.6583252, -0.2770844, -0.8013, -3.657562, -2.91301, 
    -0.06510925, 3.260681, 0.04740906, -5.038269, -3.28125, 0.2322845, 
    3.394531, 4.257553, 2.175522, -0.4299469, -5.807037, -3.66275, -1.803391, 
    -1.13385, -0.4807281, 2.677094, -1.186447, -5.757294, -2.299744, 
    -1.344269, 0.1875, -2.555466, -5.479675, -5.474228, -3.944534, -1.8302, 
    -2.563797, -1.619019, -1.540878, -2.305984, -3.092194, -3.069794, 
    -1.632294, -4.529694, -6.985947, -5.06015, -7.257813, -10.82291, 
    -14.28906, -14.48724, -14.75494, -18.4539, -21.72682, -22.67291, 
    -25.01927, -24.00703, -19.95703,
  2.735153, 3.212753, -1.837494, -1.970581, -1.81694, -5.703125, -5.725525, 
    -1.736969, 0.6387939, -2.161469, -3.615891, -1.1586, 0.0161438, 
    -2.679153, -2.798431, -2.782288, -2.484116, -1.677872, -3.756516, 
    -2.252335, 1.786728, 3.331253, 2.063019, 0.1190033, 0.1005249, -1.3237, 
    0.5276031, -2.680481, -5.642456, -5.110153, -1.463028, 1.297134, 
    -1.440369, -1.553116, -1.225266, -1.380737, -2.983856, -4.048431, 
    -0.9377594, 1.633072, 3.028122, -2.435425, -3.279953, 1.763794, 4.978134, 
    3.559906, 0.0617218, 2.83255, 6.604172, 9.894531, 11.04688, 6.971359, 
    3.661194, 4.863541, 6.347397, 5.944016, 5.272659, 4.598953, -0.9026031, 
    -5.497391, 0.0236969, 2.507813, -1.011444, -0.416153, 2.853134, 3.008087, 
    0.5984344, 1.999222, -1.407562, -4.231522, -5.859634, -2.736984, 
    2.661469, 1.999741, -1.376816, -3.350266, -3.227859, -0.4304657, 
    -1.483597, 0.359375, -0.271347, 1.938278, -0.734375, -3.114319, 
    -1.652863, -1.643494, -3.922653, -3.892441, -1.488541, -2.625259, 
    -3.375778, -3.612762, -6.4086, -9.179169, -5.739838, -2.6922,
  2.982803, -2.087769, -2.720566, -1.935944, 1.322922, -0.07577515, 2.1875, 
    -1.031769, -3.119019, -3.113281, -4.277603, -3.857559, 2.035156, 
    0.1848907, -4.791138, -2.216919, -1.654434, -2.227615, 0.1658783, 
    -2.024734, -2.940353, -5.128128, -4.489578, -3.577332, -2.068481, 
    -0.6364594, 0.8656311, 2.846359, 0.7963562, -0.6244659, 4.335159, 
    6.724991, 6.842712, 2.295059, 1.089066, 1.485672, 0.7273407, 2.860687, 
    6.153381, 6.687241, 2.850266, 5.658081, 5.54245, 4.849213, 5.360153, 
    5.882019, 4.487762, 4.70546, 6.320572, 7.683334, 7.200531, 8.870041, 
    5.284637, 3.579437, 6.132553, 4.033325, -3.946609, 0.8927155, 4.785156, 
    0.08906555, 3.618484, 2.833084, 0.8184967, 2.740616, -0.3036499, 
    -2.423431, -0.7411499, -2.388809, -3.894791, -5.359375, 0.9406281, 
    4.491394, 1.150513, -1.136978, 3.066666, 8.084885, 7.850784, 6.398178, 
    7.502869, 2.655731, 1.288284, 3.777344, 6.742706, 7.999222, 4.937759, 
    3.769012, 1.335938, -1.710419, -1.229691, 0.568222, 1.996872, 0.423172, 
    -0.2533875, 0.6658783, 4.262238, 6.862762,
  0.1484375, -0.4557343, 0.6419373, -0.1979065, 1.435425, 0.9174347, 
    -0.15625, -3.792191, -3.272659, -1.33255, -1.219528, -7.608856, 
    -4.001572, -4.273697, -3.639053, -1.500259, -2.223953, -0.7026062, 
    2.515625, -1.444534, -0.6002655, -1.138809, -0.1046906, 5.076035, 
    8.469009, 8.574478, 4.641403, 4.7323, 6.681519, 4.978378, 2.228119, 
    6.739319, 4.988541, 3.690109, 7.280991, 5.761719, 2.585678, 5.71666, 
    6.396088, 3.63829, 2.353119, -1.541656, 5.361725, 4.086456, 4.134888, 
    4.703644, 8.46875, 5.080475, 4.257034, 3.691147, 8.055984, 9.630997, 
    5.847916, 5.1138, 1.791672, 4.058594, 2.447144, 1.168747, -0.06796265, 
    1.708862, 1.231781, 1.460419, 3.500259, 2.812759, 0.7419128, -3.866409, 
    -1.370575, -1.271881, 0.5966187, 3.832291, 1.577072, -0.2354126, 
    4.469788, 4.635162, 10.61797, 15.91771, 16.68073, 15.50652, 8.171097, 
    2.546875, -1.453644, -0.7747498, 7.985413, 5.809906, 0.5471344, 1.978897, 
    0.5677032, -2.152084, -2.921356, -1.189575, -3.745316, 2.639847, 
    1.370575, 0.2408752, 2.350266, 3.387756,
  2.104431, 3.115097, 2.716675, 2.462769, 5.631775, 0.6739655, 0.0697937, 
    -1.795837, -4.223434, -7.177612, -5.181259, -2.153381, 2.171356, 
    1.136719, -2.650787, 2.640366, 5.076553, 7.133865, 6.711975, 5.029678, 
    12.93802, 11.42188, 6.965622, 9.215118, 9.30365, 11.76172, 10.33853, 
    11.69453, 8.265366, 4.308594, 1.783325, 3.102356, 5.116409, 11.23438, 
    6.136459, 4.002609, -1.654694, 3.512512, 8.939316, 6.429688, -1.895828, 
    -3.257019, -1.67395, -3.19635, 1.775253, 5.296875, 6.435684, 11.4026, 
    3.60495, 4.551559, 9.431244, 8.842453, 5.659897, 3.317703, -2.492981, 
    0.2661438, 4.851303, -1.119019, 0.5723877, 4.142975, 3.714325, 4.533066, 
    3.411987, -1.051559, 1.990891, 1.590881, 2.198441, -2.100006, 1.505997, 
    2.258072, -2.702866, 3.680481, 7.552094, 3.078903, 5.358856, 9.030731, 
    17.50496, 23.58749, 4.069016, -1.077866, 1.487244, 2.837753, 0.1666718, 
    1.732559, 0.7067719, 3.585678, -6.386459, -9.278381, -1.5112, 1.655991, 
    0.6658936, -3.216934, -3.457809, -1.507294, -2.188812, 0.4302063,
  2.83046, 1.494263, 2.164856, 1.557831, 3.807556, 1.129425, 2.693756, 
    -0.4085999, -4.955475, -3.315109, 4.054688, 6.577072, 1.407547, 
    -0.6536407, 7.192719, 5.6427, 2.327606, 7.937241, 9.026047, 7.1185, 
    12.13516, 7.616135, 6.887512, 10.1375, 3.746613, 9.172379, 10.8159, 
    4.304428, -0.2218628, -4.118744, 1.297653, 7.063782, 5.686188, 1.03775, 
    0.07006836, -0.4182434, -1.846344, -0.8247375, 1.798187, -8.365097, 
    -10.65181, -7.214844, -2.517181, -1.294006, 2.390106, 4.55365, 4.276306, 
    8.608078, 10.29688, 7.029678, 5.966919, -1.520569, -5.125778, -3.980469, 
    -6.923706, -4.404434, -0.3372345, -6.322403, -1.205475, 4.865356, 
    1.783859, 0.7414093, 3.77916, 2.366928, -0.954422, 0.7880096, 2.044266, 
    3.824478, 1.431763, -0.2890625, -2.895569, -1.617447, -7.278641, 
    2.781509, 7.1875, 2.516418, 5.967712, 9.641418, -1.873688, -10.9612, 
    -5.816147, -7.761719, -9.649734, -8.49791, -10.86095, -12.74376, 
    -11.33255, -11.84871, -12.62708, -10.15157, -5.146622, -2.685944, 
    -2.178909, -3.609375, -0.3335876, 2.882034,
  -1.508331, 3.148712, 7.8909, 5.413544, 2.52475, 0.3416748, -0.3606873, 
    4.501556, 1.31041, -6.419006, -1.239075, -3.556793, -7.870834, 2.691406, 
    9.165649, 7.534119, 6.880981, 9.55365, 0.1638184, -4.943756, -3.699219, 
    2.711731, 1.982574, -2.431519, -3.873718, -0.3463745, -2.500763, 
    -2.716919, -1.64975, -1.583344, 9.142975, 6.960938, 0.9789124, -6.2677, 
    -4.447144, -3.687256, -0.3999939, -3.88855, -5.832031, -2.797943, 
    -5.690887, -7.224487, -4.979706, -3.044006, 0.0682373, 0.7843628, 
    1.774475, 1.12291, 4.954681, -2.478394, -5.348434, -6.239838, -9.579422, 
    -8.032822, -10.82657, -7.371887, -5.748428, -1.153381, 2.588287, 
    7.451294, 2.951553, 1.573181, 0.5872498, -1.698181, -4.204681, -1.669525, 
    -6.916672, -6.6651, -7.130463, -10.08411, -12.32552, -9.615875, 
    -6.231262, 2.261719, -2.385437, -3.828125, -4.029694, -6.262238, 
    -4.86145, -11.12318, -13.37994, -6.470306, -16.75417, -17.73906, 
    -13.35912, -11.87917, -8.88385, -10.87241, -11.319, -5.067184, -0.910675, 
    5.649216, -0.1481781, -0.6903687, 3.829681, 0.5648499,
  2.461212, -1.368469, 1.502075, 1.27005, -0.5317688, -3.012756, 4.048676, 
    3.434357, -2.213791, -3.427094, -6.746094, 1.242706, 3.655731, 6.699738, 
    11.88907, 4.613525, 7.087769, 1.289063, -1.922394, -3.4935, -11.60754, 
    -7.480225, -8.4263, -9.932037, -8.592438, -5.085663, -4.676819, 
    -2.640106, 0.7479248, 1.093475, 0.7271118, -1.07135, -1.4888, -3.878632, 
    -6.344543, -6.707031, -4.947937, -2.487244, -4.035156, -4.570831, 
    -7.04715, -12.05652, -4.891418, -2.883057, 2.670044, 4.186707, 4.508606, 
    -2.768494, -5.795303, -5.506241, -6.432297, -9.478912, -8.952347, 
    -5.728638, -4.964325, -2.809891, -1.465622, 0.2164001, 1.845047, 
    -2.411453, -4.065369, -7.480728, -9.349747, -12.69766, -15.81224, 
    -11.93333, -10.32813, -13.80182, -10.5125, -7.181244, -7.66745, 
    -5.772659, -0.5257568, 0.1481628, -0.3877563, -2.877594, -8.6745, -10.25, 
    -9.299988, -5.20755, -16.61354, -1.904694, -14.12474, -12.3573, 
    -11.64792, -12.3, -14.90182, -18.4698, -9.62056, -5.399216, 1.594025, 
    -0.991394, -0.933075, 2.3815, 2.0737, 2.499237,
  1.773438, 5.596619, 5.159637, -0.410675, -4.231232, -5.950012, 2.523163, 
    -2.891937, -3.198944, 3.588287, 1.849213, -0.8354187, 4.929169, 9.104431, 
    8.316406, 1.876831, -1.506256, 2.262268, -5.509399, -4.3013, -5.951843, 
    -8.813553, -5.601563, -3.129166, -2.221893, -1.6138, 3.131256, 4.565369, 
    4.642181, 2.08255, -1.980743, -4.276031, -3.22995, -3.564575, -3.972656, 
    -8.897644, -8.459869, -3.2836, -0.2554626, -2.913544, -17.07056, 
    -11.41327, -3.942444, -4.45755, 2.281769, 4.398163, -2.748413, -5.910675, 
    -8.4711, -6.064072, -7.105728, -9.143753, -0.8448029, -4.462234, 
    -0.3526001, 1.432297, -1.079422, -5.395844, -5.086975, -7.853119, 
    -13.4487, -13.38985, -14.59949, -13.65572, -19.11015, -15.91537, 
    -11.48827, -11.28543, -7.352341, -6.468216, -3.005219, 1.575775, 
    -2.635681, -0.631012, -0.2583313, -6.422638, -8.170837, -11.25052, 
    -9.540344, 0.6367188, -6.328644, -2.660156, -4.178391, 0.6070251, 
    -0.2505188, -3.556488, -7.995575, -6.871613, -4.487488, -2.277618, 
    0.640625, 2.337769, 0.1473694, 0.244812, -2.70755, 4.639069,
  3.527588, 1.124481, -4.041168, -4.626587, -6.783325, -2.640869, -0.2854309, 
    -2.583588, 0.1901245, 6.397125, 0.2189941, -6.915894, 2.910416, 29.9659, 
    1.125, 1.239044, -1.979431, 1.177094, 5.595337, 1.952332, 2.610962, 
    -0.678894, 0.4424438, -0.9752655, -2.027863, -0.421875, 2.584625, 
    8.399719, 4.771606, 1.861969, -4.473694, -6.031006, -7.202606, -6.6875, 
    -7.251801, -8.250793, -10.44843, -5.793762, -3.7612, -14.53543, 
    -14.17993, 1.014069, 2.568481, 5.852844, 3.398956, -3.153656, -6.864594, 
    -6.134384, -9.915115, -8.821609, -5.914581, -3.526031, 0.6351471, 
    -3.485153, -4.035934, -5.266418, -6.616928, -10.10938, -10.48672, 
    -14.07005, -16.16978, -16.44949, -16.03595, -12.51666, -12.97108, 
    -11.79713, -6.177094, -5.197922, -5.495575, -2.561462, -0.116394, 
    4.394775, 1.225525, 2.980469, -1.213531, -11.51016, -5.674225, -9.817444, 
    -12.94193, 5.74115, -0.9541626, 4.867447, 0.6979065, 4.6604, 8.846085, 
    16.76277, 4.289825, -4.106506, -5.358063, -5.469543, -3.661194, 
    -2.905731, -0.3195496, 0.9028625, 1.716675, 2.989838,
  -1.402344, -3.070068, -6.4505, -10.41275, -3.016144, 0.03048706, -3.632568, 
    -9.113037, -4.691406, 0.7468872, -1.747681, -7.549744, -5.715347, 
    10.15729, -0.8216248, 5.909912, 2.818481, 3.343231, 2.855743, 3.081268, 
    3.420044, -1.129669, -6.046112, -1.632813, -3.147644, 4.25885, 4.453125, 
    8.122894, 6.655182, 1.790863, -3.870575, -6.701569, -6.217438, -5.939301, 
    -11.01431, -7.480194, -5.08905, -5.242188, -6.249481, -6.623962, 
    1.224457, 0.08828735, 0.9463501, 1.100769, -2.082306, -1.679413, 
    -2.480988, -3.618484, -3.010941, -3.053131, 0.5703125, -3.528641, 
    -6.304428, -2.996613, -5.817993, -5.92395, -6.419556, -5.08725, 
    -3.280701, -10.23178, -10.77237, -12.66797, -11.76434, -7.206512, 
    -6.008835, -3.355728, -6.291931, -2.697403, -1.029953, 3.828644, 
    1.035156, 3.124481, 3.380737, 3.13855, 3.329956, -4.438019, -7.224487, 
    -5.923187, 4.554169, 10.38672, 2.157806, -0.3338318, -1.894531, 
    -2.986206, 18.77396, 25.39323, -7.085922, -6.763031, -10.53047, 
    -8.211456, -4.335419, -5.54921, -0.3591156, 1.280212, 7.554413, 1.833588,
  3.238007, 0.3554688, 0.2294006, -8.402618, -1.677338, 3.703125, -5.265625, 
    -13.80444, -5.42395, -7.0047, 0.2361755, -2.855194, -2.793243, 0.0557251, 
    0.05209351, 4.609375, 2.930725, 0.7447815, 2.315887, 3.643219, 2.1763, 
    -0.002075195, -0.0703125, 3.440125, 1.152893, 2.139587, 0.02474976, 
    4.097137, 5.509094, 1.189056, -1.885925, -5.35495, -5.503632, -6.29895, 
    -7.074738, -7.105713, -4.704956, -6.875519, -5.593231, -4.094269, 
    -9.732819, -4.146362, -4.353149, -0.9205933, 2.301025, 6.258865, 
    6.328125, 7.822144, 4.848419, 0.6393127, -2.384125, -0.0791626, 2.229706, 
    -1.35025, -2.552063, -5.836975, -1.865875, 1.863037, -0.9718628, 
    -4.830475, -6.806763, -5.320313, -1.928375, 0.1729126, 1.123444, 
    -1.777863, 0.3776093, 1.534119, 3.265884, 6.444794, 7.571625, 7.395294, 
    11.14401, 5.9133, -7.186462, -3.782806, 2.191666, 13.47397, 15.78801, 
    0.5908813, 0.3020935, -0.5757751, -3.892731, -1.779419, 7.328644, 
    19.11771, -5.540878, -7.224457, 0.02368164, -3.933319, -1.317429, 
    -1.166412, 2.749207, 1.470825, 4.858597, 1.28125,
  5.783325, -1.050018, 7.857819, -5.574478, 6.985657, 5.577332, -3.722656, 
    -8.217194, -6.459106, -1.908051, 2.993225, -0.8624878, 1.814331, 
    6.924744, 6.372925, 5.723175, 1.298981, 1.335175, -0.785675, 1.339844, 
    -1.105469, 1.949219, 3.152069, -0.3070374, -1.581757, -3.292206, 
    -1.281494, -1.459381, -0.4421692, 0.4125061, -1.389587, -3.448181, 
    -5.909912, -5.397644, -2.778625, -8.488556, -12.70493, -14.29868, 
    -14.49426, -9.367447, -6.140625, -6.931793, -6.576828, -1.380737, 
    9.237747, 12.92188, 15.13463, 13.41121, 13.14609, 7.145035, 0.8117218, 
    -0.1828003, 1.699463, 1.602356, 0.6273499, 1.797638, 2.115356, 1.882568, 
    4.121857, 1.366119, 0.6570435, -1.914063, 2.173431, -2.1922, 3.577591, 
    2.891159, 4.962234, 7.336197, 9.907547, 13.97865, 13.71771, 12.60495, 
    11.69064, 4.421082, -9.8927, 1.505981, 27.67656, 13.50443, -0.4919434, 
    4.74765, 4.284622, -10.08308, -8.102875, -4.905212, -1.4487, 5.772919, 
    12.3138, -8.489838, -1.918213, -0.9260406, 1.64975, 4.863541, 5.698959, 
    6.703918, 6.790619, 8.801056,
  9.594299, 8.067963, 15.27161, 3.540619, 14.17606, 15.09088, 7.092712, 
    -1.00209, -8.555984, -8.764313, 8.736465, 5.690643, 5.049988, 8.116913, 
    11.48697, 14.73149, 8.737747, 7.291916, 1.145569, 3.371368, 4.5047, 
    5.57605, -0.1372375, -5.417969, -2.958313, -6.032288, -7.0289, -12.64063, 
    -5.077362, -2.969788, -2.942444, -2.566132, -5.594269, -7.019531, 
    -1.768738, -1.826538, -13.66406, -19.10729, -19.5789, -13.4539, 
    -2.109131, -2.140366, -3.365891, -1.951035, 3.964844, 10.55208, 5.628372, 
    1.759369, 0.5929718, -6.068222, -5.480469, -7.026031, -3.657806, 
    -3.567963, -2.859375, 2.277863, 3.208099, 3.514832, 6.052887, 7.288818, 
    3.278381, 4.279449, 7.531799, 8.248169, 8.45285, 10.53049, 14.51224, 
    15.55939, 11.10286, 12.80104, 11.99377, 11.13672, 1.7677, 1.056488, 
    -1.288544, 9.850266, 5.702866, -6.594513, 4.147141, 10.2776, -3.744797, 
    -4.213531, -0.06509399, 0.3390503, -1.316681, -1.784637, 8.297119, 
    -2.595306, 1.839294, 3.323425, 2.124725, 4.739838, 5.858078, 6.378662, 
    7.134125, 11.72684,
  4.579956, 7.547119, 1.504425, -3.788544, 5.13829, 15.77657, 3.280731, 
    7.23542, -11.55573, -20.66251, 1.616135, 1.969788, 7.132294, 6.758087, 
    10.21823, 10.49088, 9.265381, 8.191147, 7.733337, 8.412766, 8.285172, 
    3.531525, -0.3486938, -2.308075, -2.471588, -0.1002502, -1.9086, 
    -10.65886, -14.28151, -5.11145, -8.519257, -13.84062, -14.31953, 
    -15.60078, -8.454437, -5.574738, -8.209106, -0.0604248, -7.131775, 
    -8.481232, -0.06614685, 2.147919, -2.165619, -4.569534, -9.158844, 
    -12.69296, -16.17059, -16.80286, -13.85287, -13.31458, -2.971344, 
    0.2992249, 1.662476, 5.677338, 0.9786377, 2.5784, 2.959106, 2.147919, 
    4.008606, 4.680206, 2.722137, 2.522675, 7.297668, 5.145813, 7.414337, 
    7.6586, 6.695557, 10.05496, 6.218506, 5.423187, -4.271362, -6.917175, 
    -13.67136, -16.53622, -8.519272, 9.665375, 6.35704, -1.954437, 17.50598, 
    8.140625, 7.074478, -1.4198, -1.700012, -1.217468, 0.354187, 1.600281, 
    2.842712, -1.040619, -3.513794, 0.1533813, 0.5143127, 4.213531, 6.603912, 
    8.204163, 8.751556, 7.567444,
  -1.587006, 0.1106873, 7.977615, 13.02682, 19.65182, 10.77005, 13.51407, 
    13.97682, -5.722664, -18.76953, -6.295319, 5.519012, 3.482803, -3.679169, 
    -5.460938, -2.405212, -1.704681, -0.9046783, 8.686188, 7.992706, 
    1.050781, 4.091919, 5.835938, 6.167694, 7.050262, 2.982819, 8.320831, 
    -4.622131, -18.62032, -14.20494, -9.063797, -9.379692, -9.004684, 
    -19.23463, -15.80939, -9.37291, -13.63177, -12.21066, -8.050262, 
    -4.027344, -1.464584, -8.241409, -12.24896, -19.18672, -18.77187, 
    -21.14218, -24.6599, -25.54767, -20.65652, -18.48022, -14.7677, 
    -11.90314, -10.68829, -8.929169, -6.758057, -8.986725, -5.440887, 
    -4.660675, -6.579437, -6.323425, -4.386444, 1.180725, 1.662506, 2.939331, 
    2.597656, 0.7479248, -2.123718, -3.444763, -5.101807, -6.111481, 
    -10.86198, -14.35886, -19.64609, -22.73203, -25.59869, 9.855209, 
    32.88881, 8.013535, 8.779953, 17.30521, 4.151825, -2.86615, 6.859375, 
    -1.6492, 0.9924622, 5.112762, 4.594513, 0.4992371, -0.2604065, 
    -0.2713318, 0.6846313, -1.247925, -1.010681, -3.28595, -4.230194, 
    -2.313263,
  7.519531, 8.315094, 9.099213, 12.61093, 14.04582, 13.64011, 14.01692, 
    16.19089, 11.05624, 5.822403, 0.5265656, -0.4445343, -0.5041809, 
    -4.859375, -6.398438, -4.407547, -9.334885, -10.30208, -8.563278, 
    -10.45573, -0.4822845, 5.678894, 10.85364, 10.58282, 7.549225, 3.942963, 
    6.316406, -2.21405, -5.567978, -0.8348846, -2.885941, -0.6315155, 
    -9.441406, -7.472916, -9.552612, -6.967972, -5.961456, -5.544006, 
    -5.055466, -0.5940094, 0.5695343, -2.579941, -11.32864, -10.84271, 
    -7.851563, -9.985153, -6.976563, -10.10886, -11.77838, -14.41849, 
    -15.63516, -13.96771, -13.28984, -12.99583, -11.02943, -7.02475, 
    -3.773178, -4.400772, -3.883865, -3.107559, -4.580734, -5.144531, 
    -2.807816, 3.870834, -0.160675, 2.855209, 1.929688, -1.872147, 3.59375, 
    6.214584, -2.336197, -4.839325, -18.09818, -16.57578, -9.801826, 
    2.617706, 10.55441, -3.589325, 13.83672, 11.21405, 1.343231, -2.569275, 
    4.47345, 2.887497, 5.074203, 6.08255, 4.320831, 2.019531, 3.985931, 
    3.226822, 7.336716, 3.314835, 3.269531, 7.307297, 6.402863, 10.05104,
  3.604156, 3.89035, 2.106247, 6.253906, 3.9953, 1.833847, 0.3453217, 
    4.43959, 4.479431, 11.73672, -6.893478, -10.02762, -10.33723, -17.65495, 
    -3.316147, -3.497131, -10.36484, -16.15962, -16.86928, -16.83907, 
    -5.731522, -2.023178, 4.164063, 11.09244, 6.605469, 7.645584, 8.52005, 
    5.643494, 0.4919281, 3.609116, 5.385941, 0.6666718, -10.3237, -8.945313, 
    -6.78125, -3.080719, 2.160675, -2.161972, 0.3320313, -1.596878, 
    0.3177032, 1.693756, -4.705475, -5.210419, -4.099472, -0.1010437, 
    -3.1073, -3.018478, 1.879944, 2.081757, 0.5250092, 4.512238, 8.807297, 
    15.6026, 16.37761, 18.6599, 14.00912, 10.95755, 6.723434, 8.643738, 
    5.1474, 3.532288, 9.400009, 11.5724, 10.06641, 15.07526, 11.6711, 
    3.472916, 4.602341, 5.627869, -0.1989594, -3.372131, -8.566147, 6.612228, 
    26.85677, 19.04192, 10.01875, 12.58568, 14.14662, 15.99324, 1.397675, 
    3.103119, 4.328369, 7.585922, 9.703644, 1.417191, 1.816147, 3.180984, 
    0.4585876, -2.31926, 0.3859253, 2.089584, 0.0171814, 9.2211, 4.535934, 
    9.697922,
  -5.330444, -6.463562, -5.339325, -1.747375, -1.687225, -1.333069, 
    -2.324219, 0.0802002, 3.710175, 0.6026306, -13.84454, -11.0784, 
    -14.54219, -18.46718, -10.03778, -7.958328, -8.293762, -10.86563, 
    -14.42317, -13.98984, -8.821869, -0.3791656, 10.23515, 12.85027, 
    8.493744, 10.125, 2.75885, 4.5112, -3.031769, 10.70755, 10.49947, 
    6.821365, -2.413544, -2.457031, -9.932541, -5.758072, 0.4505157, 
    3.620041, 6.375519, 4.913269, 1.811447, 0.4471436, -0.4229126, -2.831772, 
    -3.38385, -3.632813, -4.644806, -4.726822, -0.007034302, -1.415375, 
    2.05365, 1.172913, -3.618759, -4.753906, -5.938019, -1.975784, 
    -0.1958313, -2.756256, -4.828384, -2.404434, 0.5002594, -0.5039063, 
    4.366409, 4.447144, 4.463806, 3.252853, -0.454422, 3.451553, -2.695313, 
    -7.556503, -11.82526, -8.088547, 6.694534, 14.06328, 18.25391, 9.640366, 
    0.2901001, -3.062759, 0.9898376, 0.923172, 0.9031372, 0.2406158, 
    2.228638, 4.145844, -3.444275, -2.251572, -2.91069, 1.46225, -4.1026, 
    -0.7752686, -3.566147, -0.5414124, -1.650528, -2.202866, -2.850525, 
    -6.846344,
  -6.736694, -5.840637, -4.811981, -3.677368, -3.985168, -4.241913, -5.0672, 
    -1.901276, -2.57135, 0.4718933, -4.141418, -9.519775, -11.74609, 
    -17.24298, -18.65808, -17.89507, -8.252335, -14.18619, -17.86537, 
    -17.19426, -17.78047, 8.002609, 17.32526, 15.83151, 6.128387, 1.1987, 
    0.9645844, 2.440109, 0.2565155, 9.096619, 6.695053, 4.025787, 4.180466, 
    3.777603, -1.986725, -5.453384, -0.5364685, 1.055466, 1.928131, 3.348953, 
    3.535156, -3.109116, 0.004440308, 0.08358765, 1.234634, -0.07369995, 
    1.916931, 1.097137, 6.849228, 6.276306, 1.345306, 1.5914, 0.03230286, 
    1.67395, -3.029938, -1.059631, 2.333588, 1.672668, -0.5223999, 
    -0.5070343, 1.308075, -3.377335, -2.07579, -1.990372, -0.338028, 
    0.1106873, 1.608597, 1.898178, -3.509888, 2.353378, 4.580734, 10.73254, 
    20.8578, 1.395309, 5.366669, 1.798691, -3.170319, 1.269272, -3.405991, 
    -0.9867249, -3.449219, -4.051041, -0.4255219, -1.581253, -1.942703, 
    -0.6143188, -2.730988, 2.178391, 1.499466, 2.43515, -3.485672, 0.444519, 
    -0.5070496, -0.2166748, -2.189575, -5.608063,
  -3.093994, -3.342194, -3.2966, -2.5448, -2.959625, -2.967194, -4.884125, 
    -4.6315, -3.584625, -2.4552, -2.920563, -6.703918, -9.814575, -10.36588, 
    -14.65079, -12.50208, -13.87317, -14.89114, -20.33568, -17.57864, 
    -16.28749, -6.873947, 5.511719, 11.13905, 3.538284, 1.728897, 5.288544, 
    7.634109, -1.710938, -3.198441, -1.304688, -2.322403, -1.563019, 
    5.780472, 5.670578, 4.456253, 4.316406, 3.905212, -1.616928, -4.420578, 
    1.00209, 0.3940125, 0.7716064, 3.15625, 4.375793, 4.461716, 7.689072, 
    7.07135, 4.648438, 4.532562, 5.104172, 6.804428, 5.72995, -2.460419, 
    -2.233078, -4.787506, -3.508331, -2.522659, 0.9752655, 0.6312561, 
    2.572128, 0.3559875, 1.356522, 0.2679749, -0.1502686, 1.815369, 3.403397, 
    2.278397, 5.504944, 8.944778, 16.76772, 18.48151, 10.16875, -3.808075, 
    -3.381256, -4.461197, -5.322144, -1.467957, -2.099747, -2.172653, 
    -4.298172, -0.228653, 0.7700653, 2.376312, -1.121353, -1.048187, 
    2.857285, 2.21225, -3.251038, 0.2552032, 1.207291, 0.2109375, 0.7521057, 
    -0.3200684, -0.4755249, -1.334381,
  -2.192444, -1.434372, 1.686188, -0.8338318, -0.5697937, -1.211731, 
    -1.131775, -3.027069, -4.369537, -3.895325, -4.546356, -8.565887, 
    -7.313019, -6.626038, -10.35782, -11.64035, -8.761993, -7.418243, 
    -17.81718, -21.49245, -20.2336, -15.84401, -2.847382, 3.859116, 6.205734, 
    1.437759, -4.497406, 8.406509, -0.7015686, -3.902344, 2.827072, 4.460938, 
    4.596863, 3.791412, 5.239838, 2.198441, 2.721344, 6.698166, 3.115631, 
    -0.6979065, -0.5559845, -0.657547, -0.264328, 0.5770874, 3.134888, 
    4.943481, 6.144272, 5.647141, 3.942703, 7.092957, 4.581253, -0.9835968, 
    -1.954422, -7.614319, -5.154678, -4.605728, -3.396622, -5.663803, 
    -2.507813, -2.022141, 0.5434875, 1.482803, 0.2036591, -2.070572, 
    -2.093216, -0.4343872, 3.534103, 4.655457, 14.34245, 10.58542, 6.648956, 
    5.973175, 6.385681, 0.3643188, -5.78595, -4.75885, -3.347137, -1.863281, 
    -3.640366, -1.224487, -1.753647, -3.898178, -1.680222, 0.8859406, 
    -1.506516, 0.5778656, 0.623703, -1.85495, 1.411209, 5.021088, -2.561462, 
    1.292435, -0.02708435, -0.140625, 0.9604187, -1.564072,
  -0.1333313, -0.9195251, 0.441925, 2.939072, 4.240356, -1.056763, -2.038025, 
    -0.8291626, -3.035416, -3.743484, -5.151306, -6.381775, -7.540894, 
    -5.315887, -8.488541, -10.18932, -7.021622, -6.918747, -12.37267, 
    -12.68333, -12.45703, -15.23047, -12.48958, -7.641663, 1.989594, 14.1237, 
    -4.165878, 3.234634, 6.394272, -6.740631, -4.910675, 0.7117157, 4.416656, 
    -0.3351593, -1.704941, 3.8927, 1.659897, 5.90625, 4.603638, 4.733337, 
    4.014847, -2.256516, -5.087769, -3.478119, -0.244278, 2.578903, 2.053391, 
    1.48671, 4.746094, 4.908585, 8.678391, 4.545563, 1.703644, 1.123703, 
    -0.2083282, 0.3486938, -1.813278, 0.2052155, 0.046875, 2.969269, 
    -1.575272, -0.4906158, -2.814056, -1.415115, -5.412491, -4.186203, 
    -3.216934, 1.848969, 9.570831, 9.893753, 3.985413, 5.179169, 3.304688, 
    1.130463, 0.9586029, 6.256256, 5.769012, 1.471359, 0.4606628, -4.579697, 
    -1.920837, -0.0320282, 3.821106, -0.940094, 1.101563, 2.638031, 
    0.02082825, -0.6781311, 1.24791, 2.414322, 2.091156, -2.144531, 3.427338, 
    -0.7145844, -0.2546844, 2.132294,
  6.209366, 4.856781, 3.88385, 0.390625, 2.16745, -0.6536407, 4.278137, 
    5.452087, -1.080994, -1.644012, -4.114059, -3.708862, -5.008591, 
    -5.141922, -6.463547, -10.67838, -8.511459, -7.157547, -10.34895, 
    -10.59166, -8.622925, -9.838531, -15.83046, -17.35156, -17.27083, 
    -11.56432, -13.47318, -5.5336, 4.53334, -0.3916702, -9.416397, -6.974731, 
    0.9640656, -0.01953125, 0.1033783, -0.7606812, -1.613022, 1.773956, 
    4.402863, 4.153641, 3.717453, -2.133591, -6.2612, -2.326553, -1.549484, 
    -1.731247, -0.3473969, -0.03463745, 1.356766, 2.708069, 3.940613, 
    2.324738, 2.422668, 1.37265, -1.599747, 1.624481, -1.494797, 3.222397, 
    -0.1437531, 0.5416565, 0.1231689, -0.161972, -5.433594, -4.695313, 
    -4.895309, -5.794266, -3.525253, -4.089325, 3.407806, 5.534378, 3.805481, 
    8.735153, 6.497131, 7.493225, 6.2211, 4.503632, 2.709381, 4.166672, 
    4.881516, 3.165634, 3.665894, 0.5705719, -0.766922, 4.754684, 4.003387, 
    0.1312408, 3.459106, 6.998444, 3.146881, 3.016663, 2.771622, -2.623688, 
    2.452866, 4.223175, 5.530197, 10.75233,
  10.06615, 16.00365, 19.96432, 6.541412, 1.376831, 2.394791, 6.054428, 
    4.7276, 4.661453, 1.296875, -2.779175, -2.65625, -4.824753, -3.81015, 
    0.8388062, -5.229675, -6.617188, -5.628128, -7.344528, -11.09583, 
    -6.083084, -3.970322, -5.4328, -6.846359, -9.152863, -4.444016, 
    -1.147644, -2.945053, 3.219528, 0.2440033, -5.420837, -5.731262, 
    -3.665115, -3.21225, -1.584106, -4.619522, -2.811462, -3.393219, 
    1.483856, 3.694016, 2.699738, 2.548691, 1.893494, 1.389832, -0.9549561, 
    -2.842972, -2.076309, -1.962494, -1.954697, -3.576828, -4.750259, 
    -0.3192596, 3.039581, 0.3627625, 1.170319, 4.785416, 2.3974, 3.234894, 
    4.046875, 4.949219, 3.753647, 2.158066, -2.458603, -5.148178, -6.184631, 
    -5.008331, -4.614853, -2.403122, 1.014328, 0.8781128, 1.932541, 2.487762, 
    1.378128, 1.350266, -0.8940125, 3.177078, 1.109116, 2.116409, 4.036972, 
    3.523178, 7.184113, 4.85704, 2.169006, 5.583862, 4.173172, 5.933075, 
    5.194794, 3.91301, 1.284378, 5.484894, 6.385941, 4.394012, 0.3955688, 
    -1.565369, 3.705215, 8.282028,
  7.922653, 8.943222, 6.570313, 3.541153, 1.597137, 5.839584, 11.45677, 
    8.050522, 8.103653, 9.887238, 2.110672, -0.376297, -4.598709, -3.00444, 
    -0.6716156, -2.380722, -4.072144, -2.369263, -2.33699, -4.283859, 
    0.4580841, -5.734116, -7.203125, -5.530731, -5.923691, -6.206253, 
    -1.414063, -5.296616, -8.358856, -6.421616, -6.772385, -6.71225, 
    -3.146866, -3.598434, -5.871613, -4.335419, -2.683334, -0.576561, 
    1.77475, 4.240616, 5.443748, 5.985161, 2.88855, 2.009903, 1.989059, 
    0.6945343, 0.4372406, 2.051041, 3.877602, 2.417969, 3.019012, 4.625252, 
    0.9648438, 0.3111877, 0.2588501, -0.6020813, 0.690094, 2.35025, 2.024475, 
    0.6437378, 0.2747345, -1.160156, -2.046875, -10.38124, -11.83229, 
    -6.961975, -6.123962, -6.291138, -4.007034, -0.666153, -2.580215, 
    -1.433319, 0.1203156, 2.166672, -1.425003, 2.352859, 4.024216, 0.8408813, 
    0.4458313, 2.866669, 2.549728, 6.151825, 7.053131, 6.646088, 6.206512, 
    5.129684, 4.79895, 5.050522, 3.410416, 0.9684906, 2.779953, 4.974487, 
    3.485153, 1.545303, 2.675781, 5.230194,
  8.626045, -1.273178, 0.8614655, 7.405991, 5.144272, 10.19349, 17.73229, 
    11.58906, 8.817711, 9.615372, 8.612762, 8.833336, 7.267967, 2.197403, 
    3.944016, 4.516159, 2.187759, 1.902084, 0.8661499, -2.480728, -0.7463531, 
    -2.454422, -4.993744, -6.226044, -6.696869, -5.731506, -7.339584, 
    -6.417709, -11.19583, -11.36095, -8.087494, -8.990875, -9.850006, 
    -9.190353, -7.647133, -9.387756, -5.687241, -1.128906, -0.08203125, 
    -6.570053, -7.321877, -3.449478, -1.396873, -5.274216, -3.909637, 
    -0.04348755, 3.168228, 0.9705734, 0.3544235, 0.9833298, 1.666672, 
    1.622131, 1.874474, 3.026299, -1.079163, -3.665359, -1.527077, 
    -0.3315125, -0.5523453, 1.025261, -0.373703, -2.620308, -4.252342, 
    -6.816673, -10.02917, -11.77006, -8.415359, -6.125, -5.305206, -5.260666, 
    -2.481766, -3.082031, -1.352341, -2.401558, -1.786713, 1.827087, 
    1.095306, -2.017448, -2.755203, -2.423706, -4.74688, -1.615623, 
    -1.646095, 0.3979187, 2.402344, -0.2434921, 1.703903, 1.62735, -1.473961, 
    -5.378647, 0.5408859, 3.109116, -2.408325, -1.129684, 0.3419266, 6.138802,
  4.197922, -1.269791, -0.657547, 3.11927, 4.570313, 7.251823, 12.69844, 
    11.3487, 7.470314, 10.47656, 9.802605, 6.228386, 4.209373, 2.336723, 
    2.326294, 3.195313, -0.4549561, -1.4552, -1.0578, -4.449997, -4.735161, 
    -4.296608, -5.784897, -6.277855, -5.429169, -5.282555, -2.950775, 
    -2.942444, -3.874222, -4.623955, -4.456772, -7.024734, -7.35807, 
    -4.409897, -5.437767, -6.634636, -5.728127, -4.324738, -1.197395, 
    -2.263016, -7.010414, -7.518753, -2.867188, -3.536461, -4.04583, 
    -4.795837, -2.437759, 0.5085907, 1.514061, 4.003906, 3.620316, 1.069794, 
    3.196869, 4.281509, 0.4763031, 0.5572968, 2.202347, 4.505203, 3.225258, 
    0.5658875, -1.652603, -0.8682327, -4.622917, -7.647659, -8.893753, 
    -10.90625, -6.469788, -5.521347, -7.023438, -5.919792, -2.575516, 
    -0.6348953, -1.901558, -0.5700531, 0.5570297, 0.3294296, -3.4888, 
    -2.964325, 3.701042, -0.7638016, -3.092712, -3.842445, -3.507034, 
    -6.074738, -4.772141, -6.444016, -5.420578, -0.9028625, -3.096352, 
    -8.119797, -6.859634, -5.337761, -3.495316, -1.21563, -0.4411469, 5.148438,
  0.5302124, 1.570835, -1.148697, -0.33255, -1.123436, -1.88932, 2.190361, 
    5.272141, 4.648438, 5.71067, 4.735931, 4.155991, 3.204681, 3.157814, 
    0.3028641, -1.020836, -1.046608, 1.296616, 0.714325, -0.765625, 
    -3.525002, -4.310158, -5.144791, -6.041924, -3.910934, -0.2070313, 
    0.5299454, 0.981514, -0.7625046, -4.072914, -5.901039, -2.279945, 
    -2.963539, -5.020309, -6.011978, -4.058334, -3.85807, -5.160675, 
    -4.054688, -0.05911255, -2.813278, -4.6362, -1.751305, -1.08802, 
    -2.341408, -1.702866, -1.521873, -1.477348, -2.334373, -0.4028625, 
    0.6367188, 0.3796844, 2.55938, 3.994789, 3.757294, 1.715103, 0.1640625, 
    1.117706, 1.471092, -2.142708, -0.3945313, 2.071358, -2.167969, 
    -4.820313, -7.02578, -5.461197, -7.210678, -6.25, -5.221352, -0.7575455, 
    1.021355, 0.3466187, 0.9635468, 1.908333, 2.244789, 2.314323, 1.389843, 
    -2.283596, -1.949219, -0.6075516, 0.8869781, 2.122917, -3.045319, 
    -1.996094, -1.206772, -2.382286, -0.09557343, -0.6999969, -1.114067, 
    -2.549744, -1.213547, -0.6812439, -1.27578, -2.292969, -3.541145, 
    -1.397659,
  -2.407291, -2.885933, -3.172394, -3.146873, -0.3442688, -2.305729, 
    -1.408596, -0.1671867, 0.955471, -0.9588547, 3.077866, 5.483593, 3.06823, 
    1.375523, 1.099998, 1.551823, -2.181767, -3.029945, -3.496353, -2.425781, 
    -3.83984, -5.196873, -3.827084, -1.58255, -0.2658844, 0.1132813, 
    -0.5249977, -0.5578117, 0.4088554, -0.004951477, -2.54974, -3.975262, 
    -3.773178, -3.694794, -3.646355, -2.486458, -0.4375, -0.4562454, 
    0.6773453, 1.376297, 0.2960892, 0.6325531, 2.922916, 1.603912, 0.0700531, 
    -0.4796906, -1.222393, -3.389328, -1.724998, -0.4799461, -0.7515602, 
    -1.396355, -2.918488, -1.179951, 1.678387, 1.802601, 1.204426, 
    -0.4403648, -0.1583366, 0.1697922, 3.12656, 2.666927, -1.076302, 
    -4.254688, -5.99453, -6.312244, -5.746353, -5.067963, -3.148438, 
    -2.021355, -1.718491, -1.191406, 1.208851, 1.257813, -2.182293, 
    -2.377605, -1.045052, -3.091404, -3.030209, -1.253906, -0.5343742, 
    -0.1304626, 0.5460892, -0.6557312, -1.297653, -2.79974, -3.385677, 
    -3.829166, -0.9783859, 0.795311, 1.864845, -1.493752, -1.645832, 
    -1.421616, -3.667969, -2.955471,
  0.8830719, 1.854687, 0.9945297, 0.1283875, -1.033855, -1.108852, -1.445572, 
    -0.5736961, -0.4364586, -1.102604, 0.4786491, 1.631252, 0.3406258, 
    -1.059635, -0.4377632, -0.01380157, -0.5687485, -0.6653671, -1.009636, 
    -1.85495, -4.04401, -3.623959, -2.014324, -3.374218, -3.687759, 
    -1.990887, -2.772396, -4.048176, -5.382813, -4.595051, -3.770832, 
    -5.485416, -6.980991, -4.467968, -4.427345, -5.692711, -4.101563, 
    1.425259, 4.746353, 5.539845, 2.701042, 0.3031273, -0.8494797, 
    -0.05989456, 2.396091, 1.70026, -1.239582, -2.539063, -2.032291, 
    -0.9184914, -1.088543, -0.3187485, 0.2247391, -1.334892, 1.209377, 
    0.7677078, -1.177341, -0.3981781, 0.2229195, 0.9749985, 1.089323, 
    0.9143238, 0.005207062, -3.417187, -3.939846, -2.716148, -2.594532, 
    -1.953907, -1.363544, -0.8531227, -2.172657, -2.826824, -1.497135, 
    -1.511456, -1.234638, -0.8442726, -4.043751, -4.110676, -2.560677, 
    -4.284374, -1.29427, -1.301823, -2.747398, -1.323959, -3.771873, 
    -3.341663, -2.708073, -2.432293, -1.578125, -1.848179, -2.491405, 
    -2.990364, -1.429169, -0.2898445, -1.158073, -1.182289,
  -0.8013, 0.6083298, 0.7682285, 0.2278652, -0.1221352, 0.4286423, 0.1843758, 
    0.9041672, 1.101042, 0.8598957, 1.231771, 1.714323, 1.35026, 0.9122391, 
    0.3208332, 0.3471355, 1.372395, 1.192709, 0.5908852, -2.352865, 
    -3.362499, -1.514063, -1.368229, -3.139843, -5.067188, -4.254166, 
    -2.805729, -5.202866, -7.394531, -5.546873, -2.762501, -3.008335, 
    -4.152344, -4.132549, -3.827343, -3.305992, -2.571095, -1.513805, 
    -0.8177071, 0.2260399, -1.505466, -6.253647, -7.135159, -4.078384, 
    -2.308853, -1.06979, -0.6690102, -0.9578133, -0.4476585, 0.1664085, 
    0.1072922, -0.8885422, -1.878647, -2.49427, -4.070572, -3.845053, 
    -3.248697, -2.733854, -1.595053, -2.440886, -1.258856, -0.2645817, 
    -1.724739, -3.467709, -3.830469, -3.063801, -1.999218, -1.025257, 
    -1.966928, -2.00703, -2.287239, -2.506248, -3.505989, -5.878384, 
    -5.224998, -3.865887, -5.418489, -5.070572, -1.746616, -0.71875, 
    -0.1786461, -1.410679, -2.122917, -2.715885, -2.761719, -2.263802, 
    -1.733334, -2.133854, -1.760677, -1.030991, -1.074738, -0.4625015, 
    0.671093, 1.255207, 1.519531, 1.160679,
  1.734114, 2.418751, 1.209375, -0.5559902, -1.585938, -1.219271, 
    -0.08176994, -0.1882801, -0.6729164, -1.198959, -1.376562, -0.7895832, 
    -1.525001, -2.026822, -2.21849, -2.000259, -0.7908859, -0.3427086, 
    -0.9026031, -2.959114, -3.48698, -3.801041, -4.035156, -4.237501, 
    -4.846354, -4.426823, -3.683594, -4.577604, -4.53203, -2.807812, 
    -1.373959, -1.093229, -3.460678, -4.75625, -4.295834, -2.740364, 
    -2.55625, -3.350521, -4.592449, -4.554688, -4.367188, -4.901302, 
    -5.155468, -5.70573, -4.977865, -4.254427, -3.96875, -3.900782, 
    -4.147917, -2.288542, -0.9476566, 0.5721359, -1, -2.797136, -2.789845, 
    -2.877604, -2.480469, -1.78776, -0.5544281, -1.054428, -1.842449, 
    -1.174219, 0.2260418, -0.8502617, -0.7856789, -1.174217, -2.169271, 
    -2.037241, -2.536718, -4.429167, -4.485416, -3.984375, -2.659115, 
    -2.450001, -3.30547, -3.604689, -3.094271, -2.913801, -1.877083, 
    -1.355989, -0.8703117, -1.609636, -1.372396, 0.4356766, 0.21875, 
    0.4075546, 0.4354172, 0.2361965, 0.3367176, -0.0007820129, -0.3804684, 
    -0.9252605, -0.4755211, -0.2911453, -0.1549473, 0.7559891,
  -0.1101551, 0.03802109, 0.01223946, -0.6210938, -1.858593, -2.126303, 
    -2.151042, -1.633333, -1.218229, -1.668229, -1.123177, 0.01640511, 
    1.158333, 1.377344, -0.04166603, -0.7453117, -0.8953123, -1.597396, 
    -1.561979, -1.649479, -1.820052, -1.876563, -1.965364, -2.052864, 
    -2.367448, -2.460938, -1.953646, -1.745573, -1.827865, -1.865886, 
    -1.712761, -2.338802, -3.896355, -3.382552, -2.185157, -1.770311, 
    -1.529948, -2.639322, -3.189844, -4.661198, -4.740104, -4.14948, 
    -3.288542, -2.820834, -3.130467, -2.781511, -2.866146, -3.086458, 
    -2.675261, -3.03125, -0.7861986, -0.4617195, -0.7695313, -0.6591148, 
    -1.318229, -1.478126, -1.276823, -0.6940098, -1.146874, -0.9000006, 
    -0.4453125, -0.9765625, -0.9825516, -1.588802, -2.334635, -2.865885, 
    -3.045312, -2.315104, -1.809115, -2.12422, -2.426043, -2.087501, 
    -1.03125, -0.645052, -0.7588539, -2.638803, -0.8302078, -0.7377605, 
    -0.02968788, -0.6713543, -0.8395844, -0.1559906, -0.5309887, -0.5848961, 
    -0.4664059, -0.5523453, -0.6893215, -0.5041656, 0.3796883, 1.017189, 
    0.9421864, 0.2213535, -0.3104172, -0.8848953, -1.449479, -0.8864584,
  -0.5361977, -0.6726561, -0.6398439, -0.7867184, -0.8299479, -0.567708, 
    -0.129427, 0.1924477, 0.008853912, -0.2679682, -0.1695318, 0.009114265, 
    0.4242191, 0.5341144, 0.2182293, -0.2106771, -0.5593748, -0.8627596, 
    -1.117448, -1.240365, -1.359895, -1.695573, -2.158334, -2.277083, 
    -2.117708, -1.62474, -1.220052, -1.028125, -0.667448, -0.4893227, 
    -0.7338543, -0.6239581, -0.1447916, 0.0489583, -0.09713554, -0.703125, 
    -0.5908852, -0.5645828, -0.6067705, -1.049219, -2.123438, -2.555208, 
    -3.136198, -3.209636, -3.461979, -3.153646, -3.294532, -3.56927, 
    -3.21849, -2.573698, -2.202084, -2.036979, -1.90625, -1.669531, 
    -1.779687, -1.70599, -1.419271, -1.047136, -0.9572916, -1.15651, 
    -1.447657, -1.626042, -2.170572, -1.733854, -1.890885, -1.907552, 
    -1.792708, -1.43151, -1.206771, -1.285417, -0.6065106, -0.01848888, 
    -0.07474041, 0.04218769, -0.3419266, -0.585156, -0.4343753, -0.598958, 
    -0.0427084, -0.1424484, 0.03229141, 0.2635422, 0.1575527, -0.07578087, 
    -0.7289057, -1.978386, -2.599479, -2.591667, -1.782291, -1.121615, 
    -0.6932287, -0.3937492, 0.146615, 0.5809898, 0.1026049, -0.2322922,
  0.2010415, 0.1429687, 0.1291671, 0.2080731, 0.1531253, 0.0958333, 
    0.08098936, 0.1039066, 0.05442715, 0.03437471, -0.006771088, -0.04166651, 
    -0.0999999, -0.3203125, -0.3476563, -0.3713541, -0.3450522, -0.4921875, 
    -0.4929686, -0.340625, -0.3252602, -0.2882814, -0.1682293, -0.04583335, 
    -0.04296851, -0.0114584, -0.2463541, -0.4307292, -0.5755208, -0.514323, 
    -0.4507813, -0.4945312, -0.3289065, -0.2059894, -0.1752605, -0.3096352, 
    -0.4356771, -0.5244789, -0.5557289, -0.6447916, -0.539844, -0.2927079, 
    -0.3023438, -0.4572918, -0.5546873, -0.5895834, -0.6312499, -0.6455727, 
    -0.5367188, -0.1781254, -0.1247396, -0.191927, -0.2710938, -0.3742189, 
    -0.3533854, -0.4361978, -0.5393231, -0.6184897, -0.7953124, -1.008073, 
    -1.172656, -0.9648438, -0.8914061, -0.8424478, -0.8242188, -0.5515628, 
    -0.8554688, -0.9041667, -0.8187499, -0.5252602, -0.3617189, -0.1682291, 
    -0.04348969, -0.1338542, -0.3130207, -0.5174479, -0.1664062, -0.0609374, 
    0.03776073, -0.06510401, -0.02265596, -0.0604167, -0.08776045, 
    -0.3083334, -0.3145838, -0.3031249, -0.5049477, -0.8789063, -1.014062, 
    -1.14427, -1.151823, -1.177083, -1.088542, -0.599479, -0.1283855, 
    0.1299479,
  -0.1846354, -0.1945312, -0.1919271, -0.1744791, -0.09140623, -0.1148437, 
    -0.115625, -0.1825521, -0.1466146, -0.1122396, -0.1171875, -0.1351562, 
    -0.1239583, -0.1052083, -0.0986979, -0.1229166, -0.1109375, -0.1156249, 
    -0.0859375, 0.04843748, 0.0817709, 0.04270828, -0.02786458, -0.08229172, 
    -0.1039063, -0.07369792, -0.1216145, -0.2507812, -0.2861979, -0.3148437, 
    -0.3041667, -0.2770833, -0.251302, -0.25, -0.2492187, -0.2856771, 
    -0.354427, -0.4085937, -0.4286458, -0.4476563, -0.3263021, -0.1960937, 
    -0.08697915, -0.03229165, 0.0382812, 0.09973955, 0.1377604, 0.1747396, 
    0.1898437, 0.1960938, 0.1919271, 0.1507812, 0.07682288, -0.003385425, 
    -0.1117188, -0.1127604, -0.09609365, -0.03151047, 0.03932297, 0.06093752, 
    0.1135417, 0.1020833, 0.09609377, 0.0002604723, -0.1557292, -0.3841145, 
    -0.5283854, -0.5916666, -0.5934896, -0.6083335, -0.4921874, -0.3054687, 
    -0.2372396, -0.1526041, -0.05937493, -0.03645825, -0.01718748, 
    -0.06901038, -0.1539062, -0.1669271, -0.2497395, -0.2992188, -0.3473959, 
    -0.3591146, -0.3786459, -0.4195311, -0.4473958, -0.4119792, -0.3041668, 
    -0.1695313, -0.1083333, -0.1497395, -0.2359375, -0.1953125, -0.1789062, 
    -0.1760416,
  -0.03281251, -0.04479167, -0.0546875, -0.06119791, -0.06041665, 
    -0.06328124, -0.06197916, -0.05026042, -0.03151041, -0.009375006, 
    0.006510407, 0.01458333, 0.01822917, 0.01380208, 0.003645837, 
    0.001562506, -0.005208343, -0.009375006, -0.006770834, -0.008072913, 
    -0.01640625, -0.02838542, -0.03776042, -0.05651042, -0.06614584, 
    -0.06848958, -0.07005209, -0.06458333, -0.05546875, -0.04739584, 
    -0.03203125, -0.02682292, -0.02057292, -0.01770833, -0.0234375, 
    -0.02135417, -0.02005209, -0.02526042, -0.02187501, -0.03411458, 
    -0.04244791, -0.04479167, -0.04453124, -0.03229167, -0.03020833, 
    -0.02526042, -0.02317709, -0.02447917, -0.02395833, -0.02395833, 
    -0.0296875, -0.03776041, -0.05182292, -0.06171875, -0.065625, 
    -0.05859375, -0.05833334, -0.05104166, -0.05182292, -0.05260417, 
    -0.06588542, -0.06796876, -0.05572916, -0.05572917, -0.05390625, 
    -0.0484375, -0.04843751, -0.05677083, -0.05729167, -0.06588541, 
    -0.07682292, -0.08281249, -0.07187501, -0.07343751, -0.08229166, 
    -0.08776042, -0.09114581, -0.1010417, -0.1065104, -0.1088541, -0.1140625, 
    -0.09999999, -0.09140624, -0.08854169, -0.08385415, -0.07057291, 
    -0.04869792, -0.04531249, -0.03932291, -0.03098957, -0.01875, 
    -0.01302083, -0.02135417, -0.02473959, -0.028125, -0.02838542,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -9.15625, -9.5672, -9.820313, -10.01511, -10.21875, -10.21304, -10.15601, 
    -10.18802, -10.25366, -10.4039, -10.61249, -10.89246, -11.29401, 
    -11.5354, -11.75076, -11.8685, -12.01303, -12.09402, -12.29843, 
    -12.56485, -12.77707, -12.8862, -12.77316, -12.625, -12.68176, -12.69403, 
    -12.85104, -12.9599, -13.18463, -13.40625, -13.75937, -14.09036, 
    -14.37628, -14.54868, -14.41534, -14.27213, -14.16925, -14.04453, 
    -13.83618, -13.5867, -13.29584, -13.02814, -12.79401, -12.73383, 
    -12.67633, -12.6875, -12.72604, -12.64273, -12.56796, -12.58334, 
    -12.74506, -12.9138, -13.2341, -13.50418, -13.74583, -13.76535, 
    -13.75964, -14.06564, -14.52344, -15.21692, -15.89609, -16.17526, 
    -16.27109, -16.40288, -16.41144, -16.22865, -16.01431, -15.51797, 
    -14.89374, -14.16797, -13.47003, -12.72003, -12.00522, -11.13049, 
    -10.54688, -10.0224, -9.413269, -8.770325, -8.170593, -7.367462, 
    -6.679169, -6.377869, -6.142456, -5.94635, -5.742706, -5.6828, -5.735687, 
    -5.943237, -6.253387, -6.442169, -6.754181, -7.136719, -7.583862, 
    -7.949738, -8.293732, -8.777863,
  -11.09323, -11.28204, -11.55341, -11.74429, -12.04739, -12.41666, 
    -12.92398, -13.43256, -13.72134, -14.05338, -14.71979, -15.30103, 
    -15.6315, -15.86017, -16.01276, -15.90286, -15.82578, -15.69608, 
    -15.60208, -15.46927, -15.45651, -15.30704, -15.12866, -14.72604, 
    -14.11667, -13.62814, -13.28357, -12.87943, -12.32449, -11.66901, 
    -11.36432, -11.64063, -11.90182, -11.6893, -11.36667, -11.04819, 
    -10.10886, -8.762756, -7.0065, -4.950806, -3.062225, -1.5047, 0.3323059, 
    2.036987, 3.088806, 3.880463, 3.922928, 2.978897, 1.997147, 1.163803, 
    -0.06015015, -0.9221344, -2.014328, -3.628387, -4.630981, -4.281509, 
    -3.316925, -2.067703, -1.615891, -1.147644, -1.352615, -1.534119, 
    -2.158081, -3.61171, -5.203644, -6.963547, -8.402878, -9.627609, 
    -10.03436, -10.21223, -9.716934, -8.331253, -5.560684, -2.528381, 
    -0.2346497, 1.434906, 3.690887, 5.05365, 6.272919, 7.546082, 8.591919, 
    8.820038, 8.208069, 6.866669, 5.887238, 4.912994, 3.427612, 1.510956, 
    -0.210144, -2.184387, -4.395294, -5.773193, -7.329163, -8.819794, 
    -10.26877, -10.79764,
  -15.0607, -14.66354, -14.00546, -13.20886, -12.74844, -12.41614, -12.23856, 
    -12.63724, -13.3302, -14.45337, -15.52316, -16.3508, -16.79895, 
    -16.43021, -15.52969, -14.63177, -13.68256, -13.28775, -12.71588, 
    -12.25989, -11.32968, -10.34921, -10.36511, -10.73959, -11.46692, 
    -12.44141, -13.65393, -14.33752, -14.36746, -14.29739, -14.07083, 
    -13.78229, -12.99011, -11.55182, -10.2742, -8.733612, -7.878906, 
    -6.443481, -5.1987, -4.529419, -3.832031, -2.131256, -1.506226, 
    -1.976807, -2.744293, -3.164307, -4.207809, -6.159897, -7.331772, 
    -9.648178, -12.06017, -12.90703, -12.84999, -11.49739, -10.56119, 
    -8.369797, -4.936203, -3.646088, -3.098694, -2.055222, -2.323685, 
    -3.495316, -6.509628, -9.640884, -11.69896, -12.9823, -13.43489, 
    -15.41614, -17.01094, -17.64401, -16.2883, -13.09583, -8.965378, 
    -6.376816, -4.263016, -1.58725, 1.068237, 4.668503, 9.691391, 14.79715, 
    19.03543, 20.65208, 19.05833, 16.29088, 14.80106, 12.61459, 10.03775, 
    6.051559, 2.868484, -0.333313, -3.595581, -7.664063, -11.5914, -13.53333, 
    -14.28021, -14.57446,
  -11.73672, -9.508606, -9.126038, -9.636993, -9.865875, -10.04349, 
    -10.82083, -11.98749, -11.9039, -12.07916, -12.80991, -13.21536, 
    -13.30313, -13.37161, -12.9263, -12.34451, -11.8367, -12.44818, 
    -11.86771, -10.44061, -9.410156, -9.483612, -9.325531, -9.241913, 
    -9.744537, -10.58124, -11.1875, -11.61353, -11.52762, -10.72916, -8.5755, 
    -7.049225, -6.38385, -6.319794, -6.610413, -7.423187, -9.066162, 
    -10.37085, -9.869781, -9.066406, -8.3013, -8.147675, -7.678131, 
    -8.224731, -9.493225, -8.665375, -7.571869, -8.438538, -7.195313, 
    -6.073959, -5.385681, -6.532822, -6.550522, -6.734116, -5.933075, 
    -3.421356, -0.8114624, 2.346878, 1.129425, -1.062759, -1.602081, 
    -2.194534, -5.220322, -9.261978, -13.26511, -15.04428, -18.22475, 
    -18.67891, -16.62057, -15.37682, -14.63672, -14.05469, -13.61797, 
    -13.94765, -15.10599, -13.12083, -5.777878, 3.401047, 10.27344, 15.64505, 
    14.43097, 15.79532, 13.02682, 7.813019, 3.065094, -1.775528, -4.11145, 
    -4.066132, -3.869812, -2.021622, -2.896088, -5.835938, -9.5289, 
    -11.04062, -12.93463, -13.0961,
  -10.05469, -8.686462, -8.989349, -8.683075, -7.379944, -6.583588, -6.87265, 
    -7.053925, -8.208069, -10.34714, -12.40497, -13.50391, -13.66745, 
    -14.67059, -15.01041, -13.95572, -12.36121, -9.378387, -7.568481, 
    -7.925781, -9.405731, -10.41251, -10.0289, -8.289581, -7.159912, 
    -7.414856, -9.385406, -11.92606, -13.51352, -14.68359, -14.09454, 
    -12.26251, -10.81824, -9.943756, -9.623169, -10.02109, -8.770844, 
    -7.539337, -5.939331, -4.076294, -3.197388, -3.376312, -1.844788, 
    -0.3778687, 0.0619812, 0.5023499, -2.126556, -5.404434, -8.33046, 
    -9.08255, -7.70546, -8.349487, -9.469269, -11.11172, -10.89192, 
    -8.047913, -4.020828, -1.270844, -0.9658813, -3.143753, -5.659378, 
    -6.969543, -7.232544, -6.748703, -8.104935, -10.09532, -12.72188, 
    -14.71719, -14.51353, -14.08827, -15.27448, -14.56979, -14.58046, 
    -13.27527, -11.99428, -9.005722, -4.318222, 2.734116, 4.937241, 6.038803, 
    3.647141, 2.006256, 1.653656, -0.4778595, -3.27681, -5.481506, -5.180725, 
    -4.407562, -5.499222, -7.056488, -8.939331, -8.688553, -9.629166, 
    -11.69037, -12.79504, -12.46432,
  -11.75912, -11.83698, -8.271088, -7.11145, -7.632294, -6.740112, -5.87915, 
    -7.364319, -11.75754, -14.44089, -14.23462, -15.87265, -16.89349, 
    -17.74921, -15.32578, -12.44662, -10.16174, -8.069794, -7.186188, 
    -7.947113, -10.4198, -9.667206, -7.941406, -9.524475, -12.84167, 
    -15.19714, -15.63776, -15.77161, -16.59061, -17.78671, -17.77994, 
    -14.48959, -10.46564, -9.532013, -8.658844, -6.609131, -4.272125, 
    -3.029694, 0.08282471, 2.889587, 3.438538, 1.533325, -1.386963, 
    0.6023407, 2.5336, 4.777344, 4.739563, 0.8000031, -3.216919, -6.683075, 
    -4.713806, -2.221344, -0.8585968, -2.730469, -3.422134, -3.619263, 
    -6.193481, -7.306244, -5.827072, -5.492966, -4.038544, -4.358337, 
    -4.848175, -6.122131, -7.332809, -6.982819, -8.442444, -8.626053, 
    -9.490891, -9.265366, -9.816925, -8.429428, -10.744, -12.02423, 
    -13.76666, -14.6776, -13.97343, -11.94974, -14.64166, -13.10208, 
    -11.86406, -6.695572, -6.193497, -5.780212, -6.060669, -5.345581, 
    -4.974747, -6.464584, -9.475266, -13.64818, -17.81017, -18.8716, 
    -17.41798, -15.92758, -16.18674, -14.50574,
  -11.53932, -8.193756, -7.73204, -8.863007, -11.61563, -12.23489, -12.65494, 
    -11.60547, -10.43854, -7.047394, -8.422638, -15.37943, -21.28931, 
    -20.91092, -15.69089, -12.4039, -13.50833, -15.01874, -18.11511, 
    -19.46014, -14.36069, -9.813263, -10.48697, -13.49374, -14.20963, 
    -15.33466, -12.96509, -12.85809, -14.5643, -14.32294, -15.40469, 
    -15.61118, -16.52214, -15.18648, -13.57892, -8.478638, -7.742706, 
    -6.492432, -7.270325, -7.462769, -7.128372, -10.19868, -11.88672, 
    -9.376297, -7.777344, -3.201309, -0.1617126, -0.5041656, -2.608078, 
    -2.467453, 1.161987, 3.317184, 4.232544, 4.643234, 3.167709, 0.4453125, 
    -1.433334, -4.21666, -6.311722, -4.724991, -2.067703, -4.214325, 
    -10.62395, -15.44244, -16.80495, -16.50522, -20.01381, -26.44193, 
    -24.57005, -28.36121, -28.89244, -33.71484, -37.63335, -36.85989, 
    -37.13698, -38.46301, -35.08879, -28.27579, -29.53334, -25.39166, 
    -15.20157, -11.95808, -10.60469, -11.68752, -12.94348, -15.33308, 
    -17.52005, -17.20651, -15.30002, -13.2724, -12.99167, -10.98517, 
    -11.90623, -13.96146, -16.30991, -15.64714,
  -12.88931, -10.58618, -9.897156, -12.82318, -16.30051, -16.85599, 
    -14.13176, -13.1815, -11.22003, -12.67474, -17.8862, -28.44402, 
    -33.31795, -31.0453, -29.08827, -25.92943, -29.53358, -37.38724, 
    -34.7065, -26.13542, -21.55547, -18.14789, -17.20235, -16.70236, 
    -13.96094, -11.54425, -9.882294, -8.04245, -5.908325, -6.980988, 
    -7.324738, -14.50313, -14.57344, -11.56589, -14.65494, -23.37187, 
    -31.4427, -32.75859, -31.35234, -30.30078, -19.36589, -17.49792, 
    -14.99922, -12.25235, -6.354675, -3.932037, -3.424469, -3.241409, 
    -2.614594, -6.372391, -8.877869, -8.374741, -5.29921, -2.670822, -4.4039, 
    -1.247391, -0.004425049, -0.5585938, -2.640106, -3.8125, -4.940094, 
    -5.902603, -10.19559, -12.45313, -14.04869, -15.53725, -19.07655, 
    -21.91277, -18.38124, -13.42526, -11.65858, -14.15314, -16.05156, 
    -14.29608, -13.84688, -16.16197, -19.46198, -16.42865, -12.075, 
    -11.18256, -14.78151, -20.83464, -23.15443, -29.67682, -34.61691, 
    -34.84193, -28.34947, -22.94896, -20.0435, -22.06561, -20.35364, 
    -19.12317, -17.25964, -14.89764, -17.4086, -17.18802,
  -40.33125, -38.49062, -31.69765, -29.43019, -34.55312, -32.8591, -31.28307, 
    -34.73463, -31.88229, -32.56979, -28.57318, -21.12291, -21.53723, 
    -24.75546, -29.69531, -30.19193, -30.98412, -31.91667, -29.58984, 
    -35.76485, -41.78542, -41.35963, -33.90704, -34.32109, -33.66197, 
    -29.71355, -23.23776, -17.76772, -11.79375, -5.942444, -6.2612, 
    -10.47162, -9.334641, -6.092453, -8.59375, -11.40495, -10.92291, 
    -14.76901, -15.29453, -10.3362, -10.44818, -10.89427, -8.159119, 
    -5.378906, -6.238281, -7.229431, -9.521347, -9.768494, -9.191925, 
    -6.644791, -6.316666, -8.62735, -9.232285, -10.34975, -11.17787, 
    -13.14818, -14.16016, -11.63541, -9.878372, -6.092453, -9.210159, 
    -8.996872, -7.342438, -9.404175, -14.01666, -13.59193, -8.614319, 
    -4.862762, -7.560425, -5.717712, -2.996887, -7.119278, -7.351563, 
    -6.975006, -5.334641, -8.738022, -10.55678, -9.309891, -7.218216, 
    -8.042709, -11.62057, -7.953903, -3.682556, -6.411194, -11.71953, 
    -12.07448, -13.57109, -23.14375, -34.06302, -39.36226, -40.30858, 
    -44.45546, -42.29115, -39.71353, -39.92058, -39.50861,
  -7.984375, -4.270844, -4.21666, -5.041138, -4.844788, -8.304947, -9.116928, 
    -6.021088, -0.7507782, -1.224472, -5.341415, -7.215103, -11.01067, 
    -6.110947, -1.375519, -1.203903, -3.2099, -3.042175, -4.134644, 
    -9.691406, -7.335419, -2.230469, -0.3809967, -3.685669, -6.6539, 
    -4.814331, -3.951828, -5.996872, -11.60391, -9.185425, -6.758331, 
    -4.584366, -1.684113, -0.4307251, -0.4739532, 0.458847, 1.567978, 
    -3.829941, -6.791931, -3.964844, -4.379166, -3.450256, -0.1690216, 
    1.383331, -3.553116, -4.345825, -3.336716, -3.275787, -1.709122, 
    -3.525787, -2.272141, -2.636459, -2.246613, -0.2434998, -2.125793, 
    -3.997131, -6.427078, -5.089066, -4.919785, -6.296875, -4.449219, 
    -6.275253, -7.672409, -8.033585, -10.2901, -14.85573, -13.52448, 
    -8.602341, -12.19739, -9.605988, -5.243484, -3.690109, -1.433075, 
    -0.686203, -0.02708435, -1.649734, -0.2502594, -1.173965, 1.128113, 
    7.272919, 3.945572, -0.6971436, -8.382553, -10.5177, -13.07996, 
    -9.114075, -4.35495, -6.1539, -4.600266, -1.470825, -2.648956, -7.127075, 
    -7.906769, -8.561707, -11.4948, -9.769272,
  -4.257553, -5.127609, -7.745056, -4.996094, -7.823181, -9.728134, 
    -5.149231, -0.6526031, -2.650513, -0.6885376, 1.339844, 4.726303, 
    7.756241, 8.469269, 3.544022, 5.391663, 6.5, 4.867447, 0.4953156, 
    3.41095, 4.037506, 2.380981, -2.7677, 0.4312439, 2.998962, 2.704178, 
    1.113007, -7.006775, -11.55052, -6.092712, -1.395309, 3.193756, 2.590363, 
    -0.5609283, -2.222137, -4.997131, -3.002594, -0.4533844, -1.351044, 
    1.281769, 2.128128, 1.561722, 2.253647, 4.849472, 2.786469, 0.6648407, 
    3.770569, -2.395844, -0.3887939, -0.1166687, 3.722931, 7.328384, 
    6.523956, 3.829941, 3.850784, -0.3526001, 0.8411407, -4.186462, -7.58255, 
    -7.507278, -3.220566, -2.8302, -5.755203, -3.726044, 2.349747, -6.140625, 
    -2.562759, 0.0625, -3.139847, -0.9536438, -0.1947937, -3.802856, 
    -1.338013, 3.537766, 3.126297, 0.5690155, -0.09165955, 4.885147, 
    10.96693, 9.14035, 2.4646, 4.163269, 3.328125, -2.871094, -6.062241, 
    -6.280212, -5.25235, -3.088791, 2.178391, 1.92395, -2.849472, -7.883591, 
    -7.643234, -2.250534, -4.976822, -8.480728,
  -8.05806, -4.008072, -0.07917786, 0.3244934, -5.399994, -3.116409, 
    6.480469, 7.054947, 4.637512, 3.433594, 3.461197, 6.735428, 2.295319, 
    -1.769531, 3.069794, 0.8843842, 2.326813, 6.230728, -0.2541656, 
    -1.203125, 2.273438, 3.025513, 0.407547, -0.2205811, -1.350266, 
    -3.365097, -0.8726501, -0.2703094, 1.293228, 0.008865356, -1.686447, 
    2.158066, 3.972916, 5.409378, 1.851547, -2.331238, -0.4039307, 3.583603, 
    7.284134, 8.664063, 8.913788, 9.630478, 7.749741, 5.767456, 8.268738, 
    14.4888, 6.747665, 4.141144, 6.922668, 9.853119, 4.445831, 5.193741, 
    5.488022, 3.794266, 4.728394, 8.263275, 3.307297, 0.7002563, 3.71875, 
    5.757294, 3.59584, 5.629425, -0.2494812, -0.7726593, 7.659897, 7.877853, 
    11.23672, 12.96249, -0.8111877, -5.889572, -2.241928, -1.185425, 
    1.360428, 0.04374695, 1.755203, 2.942184, 12.54845, 17.05234, 12.72734, 
    5.464325, 1.008606, 0.8692627, 4.624481, -0.1447754, -5.450775, 
    0.8612061, -1.419266, -1.544266, 2.583603, 0.8125, 2.249466, -0.2111969, 
    -4.724991, -0.8195343, -0.7065125, -3.829681,
  5.065369, 1.924988, -0.7916718, 2.047913, 4.8349, 12.70807, 7.256256, 
    3.407806, 6.401031, 5.617188, 3.325256, 6.059387, 0.2106628, -6.067719, 
    -0.5278625, -1.546875, -0.1367188, -0.01223755, 0.5549316, 0.6143188, 
    4.616135, 3.331757, 6.515091, 6.155991, 6.346878, 11.71173, 8.15155, 
    9.806488, 13.44376, 12.85754, 5.029419, 5.028107, 1.381256, 6.395844, 
    6.132538, 8.289337, 7.411224, 2.454193, 9.644257, 15.28229, 8.563019, 
    6.216675, 11.22656, 9.218475, 9.0401, 10.89401, 14.03203, 7.982544, 
    4.191406, 1.504944, 3.081512, 4.481262, 7.780212, 8.617706, 9.698181, 
    7.48645, 7.491669, 7.506241, 4.425537, 2.104156, -2.284637, 2.735168, 
    3.175507, 3.894012, 7.041412, 7.48645, 5.513535, 8.370331, 1.091675, 
    0.8101501, 1.217957, 4.102356, 5.834381, 5.215118, 7.545837, 10.43671, 
    16.63986, 22.5974, 16.30495, 8.305481, 0.4557495, -4.737488, -5.306519, 
    0.3677063, 2.073944, 3.812744, -1.831238, 3.510651, 5.875519, 1.447662, 
    3.117188, 1.213806, 0.328125, 6.799469, 6.763275, 2.944275,
  2.606262, -1.277344, -0.5549622, 3.574493, 2.931763, -0.0609436, 
    -0.5635376, 3.107025, -2.224731, -2.926025, 0.2789001, 7.198181, 
    6.083862, 8.082275, 3.818481, 5.692719, 3.351288, 1.350525, 5.155212, 
    6.936218, 6.630463, 6.645325, 5.865631, 3.479706, 2.312775, 6.824219, 
    8.129425, 6.829407, 5.7547, -1.443512, 3.577606, 5.046082, -1.315613, 
    2.957031, 3.892181, -1.173431, 2.800507, 0.5143433, 13.63828, 23.00287, 
    11.01068, 3.29715, 5.333069, 6.804688, 3.979675, 3.401062, 12.14218, 
    19.90417, 5.463531, 7.7052, 11.37527, 10.16147, 11.59451, 13.21509, 
    9.276306, 11.83984, 11.22656, 7.21225, 7.822144, 6.814331, 8.45755, 
    4.6604, 6.788544, 6.6604, 7.082306, 2.708099, 2.057281, 3.074493, 
    5.160156, 6.332825, 4.077606, 6.534882, 11.40469, 9.3284, 8.102356, 
    8.1604, 20.56589, 39.70496, 7.917175, -6.367432, -2.190094, -6.227875, 
    -5.494537, -4.114838, -7.710419, -5.192688, -8.046356, -2.481506, 
    -5.523438, -5.001801, -3.6315, -2.747131, -5.153625, 1.490356, 3.939331, 
    0.2122192,
  -7.130981, -7.625275, -0.08126831, -6.240356, -3.145569, -1.391937, 
    -7.0289, -7.157013, -7.638275, -8.162231, 7.27475, 6.072113, 7.071869, 
    10.68387, -2.366669, -1.308838, 4.588257, -1.734375, 0.4020996, 
    0.8815002, 1.996613, 1.673981, -6.54895, -2.339844, -6.502319, 
    -0.8374939, 3.746613, 2.8815, 0.7093506, -3.016937, 4.297119, 3.528107, 
    -3.342712, -3.32135, -2.327362, -0.5833435, 2.452087, 1.182281, 6.805481, 
    5.565887, -8.746094, -8.721375, -2.470062, -3.684113, 1.458313, 
    0.3432312, 0.4620056, -0.8716125, 1.713531, 8.515869, 15.25235, 5.509369, 
    3.961731, 6.513794, 8.6987, 8.493469, 5.285675, 2.327057, 2.522644, 
    4.754181, 5.030487, 2.7388, 5.238556, 7.770813, 8.988007, 6.423706, 
    -0.8726501, 2.463776, 0.3796692, -1.922668, 2.04895, 5.093231, 4.808594, 
    4.342163, 2.471863, 1.476563, 10.51978, 13.41278, -3.131256, -21.63879, 
    -14.41483, -8.941681, -18.45547, -21.66537, -21.52005, -16.86224, 
    -11.60703, -8.772919, -8.424225, -5.46405, -2.107819, -3.921875, 
    -3.059631, -1.14505, -2.449219, -4.63855,
  -8.033081, -5.0961, -3.0625, -2.79895, 1.356262, 2.415375, -1.783356, 
    -12.88019, -14.4151, -12.87607, -6.005981, -5.748169, -4.311462, 
    -4.651825, -3.905731, -3.5625, 0.1640625, 0.4299622, 2.703369, 1.479431, 
    -5.69455, -5.713287, -3.003906, -5.298706, -6.594269, -7.055206, 
    -10.43436, -9.056763, -4.928131, 0.3510437, 3.391663, 2.361969, 
    -3.190369, -6.494537, -1.565094, -0.3893127, -1.619263, -1.797394, 
    -2.636719, -3.868225, -5.310944, -4.489594, -8.061981, -7.244781, 
    -5.568237, -5.005463, -6.074219, -2.407806, 4.7388, 3.416656, 3.525787, 
    6.076538, 4.346619, 6.399475, 4.10025, 1.581512, 0.2346497, -1.070313, 
    -3.052368, -0.005187988, 3.079681, 4.25885, 4.656799, 1.180481, 3.655182, 
    0.0718689, -3.140381, -5.698944, -4.091919, 1.220306, 2.967712, 
    -1.391693, -1.864868, 0.9398499, -0.2718811, -7.365631, -3.263275, 
    -7.372406, -10.02762, -22.34399, -32.17265, -19.66486, -26.39218, 
    -17.02316, -16.54245, -12.43542, -9.031494, -12.22086, -7.247681, 
    -3.377075, -10.97528, -8.745056, -9.461212, -9.976563, -8.966675, 
    -4.887268,
  -3.349487, -3.651031, -3.697937, -9.797394, -1.767975, -4.126038, 
    -5.911438, -9.073944, -8.248962, -5.458313, -7.278412, -0.07318115, 
    -6.106781, -8.8013, -0.3997498, 8.374725, 2.168213, 0.9940186, -2.929169, 
    -4.040344, 0.263031, -5.444519, -4.480194, -7.192169, -12.21616, 
    -10.77707, -6.490082, -5.702606, -0.2010498, 0.3661499, -1.155731, 
    -3.990875, -2.054169, -2.380219, -4.632813, -11.72501, -9.148712, 
    -7.606781, -4.658356, -0.6208496, 3.711975, -2.369019, -7.909393, 
    -0.9091187, -6.7836, -5.917969, -6.052368, -6.996368, -6.2052, -5.84375, 
    -2.337738, 2.863281, 5.049744, 5.601563, 4.088043, -2.07605, -3.121094, 
    -5.945862, -4.891144, -4.937775, 2.963531, 4.43335, -3.7966, -8.667694, 
    -10.71121, -6.838287, -7.803894, -11.83307, -7.8237, -2.85495, -5.7771, 
    -4.931488, 4.71405, 0.08358765, -4.710144, -2.428619, -7.624725, 
    -15.0802, -9.001282, -13.24634, -23.51564, -7.747925, -2.008072, 
    -2.978912, -4.544525, -11.21066, -2.27475, -11.06927, -8.420563, 
    -9.304169, -6.007294, -7.0495, -9.181244, -5.528381, -2.877594, 3.538544,
  -0.598938, -3.728912, -4.043243, -4.517456, -3.306519, -2.137482, 
    -7.066406, -1.865601, 1.615601, 3.079681, -3.069519, -4.357269, 
    -1.223175, 0.009094238, 3.547119, 6.352081, -1.464844, -1.682007, 
    1.196869, 3.264343, 4.8013, 1.341156, -3.810425, -6.223694, -4.348419, 
    -2.645569, -3.879944, -3.344513, 2.403381, 1.575256, -0.1833496, 
    -4.098969, -7.410156, -7.699738, -9.655182, -9.065887, -5.145569, 
    -6.366425, -5.806488, -2.42395, -1.745056, -3.261444, -1.026581, 
    -4.075775, -2.403656, -6.115631, -5.588806, -7.786469, -8.671631, 
    -1.014862, 2.401031, 1.322388, 2.979431, 8.1828, 5.2052, 3.0177, 
    -0.8760376, 1.721863, 0.7692871, -7.142975, -5.0466, -12.86148, 
    -16.19687, -20.84271, -19.22708, -14.99451, -13.23047, -11.73413, 
    -10.05676, -10.22656, -5.724243, 1.765625, -4.233856, -2.451294, 
    -2.912231, 0.1164246, -5.947144, -14.03619, -1.652344, 6.070297, 
    -8.597397, 9.489075, 1.956238, 4.656769, 2.176041, -4.103394, -6.659393, 
    -6.777863, -5.171356, -13.27527, -8.828888, -8.385162, -5.489594, 
    -2.278656, 2.758606, 0.9445496,
  -0.5411377, -1.027069, -13.26172, -5.382538, 0.09060669, 3.242462, 
    1.545044, -2.457031, 0.1960754, 5.020569, -1.825012, -8.6073, -5.542694, 
    11.21745, 2.5336, 3.225006, 1.437775, 3.657013, 5.212769, 2.280212, 
    5.676575, 1.574493, -2.289063, -10.86746, -2.107269, 2.773438, 3.188019, 
    6.013306, 5.555481, 0.2098999, -1.144287, -6.172394, -9.336975, 
    -5.673187, -3.582794, -7.704681, -10.37552, -7.895294, -1.805725, 
    -1.648956, -7.4198, -3.81485, -6.849213, -3.419281, -0.6507874, 
    -0.8406372, 4.019531, 1.214294, 0.278656, 12.06119, 6.2211, 7.8815, 
    7.53595, 3.866394, 6.284363, 3.035675, -2.183319, -3.468994, -7.157043, 
    -16.19922, -24.95831, -33.00313, -25.52658, -18.83307, -17.66144, 
    -18.66534, -14.56302, -8.200531, -3.606262, -0.01171875, 0.3927002, 
    7.103668, 2.122925, 6.125519, -1.904968, -9.796631, -6.815613, -10.21042, 
    11.1651, 16.83437, -2.4133, 9.152618, 2.388, 5.938538, 7.583847, 
    10.17996, 0.1182251, -3.456787, -4.535675, -4.734619, -4.665619, -1.2789, 
    1.086456, 1.489838, 3.563049, 6.258575,
  3.15625, -0.9078369, -3.387238, -4.215118, 7.40155, 6.886993, 4.564056, 
    -2.009644, -1.282532, 7.004944, 4.212769, -6.231232, 2.197403, 14.64037, 
    8.583618, 8.215881, 7.720581, 12.08594, 1.72995, -3.718994, -0.9908752, 
    0.05258179, -0.4403687, 1.186737, 0.6489868, 6.375244, 7.225281, 
    6.714844, 5.412476, 0.5804749, -0.7908936, -6.065613, -6.958588, 
    -8.966675, -6.879181, -7.450775, -6.489044, -5.562775, -4.256531, 
    -0.7794495, -2.832825, -1.861725, -3.740356, -0.9518127, 2.513, 2.183594, 
    5.39035, 6.617706, 12.1599, 14.20651, 7.820557, -1.732819, 0.6460876, 
    -2.610168, 0.5674438, -1.41275, -8.976563, -19.33749, -19.72684, 
    -16.03412, -17.98984, -15.45728, -11.27081, -12.22107, -10.20157, 
    -5.34845, -3.133575, -1.191925, 2.055725, 8.205719, 5.436707, 10.48645, 
    9.014069, 7.128632, -2.107025, -4.559906, -6.478638, -0.5750122, 
    26.02553, 12.98048, 1.686737, 14.71172, 5.630463, -3.3367, 2.622131, 
    19.75858, -6.141663, -5.072662, 1.00885, -0.2932434, -0.01928711, 
    1.712006, 1.130219, 4.386719, 3.418488, 4.925781,
  7.7565, 2.588287, 7.858612, 2.223419, 17.44087, 10.6198, 10.66823, 
    10.43463, 7.024719, 8.9758, 11.52524, 1.791931, 1.969513, 7.5401, 
    8.600525, 14.10989, 11.94662, 7.387756, -0.212738, 0.3299255, 0.7065125, 
    -1.779144, 2.737244, 1.355469, 2.185699, 3.077576, 6.054138, 2.433594, 
    2.131256, 0.7966309, -1.389038, -2.8125, -7.664307, -7.38385, -9.317963, 
    -5.665131, -6.152344, -5.005463, -3.246643, -1.114319, -7.079437, 
    -3.7612, -0.6598816, -0.3645935, 4.963531, 5.103363, 5.091919, 3.587234, 
    2.089844, -3.103638, -0.2286377, -6.586456, -13.27917, -8.989044, 
    -7.736694, -13.95468, -15.32056, -16.64063, -8.959381, -3.6203, 
    -4.611481, -2.929443, -8.302887, -5.719543, -3.533844, 0.2661438, 
    1.38855, 6.135147, 8.497131, 9.110672, 12.86952, 11.84427, 15.25287, 
    14.2883, -2.964844, -6.483337, -13.18256, -1.486191, 20.88803, 7.581268, 
    9.933334, 5.247406, -9.2966, -12.32578, -4.238281, 16.31824, -2.089081, 
    -6.534912, 3.998688, 1.118988, 4.166138, 5.457031, 6.135956, 10.27316, 
    7.147675, 8.32605,
  7.48175, 4.936218, 8.925232, 8.828674, 13.92317, 8.917709, 8.27005, 
    1.650772, 4.749222, 21.4987, 15.8065, 5.213287, 6.012482, 3.571106, 
    1.424988, 5.539063, 1.648178, -0.7338562, -3.768738, -2.974457, 
    0.2914124, 2.389832, -0.08856201, -1.345306, 2.265625, 2.453674, 
    -2.216644, -7.186462, -7.397644, -2.291412, -6.273438, -4.993744, 
    -5.710938, -5.928101, -3.538544, -4.642426, -2.174469, 1.117981, 
    0.8158875, 4.68045, 7.32785, 9.811462, 2.7901, -5.638794, -4.030457, 
    -6.452072, 2.837753, 9.146103, 2.274216, -4.754944, -0.6434937, 
    -6.827087, -13.99741, -12.48491, -13.01379, -9.831238, -8.907318, 
    -4.768768, -0.5776062, 0.6895752, 3.3909, -0.2846375, -1.608856, 
    -0.8273315, 0.265625, 7.694794, 8.782547, 13.44922, 14.08775, 16.20546, 
    17.14192, 13.38098, 17.79819, 10.82397, -7.315887, -15.99583, 1.510155, 
    18.25287, 6.170837, 10.55989, -0.3648376, -11.20103, -10.40001, 
    -7.001816, 1.333069, 2.082825, 12.23669, -0.8533936, -2.624481, 
    -0.3388062, 4.344269, 5.296356, 4.152084, 10.33984, 8.507568, 10.44089,
  11.55936, 9.945068, 9.310669, 4.744537, 8.813278, 3.201569, 0.481781, 
    -5.905731, -6.947128, 5.629166, 5.801559, 3.060394, 5.035431, 0.2825317, 
    -7.157547, -2.82135, 0.2296753, 0.1984406, -0.7604218, -3.767975, 
    -5.556763, -0.8288879, -4.325531, 3.016663, 4.319763, 1.060944, 
    0.7158813, -9.752869, -10.69427, -0.1648254, -1.114075, -1.038025, 
    -3.421356, -3.037506, -2.736206, 0.9567871, 8.354431, 23.05052, 3.478127, 
    1.891144, -0.1971436, 8.738281, 4.874481, -5.335159, -9.773178, 
    -13.45964, -9.551041, -9.125793, -14.13228, -17.09425, -19.54295, 
    -14.28517, -17.55495, -21.73933, -20.87003, -17.58099, -12.50522, 
    -9.317444, -3.530487, -3.562225, 1.571106, 2.309387, 5.574219, 8.134125, 
    10.5289, 12.00937, 13.04114, 13.4982, 17.81302, 15.33023, 13.34662, 
    11.92734, 5.393494, -2.443237, -3.773697, 5.728119, 11.25548, 1.420303, 
    16.76277, 5.745834, 2.681, 12.29713, 15.33151, 4.706512, -0.1513062, 
    -8.144531, 2.8927, 4.348175, 0.8356934, -0.3851624, -0.1953125, 3.820068, 
    5.117462, 8.410675, 9.908325, 9.750275,
  -1.850525, 2.058868, 4.884369, 2.225525, 10.22083, 6.215363, 7.915359, 
    11.35234, -3, -13.51459, -11.93517, -0.1471405, -0.8981628, -2.688797, 
    -8.137238, -1.686722, 5.482025, 10.12579, 3.435684, -0.890625, -6.354431, 
    -4.600021, 1.508072, 0.1109467, -0.8132935, -9.502884, -6.123703, 
    -1.911972, -22.31093, -11.77264, -6.953125, -10.09506, -9.541412, 
    -5.465637, -7.052612, -1.451035, 0.7375031, -2.727081, -10.14401, 
    -15.64558, -8.125778, -5.454163, -4.193237, -7.752869, -13.55312, 
    -19.8461, -23.95911, -27.18256, -27.73856, -22.55861, -18.72397, 
    -17.88101, -14.91666, -12.16769, -9.573425, -9.594543, -5.430481, 
    -5.100525, -3.876038, -3.705475, -0.7864685, -2.219788, -0.7765503, 
    0.5617065, 0.1369629, 4.751068, 3.329681, 0.1315308, -1.193207, 
    -3.496613, -6.848724, -6.909607, -16.20261, -9.153641, -5.680206, 
    8.692703, 18.38568, 7.549225, 18.93593, 8.258072, 25.42682, 15.84322, 
    2.809875, 0.07293701, 4.438538, 1.734619, 4.508606, 4.294769, 0.6895752, 
    0.05783081, -0.359375, -0.2851563, -0.0249939, 0.4156189, -0.4172058, 
    -2.097656,
  2.655472, 0.07421875, 7.686462, 12.38515, 16.71666, 10.16641, 3.246353, 
    -8.978897, -21.18594, -30.59557, -26.57213, -11.46016, -5.041931, -6.75, 
    -12.25156, -13.42447, -4.227615, -1.066681, 0.1112061, -1.614319, 
    -2.871353, -6.144531, 3.219528, 1.638809, 5.694534, -9.465622, -26.625, 
    -8.396095, -22.04713, -18.00755, -18.27396, -4.961456, -0.01641083, 
    -7.807556, -8.777863, -3.7836, 2.137253, -1.884903, -9.435928, -10.03645, 
    -11.49687, -10.56276, -11.43906, -13.26563, -16.5625, -18.87656, 
    -28.42813, -33.26822, -34.35858, -29.02007, -31.98776, -25.20703, 
    -22.47658, -20.87866, -18.05573, -16.65573, -12.74768, -8.940887, 
    -9.407043, -9.210938, -10.08359, -8.526276, -10.47214, -9.764832, 
    -6.31955, -5.142181, -2.75235, -2.045837, -2.87735, -4.083069, -7.623947, 
    -3.559647, -18.51407, -22.51848, -20.74922, 1.058594, 43.88203, 8.055206, 
    6.355209, 35.05754, 14.69453, 3.792206, 1.905472, -1.041412, 0.263031, 
    7.106247, 4.516663, 3.239075, 0.9450684, 2.999481, 1.283325, -2.180969, 
    1.397644, 1.622406, 1.717712, 2.798706,
  2.831512, -4.076035, 8.2034, 13.6888, 0.4755249, -4.623184, -14.57187, 
    -21.98567, -20.70442, -17.28984, -21.64088, -22.35493, -15.00729, 
    -12.78723, -8.961975, -15.08646, -12.4664, -9.750778, -10.76146, 
    -9.765106, -6.967712, -4.362503, 4.870575, 7.827606, 4.463013, 0.3205719, 
    -1.125275, 6.357819, -9.579437, 0.8697815, -0.03515625, -1.800262, 
    -2.20079, -0.3117218, -0.9903564, 0.9950562, 3.449997, 0.4695435, 
    -3.108856, -7.371094, -12.07579, -11.95338, -9.835938, -9.115616, 
    -12.20338, -7.909363, -4.560928, -5.414841, -4.914322, -3.554947, 
    -10.90416, -10.28151, -16.04271, -17.35443, -17.1526, -16.77605, 
    -11.4435, -6.158844, -4.9263, -3.964066, -4.102341, -3.444534, -1.702606, 
    0.07603455, 4.996613, 8.700256, 8.585159, 7.907547, 2.664581, -3.472137, 
    0.5442657, -0.7986908, -3.638031, -1.694534, 3.094788, 16.59635, 
    31.24844, 11.63802, 18.17813, 28.33281, 1.944275, -1.176041, 3.210419, 
    3.745834, 7.375, 8.582291, 9.068756, 8.707031, 6.384628, 5.172394, 
    2.9646, -1.440643, -0.354187, -2.2836, 5.058853, 1.983078,
  -7.282547, -9.767456, -6.476059, -5.614319, -4.806, -3.565369, -8.049744, 
    -11.35208, -9.783081, -17.95964, -32.06978, -17.95313, -16.17136, 
    -12.30026, 1.640106, -4.245575, -8.579941, -5.219009, -3.001053, 
    -7.427856, -5.587769, -2.740112, 7.610428, 7.466141, 3.021881, 
    -0.4124908, -5.154434, 0.504425, 0.467453, 9.096603, 9.830994, 5.363541, 
    -3.467957, 0.3721466, 8.45079, 6.386719, 5.441147, -5.947922, -5.233322, 
    -5.395309, -6.276031, -5.640884, -9.254425, -9.037491, -10.57968, 
    -1.567719, 0.5622406, 3.489594, 7.788284, 8.737762, 8.259369, 8.746353, 
    10.90755, 14.27995, 19.58673, 20.85989, 18.92084, 16.54375, 14.6091, 
    12.90468, 2.905212, 1.234634, 1.567444, 4.147659, 6.380981, 6.714584, 
    5.12265, 0.4320374, -0.8223877, 2.230728, 7.595047, 0.8364716, 3.921616, 
    10.96225, 27.14792, 22.51485, 28.62968, 22.58203, 10.30626, 11.89401, 
    2.404953, 4.312241, 2.103897, 6.864838, 12.00157, 5.636459, 4.790115, 
    1.251038, 1.078918, -1.240875, -4.775253, -6.505203, -4.509369, 
    -7.334381, -6.378387, -6.5625,
  -8.04245, -11.09557, -9.88855, -8.998169, -8.597397, -6.002075, -7.386185, 
    -8.173187, -8.014313, -11.83098, -15.05156, -12.0435, -18.93176, 
    -10.63802, 0.2770844, -0.3020782, 0.8440094, -0.1229095, -3.670837, 
    -7.935944, -6.268738, 5.004425, 4.621353, 6.537506, 8.810165, 6.355209, 
    -2.128906, -1.697144, 10.05286, 4.190353, 1.980209, 8.931, 1.1698, 
    7.453125, 5.347397, 2.263794, 0.5848999, -3.299484, -5.269272, -2.0289, 
    -1.264328, 0.046875, -0.4398499, -0.686203, -1.205994, 0.9427185, 
    -1.577606, -0.4489594, -0.1578217, 5.777344, 5.928909, 9.429428, 
    3.314072, 8.632294, 10.97136, 11.63568, 12.14531, 12.25417, 8.408325, 
    3.701309, 1.257019, 0.0236969, 0.4054718, 3.777603, 6.663025, 0.1596375, 
    -2.726303, -3.105209, -6.212234, -6.451035, -5.536987, -6.648697, 
    7.984116, 25.92422, 10.83438, 3.466415, 1.480209, 4.528122, 2.064575, 
    3.514313, 3.263535, 1.027863, 1.911469, 4.036728, 1.065369, 4.032288, 
    2.772659, 1.693237, -0.2984467, 2.241394, -2.791672, -1.995316, 
    -4.760162, -6.592194, -6.843491, -7.1138,
  -6.729431, -8.072403, -10.42395, -9.527344, -7.733582, -7.085678, 
    -5.371094, -6.701035, -7.146088, -6.019531, -6.940887, -12.51094, 
    -14.31641, -13.26457, -8.330734, 1.546082, 4.641678, 2.509125, 0.9750061, 
    -7.185669, -12.66953, 4.882034, -1.224213, -1.805725, 9.665894, 2.848694, 
    -0.359375, -5.478378, 1.257294, -0.9921875, 0.4385529, -0.1083221, 
    6.249741, 5.987762, 2.220566, 7.226044, -0.2906189, 0.3731842, 2.674225, 
    7.695053, 4.762756, 3.244797, 3.373688, 6.235931, 4.146088, 5.825775, 
    7.24791, 5.632813, 5.994797, 7.795837, 8.691406, 4.725266, 7.06459, 
    5.558853, 7.789063, 2.577866, -1.106506, -3.953644, -3.50885, -1.820313, 
    -2.80365, -3.457291, -0.5513, 3.003906, -2.313797, -3.344269, -6.316406, 
    -8.04921, -11.06615, -4.950531, -1.645828, 11.10234, 25.7849, 12.84036, 
    2.439056, 5.611984, 9.135941, 8.757294, 9.264069, 9.061188, 8.223709, 
    9.516922, 1.886719, -3.315613, -1.918228, 4.949219, -1.052338, 9.155457, 
    6.495834, 6.009903, 0.1898499, -3.168747, -4.631256, -4.649994, 
    -6.076309, -6.347916,
  -4.329178, -3.983063, -4.692184, -6.787506, -6.858337, -6.928116, 
    -5.181519, -4.105988, -4.849472, -5.075256, -6.354431, -9.108078, 
    -8.114853, -6.99791, -9.346085, -0.4648438, -1.308868, -3.809891, 
    -5.711197, -4.639587, -9.269531, -10.87189, -2.556503, 2.489075, 
    7.515625, 9.445831, 2.286972, 0.2484436, -2.654678, -1.66954, -2.068497, 
    -2.414841, 2.221878, 5.304428, -0.6062469, 6.213806, -0.5716095, 
    -0.8929596, -0.4263, 1.465897, -0.5223999, 0.1231689, -0.1927032, 
    3.624741, 2.515625, 4.261978, 2.975784, 3.365891, 5.780212, 5.495575, 
    3.622391, 3.759628, 5.589066, 5.985947, 2.443497, -1.538284, -2.846863, 
    -5.701294, -6.229675, -7.162491, -3.604431, -0.3039093, 1.540359, 
    2.092194, 2.042969, -0.8729248, -6.203384, -8.624741, -5.318497, -1.8526, 
    9.756508, 18.37656, 18.84608, 4.271088, 4.849487, 5.951828, 5.512497, 
    10.41719, 10.20052, 5.530731, 5.475784, 3.454422, 3.695313, 3.383591, 
    -2.905991, -3.759644, -3.275528, 3.003372, 3.191132, 9.529434, 2.444794, 
    -2.322647, -3.600266, -4.740891, -3.877869, -4.855728,
  -1.629684, -0.9260406, 0.2661438, -2.358063, -3.776031, -3.676041, 
    -3.792191, -4.488022, -3.355728, -3.936722, -5.075256, -8.263794, 
    -8.529419, -5.397659, -3.287247, -2.807556, -1.930481, -5.034897, 
    -5.595566, -6.032288, -8.592712, -10.33438, -6.686966, -3.834381, 
    0.8427124, 5.527344, 3.652084, -6.138016, 2.199997, -0.06770325, 
    -0.05781555, -4.423172, -4.711716, 1.57058, 0.380722, 1.618225, 3.11145, 
    -1.54895, -0.4736938, 1.303116, 0.296875, 3.59166, 2.897385, 1.398956, 
    2.227356, 3.416672, 1.015366, 2.080475, 3.670303, 5.311462, 6.944016, 
    7.243484, 3.1362, 1.615891, 3.152603, -0.1145782, -0.8156281, -4.554688, 
    -2.063278, -0.9411469, 0.978653, 2.697647, 0.4156342, 1.502609, 
    -0.9338531, 0.5463562, -2.323441, -4.2547, -4.697922, 1.218231, 2.17421, 
    5.644531, 6.183594, 2.713547, 2.668228, -0.2791748, -0.28125, 2.398438, 
    4.787766, 3.003372, -0.2260284, 0.4645844, 3.771866, 0.9968872, 
    -0.5843658, 4.384125, 1.972916, -4.344009, 2.277603, 4.598434, 4.613281, 
    2.38385, -2.851563, -1.538025, -1.365356, -1.169006,
  0.4598999, 0.6546936, 2.416931, -1.677597, -1.44635, -3.552872, -3.597916, 
    -3.674744, -0.776825, -0.5351563, -4.282028, -7.521347, -13.19531, 
    -8.782303, -3.260941, -6.557541, -5.378647, -4.96875, -7.958588, 
    -5.470825, -4.824478, -5.178391, -6.286987, -5.593491, -10.92891, 
    0.1015625, -1.880203, -8.113281, -0.3986969, 9.172661, 7.97995, 3.155724, 
    0.5567703, 0.04401398, 3.162766, -0.5955658, 0.2416687, -1.651566, 
    0.4791718, -1.724747, -1.956238, 1.036453, 1.880737, 1.551041, 1.86145, 
    0.6408844, -0.478653, 0.5690155, -0.5749969, 0.3742218, 3.159637, 
    3.364578, 0.7476654, 4.77916, -0.0255127, -1.96875, -3.063812, -5.811981, 
    -3.099213, -5.688812, -1.984634, 1.90834, 6.512238, 1.640884, -1.423691, 
    1.770569, 4.0224, 3.604691, 3.214066, -4.745834, -0.5111847, 1.117966, 
    -3.066406, -3.664322, -0.7156219, 1.595047, 4.61615, 1.166656, 1.00235, 
    0.5390625, 0.8062439, -2.380722, -0.2848969, 1.295059, 1.160934, 
    1.732819, -0.7270813, 0.4997406, 0.5880127, -1.498962, 2.125, 3.617188, 
    6.718491, 5.595047, 2.135422, 1.005997,
  8.474472, 4.164322, 2.932037, -0.5031128, -0.4968719, -1.014847, 2.703125, 
    0.1338501, -1.507813, 6.206772, 1.695831, -3.065887, -6.241135, 
    -6.197662, -8.226044, -9.195313, -8.418243, -5.434387, -1.512497, 
    -3.317978, -2.439316, -2.674728, -11.09921, -7.794006, -7.110413, 
    -7.812759, -10.63359, -14.60652, -3.804947, 9.248955, 6.16433, 5.030205, 
    3.617714, 0.1906281, 3.757294, 2.131248, 3.844009, -0.08879852, 
    -1.306252, 0.8825531, 0.0700531, 1.989578, 3.246353, 2.697655, 3.490364, 
    -1.851563, -0.816925, -1.418228, 1.231255, 2.732025, 3.897133, -2.298172, 
    0.0007858276, -0.4507751, -3.871353, -2.18515, 0.3554688, 1.18203, 
    -1.338806, 3.276047, 0.816925, 0.9335938, 5.057037, 6.514587, -0.3135376, 
    0.7341156, 4.496613, 8.345322, 6.490891, 0.6875, -1.663544, -2.419006, 
    -2.561195, -4.8862, -1.338547, -0.9945221, 0.2440109, 1.536201, -1.2099, 
    0.7020798, 1.298958, 0.8091125, -0.221611, 4.236977, 2.949745, 1.166153, 
    2.655991, 4.25338, 1.695831, 1.31823, 4.488274, 1.229691, 10.44141, 
    12.931, 18.42813, 20.9323,
  17.019, 18.73985, 10.31328, 4.865105, 4.770576, 3.09948, 6.778389, 
    7.310165, 9.029945, 13.86015, 9.12291, 5.060684, -0.9281158, 1.421616, 
    -1.24662, -4.03672, -2.259109, -2.191406, -3.681244, -6.534645, 
    -6.354416, -6.782547, -5.253128, -6.961716, -9.973175, -8.923172, 
    -8.559631, -11.21015, -3.432816, 0.5041656, 2.225266, 3.044792, 2.927345, 
    2.704422, 3.964577, 3.633858, 0.8562469, 2.27005, -0.1346359, 1.626816, 
    1.820053, 1.302864, 4.504166, 1.88073, 1.822914, -1.821617, 1.233856, 
    -0.2242203, -4.498955, -0.734642, 1.914848, 1.868752, -0.9554672, 
    -1.391403, -2.549736, -0.4770813, 0.1755142, 2.887238, 2.415108, 
    -0.04557037, 1.942451, 2.380989, 2.703392, 3.398697, 2.60807, 1.595322, 
    2.29583, 5.20417, 4.921089, -0.2919159, 2.435417, 0.6291656, -5.825264, 
    -3.046875, -3.275002, -1.318748, -0.579689, -1.428383, -0.3184891, 
    2.498695, 0.5679703, 1.571609, 3.935677, 2.261719, 1.417969, 4.542969, 
    2.500259, 1.459892, 2.249222, 2.324738, -0.08802032, -0.006507874, 
    4.340103, 8.955727, 15.83047, 20.02657,
  14.8862, 7.006775, 3.977089, 6.730469, 1.642189, 1.205467, 4.934898, 
    4.878647, 9.210678, 14.2888, 11.325, 10.18125, 4.669533, 2.327087, 
    2.343231, 1.855469, 0.6330719, 0.2020798, -0.3291626, -1.706253, 
    -1.291405, -3.302605, -4.028648, -5.9375, -6.542709, -8.573959, 
    -9.089844, -6.937759, -4.321617, -8.436722, -4.6362, -2.073959, 
    -4.098961, -6.705734, -5.31823, -2.711197, -0.8606796, -1.595833, 
    -1.603912, -0.1828079, 2.299744, -1.430992, -1.980988, 1.588799, 
    3.087494, -0.0627594, -2.093231, 0.8880234, 0.3736954, -2.055206, 
    -1.164589, -1.583595, -2.208336, -0.8265686, 0.2679672, -0.1351624, 
    -1.624733, 0.7361984, 0.7432327, -0.3197937, -0.705986, -2.879166, 
    0.3651047, 3.4039, 1.331245, -2.904427, -1.347397, -1.137505, -0.6705704, 
    -2.385155, -1.067451, 0.9640579, -1.716408, -2.458069, -1.518745, 
    -3.475258, -3.630989, -1.951569, -3.047134, 1.521355, 0.9752579, 
    2.675522, 4.339584, 0.3778687, 1.385162, 3.980209, 5.337761, 5.111977, 
    2.735939, 1.922394, 1.77578, 4.994537, 4.532028, 5.613022, 15.73177, 
    16.14219,
  2.414063, -0.008590698, 4.669533, 7.297134, 3.955215, 3.683594, -0.7580719, 
    -4.233074, 1.261978, 8.041145, 3.434113, 2.46328, 1.666145, -1.187241, 
    -1.697136, -3.670052, -5.913536, -5.828125, -1.032288, -1.835938, 
    -3.710419, -2.729172, -6.526558, -6.588799, -4.329689, -4.195839, 
    -5.214844, -4.718491, -5.86042, -8.323959, -6.899216, -5.93177, 
    -8.354431, -6.905991, -8.460678, -7.690887, -2.060936, 0.4325485, 
    0.4802094, 1.861198, 1.068748, -0.1273499, 0.8557358, -0.8026047, 
    1.113022, 0.4463501, -2.617447, -2.957558, 1.049217, 0.09140778, 
    -3.258331, 0.3742218, 1.552086, 0.7898483, 0.5697861, 1.167709, 
    0.5333328, -1.679947, -2.555992, -0.5854187, 1.164841, 2.941925, 
    0.455986, -0.6119766, -3.247917, -4.165886, -2.687756, -4.728645, 
    -4.846619, -5.902863, -5.725517, -4.808853, -2.88047, 0.001304626, 
    -0.9713593, -2.06094, -2.269276, -2.482292, -2.103653, -1.523438, 
    0.8234406, 0.7177124, -1.458595, 1.054955, 1.363281, -0.4835968, 
    -3.399734, 0.7541656, 0.901825, -2.107033, -0.1541672, 2.744011, 
    5.324997, 2.490364, 1.236458, 4.675522,
  0.1679688, -2.700001, -2.908852, -0.08463669, -4.019531, -2.560936, 
    -1.468227, -1.532028, -0.06041718, -0.4544258, -2.716408, -2.739582, 
    -1.842186, -3.507553, -3.626564, -3.608593, -5.416664, -7.452862, 
    -4.287762, -6.103905, -6.811718, -4.59375, -4.300781, -3.427086, 
    -1.461205, -0.1630249, -0.589325, -1.848694, -4.141663, -2.440102, 
    -1.428909, -4.334892, -5.948181, -5.523438, -7.221092, -8.15078, 
    -5.752861, -3.753906, -2.947136, 0.203907, -0.2799492, -2.482552, 
    0.1153641, -0.8976555, -0.8447914, 1.061459, -2.171875, -3.915623, 
    0.2411461, -0.1065102, -0.3085938, 1.078125, 1.846092, 0.7718735, 
    -0.4776039, 1.234375, 1.603382, -1.565102, -0.1945305, -0.2304688, 
    1.038021, 0.6966133, 2.291405, 1.087502, -0.7450485, -2.637241, 
    -2.683071, -5.346355, -4.636719, -5.916405, -7.504951, -4.972656, 
    -1.86224, -1.046352, -1.248695, -3.334377, -3.246613, -3.728905, 
    -3.287762, -2.010418, 0.8260422, -1.083855, -3.003906, -1.467705, 
    -0.4986992, -1.970051, 0.5039063, 0.4656258, -2.015625, -1.832813, 
    -1.751041, -0.3908844, 1.640625, 0.549221, -2.880207, -0.04531097,
  -0.8468761, -3.467188, -3.675522, -1.140884, -0.7718773, -2.229948, 
    -2.283855, -4.440365, -2.470312, -3.934637, -4.443748, -3.253643, 
    -3.641146, -5.066406, -4.745571, -3.015625, -4.687759, -5.978645, 
    -3.284374, -3.596615, -4.427864, -3.278645, -1.457291, -1.797134, 
    -0.7559891, -0.9223976, -0.5286446, -1.923439, -3.339844, -5.40469, 
    -4.119007, -5.84922, -5.477081, -4.885155, -4.010937, -4.739063, -5.1138, 
    -4.492451, -3.270836, 0.4924469, -0.685936, -3.271873, 0.3020859, 
    0.5838509, -0.7166672, -0.1184883, -0.8919258, -1.875782, 0.05703354, 
    -1.012501, -2.201824, -2.045834, -1.822914, -1.900261, -1.266148, 
    -0.6736984, 0.6408844, -0.3382835, 0.2645836, 0.9734383, 1.582813, 
    1.38932, 1.190104, -1.029167, -2.152082, -3.255989, -2.195576, -1.585938, 
    -2.570313, -3.319012, -3.044792, -2.497658, -0.1705704, -0.879425, 
    -0.7596359, -1.115883, -1.109896, 1.077347, 0.5533829, -0.2026024, 
    0.03619766, -0.5013008, -0.767189, 0.3968773, -2.224998, -1.448177, 
    1.691925, 1.176304, -1.751823, 0.04401016, -0.183075, -1.118229, 
    -1.035156, 0.9911461, -0.7276039, -0.5351563,
  1.816927, 0.1351566, -0.3851566, -1.412762, -2.340885, -1.512501, 
    -2.847136, -3.792187, -3.856771, -1.275782, -1.254686, -1.942709, 
    -1.539843, -1.285418, -1.430468, -2.337761, -2.488802, -1.330469, 
    -0.1833344, -1.707291, -3.435938, -1.735678, -1.340626, 0.4882813, 
    0.7624989, 0.1140614, -0.3768215, -1.138542, -1.870052, -3.863802, 
    -4.590103, -4.389585, -3.47422, -2.295574, -3.005989, -2.557552, 
    -2.785679, -2.814583, -1.068748, -0.1315098, -0.1695309, 0.2911453, 
    -0.07291603, 0.8786469, 0.7414055, 0.1427078, 0.2005215, -0.04374886, 
    0.2789059, -0.3416653, -1.335157, -0.9273434, -0.3828125, -0.5213547, 
    -0.6937485, 0.2015629, 1.907553, 2.389582, 0.922657, -0.2369804, -0.625, 
    -1.26927, -2.104427, -1.722395, -1.78698, -2.926043, -3.376041, 
    -3.291668, -2.748959, -2.371614, -1.212238, -0.6283855, -0.3591156, 
    -1.59453, -0.8367195, -0.5442696, -0.7489586, -1.746094, -1.783854, 
    -1.409115, -1.121353, 0.05416679, 2.11146, 1.201302, -0.7304688, 
    -0.4552078, 0.7640629, 0.8598957, 0.3335934, 0.7877598, 1.403126, 
    -1.039843, -1.108595, -0.4390621, 0.8875008, 2.284636,
  -1.827343, -0.5635414, 0.001301765, 0.620573, 0.4874992, -0.4471359, 
    -1.949219, -2.108854, -2.425261, -1.909375, -1.520312, -1.252865, 
    -1.064584, -0.75599, -0.7692709, -1.014323, -1.186978, -0.4260426, 
    -0.5023422, -1.419271, -0.8635426, -0.1914063, -0.6299486, -1.111198, 
    -1.194271, -1.050001, -1.814584, -2.329428, -2.453124, -2.240104, 
    -2.266928, -2.46302, -1.992449, -2.199219, -3.391145, -3.056252, 
    -2.390886, -0.2486992, 1.557032, 1.451042, 1.843229, 1.548697, 0.1687508, 
    -0.3773441, 0.370573, 0.7145844, 0.9789066, -0.5177097, -0.457552, 
    -0.7380219, -0.8877602, -0.5059891, -0.2614594, 0.2843761, 0.422657, 
    -0.4697914, -1.38698, -0.901041, 0.3091164, -0.1828117, -0.8127604, 
    -1.084896, -1.075521, -1.16875, -0.4846363, -1.541405, -3.323439, 
    -2.706511, -2.097135, -1.164844, -1.34974, -1.021614, 0.2036457, 
    0.764843, -0.5997391, -2.259113, -3.292448, -2.971875, -2.633855, 
    -1.287761, 0.1437511, 0.5533848, 0.2364578, -1.165886, -0.5028629, 
    0.05677032, 0.1046867, 0.07343864, -0.1434898, 0.5606766, 0.9921875, 
    0.7557297, -0.1151028, -1.167187, -1.54974, -1.119532,
  -1.330209, -1.376822, -0.7166667, -0.7263021, -0.7669272, -0.5299482, 
    -0.8895836, -1.295313, -0.973177, -0.7203126, -0.6713543, -0.7763023, 
    -0.8453126, -0.850781, -0.893229, -0.5585938, -0.4203129, -0.5130205, 
    -1.047656, -1.511459, -1.116926, -0.7049484, -1.14375, -1.929427, 
    -1.701562, -0.9924479, -0.4416666, -0.5752606, -1.144531, -1.042448, 
    -0.7848959, -0.6335936, -1.065364, -1.223699, -1.660156, -2.040105, 
    -1.895833, -1.280209, -0.4070311, 0.03932285, -0.4247398, -0.7041674, 
    -1.236458, -1.4375, -0.8895826, -0.5231771, 0.6895828, 1.476042, 
    1.002604, 0.4049482, 0.0354166, -0.6963539, -0.9893227, -1.152083, 
    -1.575781, -2.059896, -1.610938, -0.4919271, -0.488802, -0.6190104, 
    -0.9463539, -0.9085937, -1.010417, -1.058333, -0.9796877, -1.526563, 
    -1.923959, -1.744532, -1.150521, -0.9333329, -0.614584, -0.6312504, 
    -0.9507809, -1.057032, -1.982291, -2.228125, -1.904167, -1.647917, 
    -1.939062, -1.206771, 0.2223959, 0.214323, -0.119792, -0.30651, 
    -0.5770836, -0.8500004, -1.023958, -0.6807289, -0.1239586, 0.07656193, 
    0.270833, -0.0666666, -0.5343752, -0.6783857, -0.4953127, -0.7549486,
  -0.03958321, -0.0270834, 0.1039062, -0.2317708, -0.2726564, -0.4382811, 
    -0.6674478, -0.4380209, -0.4010417, -0.6020834, -0.8838542, -0.7059894, 
    -0.370573, -0.191927, -0.3268228, -0.4489584, -0.4710937, -0.217448, 
    -0.1442707, -0.08541679, -0.09843755, -0.4533854, -0.4059896, -0.4320312, 
    -0.4614584, -0.3260417, -0.4018228, -0.6307292, -0.7395835, -0.5859375, 
    -0.6671875, -0.917448, -0.9122398, -1.215365, -0.8914061, -0.8890624, 
    -1.158333, -1.320833, -0.8859372, -0.3742189, -0.09453106, -0.2929688, 
    -0.4554687, -0.6252608, -0.7315102, -0.3619795, -0.6937499, -1.066146, 
    -1.188281, -0.6747398, -0.1260417, -0.2242188, -0.7361979, -0.8783855, 
    -0.9979167, -1.069531, -1.149219, -0.9351563, -0.6083331, -0.5544271, 
    -0.6815102, -0.8078125, -0.4947917, -0.3140626, -0.1390624, -0.05338526, 
    -0.3984375, -0.6044273, -0.729948, -0.9549477, -0.9041669, -0.9242187, 
    -1.017969, -0.6182292, -1.091927, -1.423437, -1.403125, -1.011198, 
    -0.7434895, -0.2885416, 0.0739584, -0.09348965, -0.4151039, -0.3872399, 
    -0.2596354, 0.1627603, 0.3763022, 0.3289061, 0.6351562, 0.5713539, 
    0.2789061, -0.2106771, -0.2994792, -0.4065104, -0.5117188, -0.239583,
  0.0106771, 0.1434896, 0.04557288, -0.09583342, -0.2359375, -0.2440104, 
    -0.2638021, -0.1953125, -0.1927083, -0.1130208, -0.05520833, 0.03802073, 
    0.06171882, 0.03463542, 0.01614583, 0.005208373, 0.01406252, -0.03828126, 
    -0.1286458, -0.1330729, -0.1114584, -0.09557289, -0.1265625, -0.0703125, 
    0.01953125, -0.01197916, -0.1098958, -0.1572917, -0.1554688, -0.07291663, 
    -0.08333337, -0.09479165, -0.08255208, -0.1111979, 0.005729198, 
    0.04505205, -0.1049479, -0.1567708, -0.2567708, -0.2674479, -0.2921875, 
    -0.2986979, -0.2072917, -0.1049479, -0.0617187, -0.1005208, 0.02161455, 
    -0.1447916, -0.2692708, -0.3773438, -0.2916667, -0.2776041, -0.2992188, 
    -0.1768228, -0.2169271, -0.2494792, -0.2533854, -0.2624999, -0.3328125, 
    -0.2499999, -0.1385417, -0.1078125, -0.116927, -0.07864583, -0.05026042, 
    -0.08203125, -0.1630208, -0.1424479, -0.1320312, -0.2947916, -0.2179688, 
    -0.165625, -0.1588541, -0.225, -0.1757813, -0.373698, -0.3192708, 
    -0.3377604, -0.1809896, -0.171875, -0.2075521, -0.2632812, -0.1747396, 
    -0.1640625, -0.1346354, -0.08749998, 0.02942705, 0.08854163, 0.1117187, 
    0.1510416, 0.0953126, 0.1117188, 0.1419271, 0.08697915, -0.07656252, 
    -0.08880198,
  0.0078125, -0.007031262, -0.01276042, -0.01276042, -0.004947916, 
    -0.004947916, -0.005729169, -0.004427075, -0.006770834, -0.01432292, 
    -0.02213541, -0.034375, -0.03020833, -0.02630208, -0.01510417, 
    -0.001822911, -0.006510422, -0.008593753, -0.025, -0.02578125, 
    -0.02630208, -0.007031247, -0.0007812381, 0.01145834, 0.006510422, 
    -0.0007812455, -0.02109376, -0.02369791, -0.01432291, -0.01380208, 
    -0.03411458, -0.03932292, -0.04765625, -0.03880209, -0.02864583, 
    -0.02369791, -0.0078125, -0.02916667, -0.04270834, -0.04713541, 
    -0.07421874, -0.07604167, -0.06067708, -0.04531249, -0.02682292, 
    -0.01171875, 0.001302093, -0.008854166, -0.0234375, -0.01536459, 
    -0.02213542, -0.0234375, -0.03619792, -0.04947916, -0.04322918, 
    -0.03255208, -0.01848958, -0.005989581, -0.001041666, 0.004166663, 
    0.005468741, 0.01510417, 0.01536459, 0.01276042, -0.0109375, -0.03072917, 
    -0.02161459, -0.01067708, -0.01354167, -0.04244792, -0.04661458, 
    -0.04036459, -0.05052084, -0.040625, -0.040625, -0.04609375, -0.04453125, 
    -0.04973958, -0.03567709, -0.04270834, -0.07109375, -0.05989583, 
    -0.04453124, -0.02291667, -0.03333333, -0.03567708, -0.05286458, 
    -0.05989583, -0.04739584, -0.03723958, -0.03567708, -0.03697917, 
    -0.001822919, 0.03203125, 0.03151042, 0.01328124,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  -13.5979, -13.19714, -12.85965, -12.7229, -12.53696, -12.42682, -12.26822, 
    -12.01901, -11.80627, -11.66797, -11.61118, -11.58905, -11.35703, 
    -11.04141, -10.78464, -10.68127, -10.65051, -10.90964, -11.27499, 
    -11.63019, -12.04272, -12.41144, -12.91718, -13.29868, -13.57578, 
    -13.8125, -13.83435, -13.67578, -13.58542, -13.37033, -13.16537, 
    -13.03595, -12.90808, -12.69376, -12.34634, -11.95782, -11.54062, 
    -11.17447, -11.12915, -11.21899, -11.20572, -11.18228, -10.96094, 
    -10.72293, -10.59637, -10.54947, -10.75729, -10.99426, -11.37268, 
    -11.55807, -11.57239, -11.51016, -11.29037, -10.9263, -10.44348, 
    -10.18384, -9.941162, -9.898438, -10.27551, -10.87189, -11.64661, 
    -12.18933, -12.75104, -13.33957, -13.92657, -14.68829, -15.49478, 
    -16.33673, -16.82031, -17.35312, -17.94168, -18.16431, -18.44324, 
    -18.73462, -19.00677, -19.22708, -19.51587, -19.87759, -20.1409, 
    -20.34271, -20.52814, -20.5224, -20.49167, -20.45575, -20.43384, 
    -20.22162, -20.08047, -19.72995, -19.12033, -18.46744, -17.80914, 
    -17.14844, -16.26846, -15.34607, -14.63541, -14.09479,
  4.636719, 2.492462, -0.2486877, -2.956512, -5.634888, -7.459137, -8.830475, 
    -9.827606, -10.45496, -10.50674, -10.3349, -9.996094, -9.807526, 
    -10.22086, -10.73904, -11.37473, -11.74271, -12.18802, -12.69974, 
    -13.10599, -13.29688, -13.49454, -13.60025, -13.31848, -13.28098, 
    -13.61301, -13.65625, -13.58044, -12.99271, -12.01797, -11.08255, 
    -9.800781, -8.494019, -7.6362, -7.013275, -6.660675, -6.540375, 
    -5.813812, -4.509125, -2.780212, -1.62265, -0.7546692, -0.1453247, 
    -0.1278687, -0.2859497, -0.2539063, -0.1177063, 0.174469, 1.040894, 
    1.072388, 0.809906, 0.8028564, 0.3408813, -0.9083252, -2.618744, 
    -3.841675, -5.69635, -6.963531, -8.410431, -9.280731, -9.538788, 
    -9.254944, -9.420593, -8.894257, -8.333344, -7.292206, -6.722656, 
    -7.048187, -7.9953, -8.888306, -9.407532, -9.971863, -10.90286, 
    -11.73828, -13.1315, -14.43619, -14.76328, -14.34662, -13.70755, 
    -13.08282, -13.9198, -14.80807, -15.92709, -16.68671, -16.14584, 
    -14.50052, -12.24219, -10.56274, -8.215881, -5.263275, -2.192719, 
    0.4606628, 3.324768, 5.477081, 6.420837, 5.961456,
  -1.911194, -3.332031, -4.4198, -4.916901, -4.9729, -6.136719, -7.735657, 
    -9.47995, -11.24869, -13.01929, -14.26639, -16.18777, -17.39349, 
    -18.10104, -17.9646, -17.4487, -16.74295, -15.39505, -13.99271, 
    -13.11169, -12.58331, -13.18256, -14.26251, -13.57501, -12.43332, 
    -11.71353, -11.02319, -10.37241, -9.513794, -7.747406, -6.387512, 
    -5.445068, -5.319, -5.292694, -6.664581, -8.31485, -9.2901, -9.791931, 
    -8.988037, -6.852325, -5.641937, -4.890869, -4.063293, -3.145294, 
    -1.331787, 2.206268, 5.24115, 6.709625, 6.119537, 3.891388, 1.955475, 
    -0.2882996, -1.77005, -2.188538, -1.009399, 0.6726685, 2.820557, 
    4.562775, 3.969788, 1.722656, -0.7296753, -3.367188, -4.564056, 
    -3.898438, -3.54895, -1.401825, 1.308319, 1.927063, -0.2976379, 
    -3.685913, -5.633087, -5.529419, -5.23645, -6.315887, -7.875, -8.945038, 
    -9.374207, -10.54037, -11.04843, -10.59973, -9.17865, -8.11145, -7.6492, 
    -7.313812, -3.0242, 2.023163, 7.841156, 12.8573, 14.50546, 13.07864, 
    9.540619, 7.085144, 6.482025, 5.806488, 3.493225, 0.2184753,
  -13.55417, -15.25598, -14.67578, -11.94376, -8.574463, -6.458832, 
    -5.667969, -5.773438, -6.194794, -7.96225, -10.55441, -12.23956, 
    -12.74844, -11.91901, -12.07578, -9.633331, -7.907532, -8.045593, 
    -8.777893, -9.911224, -10.72733, -11.97891, -14.24429, -14.306, 
    -14.62372, -14.11771, -12.27631, -12.66797, -13.23386, -13.82837, 
    -13.09244, -12.82864, -11.92862, -11.31277, -11.28619, -12.22812, 
    -14.48151, -16.11951, -16.28073, -15.93826, -14.71979, -11.56039, 
    -8.280975, -3.742981, -2.396606, -4.152344, -8.158844, -7.297638, 
    -5.516937, -4.398438, -5.104156, -6.679443, -8.078888, -9.855469, 
    -8.242432, -3.576813, 4.615356, 9.233856, 10.60052, 9.044769, 3.6138, 
    -2.120819, -1.735931, -0.3609314, 1.931488, 5.94455, 10.37473, 14.42188, 
    13.52863, 6.9841, -0.258606, -3.892181, -3.345551, -3.553131, -5.761963, 
    -9.951294, -11.44611, -11.13565, -9.7883, -10.00833, -12.12891, 
    -13.37866, -14.43387, -13.73721, -9.224213, -5.132263, -1.7164, 
    -0.09063721, -0.9265747, -0.9338684, -3.42215, -5.43985, -6.014832, 
    -7.893219, -10.72342, -11.51666,
  -14.52866, -17.47916, -17.66119, -15.50311, -11.11093, -7.806244, 
    -7.605988, -6.68985, -7.330719, -7.742432, -8.490875, -6.434875, 
    -5.378113, -8.264587, -9.931, -9.2388, -7.690125, -4.802368, -3.860138, 
    -3.998444, -5.654419, -5.167694, -5.246094, -7.639038, -9.238556, 
    -8.034363, -8.854431, -10.51614, -10.03201, -10.03152, -10.64166, 
    -11.27448, -10.69635, -9.969299, -8.782043, -8.003906, -6.679169, 
    -8.154694, -9.997894, -11.96222, -14.23648, -16.34973, -16.32422, 
    -17.61691, -18.59482, -19.86121, -19.52216, -21.12527, -18.806, 
    -15.08957, -8.894012, -4.097656, -4.875793, -7.113831, -6.677612, 
    -4.867981, -3.266388, -3.463531, -4.572113, -6.92395, -9.758331, 
    -11.24039, -9.189575, -8.277618, -7.484375, -6.520294, -6.649506, 
    -4.090637, -3.060944, -2.278381, -3.68515, -9.317719, -9.231262, 
    -10.54245, -13.51407, -10.98203, -3.869019, -4.210175, -8.663788, 
    -10.38541, -11.53802, -12.2724, -9.769012, -8.092712, -6.820068, 
    -5.231262, -4.457794, -4.363281, -3.481506, -3.683319, -6.563019, 
    -6.212769, -8.511719, -6.806488, -6.413788, -9.677094,
  -14.43857, -18.68411, -10.01694, -6.12915, 0.3093567, 4.460693, 2.966125, 
    -3.817963, -9.296875, -11.09064, -10.71118, -11.21146, -10.64896, 
    -9.494537, -6.471893, -4.305969, -2.050781, -0.3544312, -2.58725, 
    -4.279968, -3.891937, -6.417725, -12.05313, -17.52448, -15.69296, 
    -14.15442, -14.51434, -15.0849, -12.78543, -8.590118, -5.876556, 
    -6.322937, -6.070557, -6.274506, -4.789307, -4.45755, -6.595032, 
    -7.978119, -8.293518, -7.2453, -9.268768, -13.88516, -19.16379, 
    -18.47501, -14.63544, -13.11093, -13.3013, -15.47919, -15.14191, 
    -12.93463, -8.436462, -5.346619, -5.208069, -8.842957, -9.232025, 
    -4.985443, -3.47345, -3.992706, -6.384613, -9.970306, -12.89999, 
    -14.98828, -17.46823, -20.7789, -24.15833, -25.04871, -21.53387, 
    -19.46927, -22.7164, -26.70079, -24.36278, -18.76483, -22.38098, 
    -23.37552, -25.70862, -22.42056, -14.55026, -7.993744, -10.12943, 
    -10.36771, -10.0177, -8.893494, -9.223419, -9.743225, -13.82681, 
    -16.21042, -12.9086, -9.5784, -7.060425, -7.185394, -10.53464, -14.24481, 
    -15.53906, -12.66431, -8.712738, -9.744019,
  -17.8013, -17.03049, -14.48438, -15.28308, -18.17499, -25.27267, -32.67917, 
    -35.19141, -33.91431, -26.62811, -24.59845, -23.76926, -21.53021, 
    -16.80624, -13.50052, -13.94949, -17.32211, -19.3349, -18.19193, 
    -13.82916, -10.61014, -11.42136, -13.49533, -14.86224, -15.16406, 
    -12.84634, -17.46484, -21.34949, -19.06744, -12.74142, -9.670319, 
    -10.59427, -15.35001, -14.87552, -9.086212, -4.262238, -12.40964, 
    -21.31042, -26.11902, -23.07629, -20.06433, -21.21901, -20.73904, 
    -14.64479, -4.154419, 1.136459, -1.835678, -4.336472, -8.393753, 
    -7.172394, -0.9682159, 1.0336, 1.970825, -0.0385437, 3.026825, 7.507813, 
    9.1521, 2.629944, -6.811188, -9.03125, -10.76511, -13.05209, -21.26457, 
    -27.30859, -28.8, -23.69505, -14.02162, -13.74323, -17.02266, -20.35416, 
    -20.0388, -18.9828, -22.58229, -26.74454, -31.17267, -34.06563, 
    -34.54271, -34.34428, -38.13751, -48.42812, -46.26511, -36.68724, 
    -29.77032, -31.67474, -40.62109, -41.96146, -37.65469, -33.35156, 
    -32.45419, -30.40079, -26.42892, -23.64426, -22.38748, -22.62241, 
    -23.31641, -21.22214,
  -45.56122, -41.55704, -37.40625, -41.80807, -46.39764, -50.70181, 
    -50.73907, -45.42969, -43.2151, -48.81042, -51.22136, -52.46744, 
    -54.08696, -55.30443, -49.61978, -42.04376, -38.38072, -37.47945, 
    -36.29428, -38.20079, -35.39661, -32.40598, -35.57162, -36.72083, 
    -34.36069, -31.99062, -26.83333, -24.01746, -18.46536, -13.64844, 
    -12.92265, -12.89948, -15.12448, -14.80652, -10.22736, -5.910934, 
    -6.628128, -3.190887, -6.172913, -6.076294, -4.079681, -2.289322, 
    -0.4466248, 1.219528, -0.2184906, -5.676559, -11.47214, -13.25755, 
    -9.867966, -10.06276, -10.31796, -7.352341, -4.797653, -8.427078, 
    -6.232285, -3.199997, -2.926041, -7.45079, -15.2263, -14.43985, 
    -4.313293, -1.818497, -2.543228, -0.9794159, 1.535675, 2.712509, 
    1.388535, -1.046082, -3.154419, -5.873444, -7.088547, -6.211975, 
    -7.335419, -6.830475, -7.5961, -13.375, -18.96562, -16.54428, -13.84271, 
    -13.15416, -11.9828, -11.925, -11.00781, -17.34975, -22.67865, -30.82292, 
    -36.56406, -43.8078, -48.74426, -46.70729, -44.53645, -45.94141, 
    -50.47137, -52.10675, -54.07291, -51.44193,
  -22.88957, -21.26277, -16.77423, -16.6375, -21.87578, -21.72423, -18.05365, 
    -13.15781, -13.3336, -15.40546, -18.66953, -12.8284, -10.25548, 
    -7.590622, -6.834122, -6.356522, -9.484894, -9.985931, -10.98671, 
    -8.163544, -7.844528, -11.11952, -17.37578, -18.63646, -12.36433, 
    -8.456253, -10.21327, -12.42319, -13.02553, -11.7948, -8.276047, 
    -4.01796, -1.915634, -6.850784, -6.902603, -9.645584, -7.569275, 
    -2.591415, -7.313538, -14.50052, -13.38905, -5.275269, -6.334381, 
    -11.3573, -12.95859, -13.89505, -13.95444, -8.297913, -6.482819, 
    -12.06302, -17.05443, -13.52682, -5.766403, -9.615631, -11.58229, 
    -7.195313, -0.9648438, -5.938278, -13.16953, -10.56354, -5.29686, 
    -8.70755, -9.936462, -2.275269, -1.692963, -3.740891, 0.7083435, 
    1.206253, -0.8562469, -0.7335968, -0.3403625, -2.913025, -7.016663, 
    -6.293243, -2.834885, -6.696869, -8.394791, -13.19844, -12.02057, 
    -9.996094, -14.27838, -16.06458, -17.24504, -17.3474, -10.5909, 
    -9.851822, -8.086975, -10.92578, -14.42422, -14.84766, -17.76198, 
    -28.86952, -31.73878, -30.24113, -23.47031, -22.25209,
  -18.94766, -11.38985, -7.449478, -8.763809, -6.722916, -1.157288, 
    0.5122375, 1.911194, 3.649734, -0.1820221, -10.81667, -11.43517, 
    -10.21251, -7.679947, -5.067184, -9.576569, -8.989853, -5.937759, 
    -2.858337, -7.980209, -9.197388, -8.893234, -8.779175, -3.647644, 
    -3.224991, -4.041138, -10.91458, -14.13203, -12.8922, -8.420578, 
    -5.245834, -5.338806, -3.024216, -3.594269, -5.209122, -9.595047, 
    -4.791412, -3.040619, -4.282028, -9.414063, -7.802078, -6.156525, 
    -1.291153, -8.424225, -10.16119, -2.724487, -2.697922, -2.248428, 
    -2.305466, -1.398956, -7.717712, -3.973694, 2.042969, -3.86145, 
    -6.552078, -2.422928, -0.5734253, -5.611465, -4.517715, -0.5924683, 
    0.2174377, -4.693756, -2.032547, -1.655731, -4.921097, -6.280457, 
    -0.1598969, 2.428131, -2.471085, -6.631516, -1.403915, 0.5619659, 
    0.7239532, 5.594788, 3.159103, -4.452866, -11.82864, -11.6974, -13.25781, 
    -4.181274, 2.351807, 2.028656, -8.394272, -16.89558, -12.57629, 
    -7.451553, -4.162247, -7.661453, -8.245575, -4.173691, -10.28906, 
    -14.99739, -10.60234, -5.149994, -10.46327, -17.36642,
  -3.976563, -7.9552, -5.402328, -3.351563, 2.469788, -0.0304718, -9.653107, 
    -8.986465, -5.235687, -5.890106, -6.304413, -6.108322, -2.892441, 
    -4.605484, -8.787491, -3.919022, -0.06640625, 3.286209, 1.765884, 
    1.434372, -2.141403, -5.913788, -8.340103, -7.935425, -5.507553, 
    -6.123962, -9.533844, -5.741653, -1.844009, -1.088287, -4.358322, 
    -7.748169, -5.355743, -2.690887, -2.927353, 4.802872, 2.606781, 
    -0.5211029, 1.091919, -1.757568, -6.559906, -7.242706, -2.95575, 
    4.680969, 6.9487, 4.119019, 9.094788, 1.142181, -5.978149, -0.1138, 
    -1.573425, -4.448181, -4.409882, -10.8862, -14.68594, -11.68567, 
    -5.905457, -3.759628, -4.501831, -6.760925, -8.169266, -4.608582, 
    -1.308838, 0.3151093, -3.493225, -5.517975, -4.128632, 2.052078, 
    -0.7122345, 1.375275, -0.433075, -1.610947, 0.6575623, 2.649719, 
    -5.210175, -10.50105, -6.690628, 6.728897, 6.360931, 8.808594, 7.560944, 
    5.030457, 0.660675, -3.184631, -8.9151, -6.833588, -6.14505, -6.374756, 
    -4.546112, -0.7890472, -1.402344, -5.041138, -4.270828, -2.905991, 
    -9.410416, -7.870834,
  -0.6851501, -5.362244, -2.494537, 1.798706, -1.732025, -1.813263, 3.920044, 
    10.22083, 5.820862, -1.106537, 4.086975, 10.48514, 8.199768, 1.675018, 
    -3.267731, 0.5716248, 3.255981, 0.2304688, -2.040863, 1.773956, 7.701019, 
    1.983093, -1.551056, 4.003632, 6.050537, 4.563293, 3.82785, 7.020569, 
    4.532532, 9.479401, 11.66147, 8.102356, 11.00391, 10.12238, 5.237244, 
    7.710175, 17.31824, 12.97632, 7.865631, 4.2547, 2.157806, 8.854675, 
    6.88385, 3.279938, -1.948975, -0.3617249, 7.944519, 8.85495, 0.6820374, 
    5.387512, 7.199738, 1.286743, -2.692688, -5.192444, -0.09609985, 
    4.413544, 4.259125, 3.564056, 3.816162, -1.704163, 0.6065063, 6.731506, 
    -0.5640564, -5.155182, 2.181793, 1.065094, 2.308075, 3.625519, 3.964325, 
    4.803375, 1.944, -1.805481, 4.174225, -0.524231, -3.134644, 2.304688, 
    11.7164, 27.99036, 23.37317, 11.15784, 6.960938, 7.501038, 7.9953, 
    7.438293, 5.627075, 7.566406, 5.745819, 0.3994751, -4.321625, -3.134369, 
    4.024994, 3.609894, 2.945587, -2.113525, 0.1947632, 3.337494,
  -0.3820496, 5.4841, 11.52292, 3.810425, 5.330475, 11.05338, 8.374237, 
    9.843475, 9.082031, 6.68335, 10.31119, 12.19662, 6.672638, 3.175262, 
    3.954407, 10.72577, 7.880981, 0.5721436, 1.351837, 6.359894, 9.949738, 
    8.322906, 7.066406, 12.7052, 17.02579, 15.62656, 17.23569, 16.42944, 
    15.97318, 19.05835, 18.5401, 21.62213, 24.95496, 20.38617, 20.49844, 
    23.14948, 19.68073, 9.742462, 15.04895, 16.90311, 8.078369, 6.229431, 
    2.345062, 2.102081, 2.283844, 7.184662, 20.38907, 17.05963, 15.87344, 
    15.58853, 18.79871, 10.87683, 10.80389, 10.18726, 16.04141, 21.39999, 
    11.05026, 0.8544312, -1.664307, 3.414063, 2.460144, 0.8815308, 0.3424377, 
    6.348694, 9.016937, 2.06485, 1.980225, 1.425507, 2.223419, 9.759644, 
    8.825256, 10.93124, 17.50833, 11.70236, 13.94272, 22.3367, 25.29166, 
    37.25807, 35.68073, 9.179443, 10.91043, 6.941132, 0.53125, 5.179688, 
    4.420563, 7.211487, 7.990631, 0.8731689, 2.070831, 7.427582, 4.378113, 
    1.983093, 6.553131, 5.790863, 2.698181, 2.095032,
  -3.24765, 1.371887, 11.8862, 14.08072, 11.96561, 6.255463, 6.450256, 
    7.378113, 7.097931, 5.411987, 6.288788, 9.278137, 13.74948, 19.66669, 
    10.04062, 13.86435, 14.90988, 5.536743, 14.59869, 10.71121, 8.394775, 
    11.92734, 8.054169, 11.45679, 8.218506, 7.067719, 11.14246, 7.985687, 
    10.24191, 12.80392, 14.28827, 15.19556, 6.081757, 10.70572, 15.48386, 
    12.71249, 10.41275, 12.54349, 29.38593, 36.28281, 12.75287, 3.537231, 
    -0.799469, 3.693756, 3.361206, 4.812225, 14.68411, 19.75964, 15.18829, 
    10.03699, 7.874451, 11.09686, 15.67554, 18.40417, 16.44949, 16.7453, 
    10.52084, 3.863037, 4.767181, 3.534119, 0.7437439, 4.939575, 3.264557, 
    2.888031, -0.2437439, 0.7987061, 4.934387, 4.999237, 1.713806, 8.645569, 
    4.496368, 5.855194, 11.7388, 6.96875, 8.060699, 8.621368, 19.28049, 
    33.22293, 13.38074, 0.8551941, 3.857025, -2.0466, -4.154694, -2.558075, 
    4.564331, 1.738281, -3.617188, -0.2888184, 2.622375, 3.290375, -1.075012, 
    3.417969, 6.902618, 8.856262, 6.083069, 0.9489746,
  -0.7690125, 3.314056, 5.125, 3.67395, -0.2520752, 0.940094, -1.525787, 
    -3.506775, -0.6653442, -1.188019, 9.3974, 13.65155, 5.432312, 8.753387, 
    4.265869, 7.645844, 9.393219, 5.023163, 7.9776, -0.7645874, -1.652863, 
    2.422638, -4.855469, -5.400238, -7.953125, -1.685944, 0.8145752, 
    -5.534119, -0.475769, -3.61145, 7.078888, 12.90625, 3.29895, 7.113556, 
    2.1922, 0.3528748, 11.22293, 15.44113, 21.58594, 15.71902, 2.297668, 
    -8.660156, -5.77005, -4.65625, 1.220581, 8.514343, 6.029419, 5.509613, 
    3.754944, 5.832031, 4.279938, 9.060944, 9.167969, 3.445831, 5.908325, 
    4.018219, -0.2166748, 5.547668, 6.4039, 5.978638, 0.1984253, 1.688019, 
    7.856262, 2.822632, 7.523438, 6.622131, 1.274994, -0.5273438, 1.500793, 
    -2.243225, -0.4710999, -0.8234558, -4.645325, -2.246368, 4.641663, 
    0.7984619, 6.551575, 6.518219, -8.478912, -14.45053, -15.27292, 
    -9.968475, -15.83203, -11.3284, -7.017456, -12.53934, -15.71249, 
    -9.210938, -0.5739441, -2.508087, -3.896088, -1.666931, -5.302582, 
    -1.527344, 0.9817505, -5.259369,
  2.571106, -0.4114685, -2.95105, 0.7140503, 2.163269, 0.7992249, -1.570831, 
    -15.70676, -28.4534, -10.21094, -2.181244, -2.273956, -7.088287, 
    -6.543762, -6.334625, -5.252594, -0.5604248, 0.8052063, 0.04504395, 
    -9.018463, -9.2948, -5.797638, -2.777069, -9.22345, -10.10468, -7.287506, 
    -6.997131, -4.911194, 0.7489624, 0.7276001, 8.691681, 3.919037, 
    -5.421082, -6.826324, -3.180756, 3.172913, -1.736206, -0.3812561, 
    6.527344, -0.8104248, -9.465881, -15.19583, -9.148193, -3.073456, 
    -2.659912, -1.618225, -3.982574, -1.762756, -2.760681, -0.2505188, 
    -0.6906433, 2.532562, 0.2036438, 2.629944, -4.125519, -6.549469, 
    -3.887268, 5.104401, 5.194519, 2.547394, 2.431, 0.151825, 6.079437, 
    4.545593, 4.090637, -1.984131, -10.92526, -5.958862, -3.8685, -6.765625, 
    -4.721863, -2.32135, -7.48645, -0.9286499, 3.729431, -4.264343, 
    -5.082794, -7.557556, -10.39246, -18.83438, -21.55338, -14.33179, 
    -23.2406, -18.27344, -17.42682, -14.02759, -13.02863, -14.30157, 
    -7.002106, -4.0896, -3.356506, -3.878113, -4.331238, -4.556244, 
    -2.372131, -0.2458191,
  -3.50885, -3.713013, -1.238556, -6.788025, -3.33725, -7.296875, -11.944, 
    -24.79608, -26.28752, -14.49554, -12.26746, -7.836182, -8.365356, 
    -8.492432, -7.777344, -10.28021, -8.702606, -6.928131, -7.186188, 
    -7.723969, -8.657562, -7.285675, -10.74191, -7.193726, -5.840363, 
    -3.493225, -3.515869, 4.884369, 8.94635, 4.671356, 1.880463, -5.308594, 
    -14.62372, -8.835175, -5.483063, -2.058075, -1.25885, -2.617981, 
    -3.247162, -6.914581, -11.81458, -16.10101, -3.94635, -0.9049683, 
    -0.497406, -1.651825, -4.226563, -7.997681, -7.393738, -8.971069, 
    -9.985168, -9.892181, -11.05157, -9.86615, -2.306519, 7.925781, 8.447144, 
    12.15079, 11.03384, 4.9021, 4.784637, 3.7164, 0.3999939, -5.45105, 
    -5.841919, -11.08127, -8.673431, -10.48099, -12.11771, -6.914063, 
    -6.20105, -5.2724, 0.2166748, -2.200531, -9.492188, -4.685944, -4.646606, 
    -8.281799, -0.5036621, -3.581787, -26.0737, -8.786469, -17.48256, 
    -24.6078, -17.59479, -9.912994, -4.884125, -2.191406, -0.772644, 
    -0.2744751, -1.565613, -1.341644, -2.332825, 1.94635, -3.515625, 0.3364563,
  -3.829407, 0.52005, -11.51718, -5.6362, -4.087738, -7.694519, -15.92343, 
    -13.93854, -7.688812, -10.00626, -7.844513, -9.861725, -8.015625, 
    -3.709625, -3.366913, -5.841125, -8.371094, -6.169769, -4.0466, 
    -0.6455688, -5.253906, -10.56226, -10.62943, -1.992432, -0.7229309, 
    4.780212, 2.765381, 6.171875, 6.136993, 0.6411438, -5.188538, -7.592712, 
    -5.701813, -4.210693, -4.334106, -2.917969, -1.257294, -5.03125, 
    -3.271362, -3.44455, -5.823456, -3.100006, 3.59375, 3.124756, 5.389862, 
    -6.138, -10.68542, -12.59686, -10.94165, -10.49973, -7.191681, -11.12369, 
    -4.974457, -1.916656, 6.118744, 16.16327, 14.69272, 9.09375, 11.34558, 
    12.48541, 6.018738, -4.722137, -14.34244, -17.44193, -18.07291, 
    -20.92371, -20.57733, -19.13986, -8.195038, -6.855469, -0.4054871, 
    4.582825, -4.736694, -5.870056, -1.043732, 4.802063, -4.079681, -7.88385, 
    21.00131, 3.810684, -15.62762, 12.11954, 7.414581, 7.638794, -4.516663, 
    -3.125763, -0.7223816, 5.918488, 1.184631, -10.13931, -10.10416, 
    -5.101807, 0.6640625, 4.088013, 2.756256, 3.199493,
  -2.4953, -6.716675, -10.80341, -3.945313, -2.262756, -9.760681, -11.52914, 
    -6.05365, -8.760925, -7.194275, -5.889832, -10.47214, -13.66432, 
    -5.165619, -1.120331, 3.322144, -4.934387, -7.835938, -6.24115, 
    -5.297913, -5.059357, -9.43515, -6.335419, -5.133331, 1.2659, 5.977631, 
    13.68152, 8.722931, 5.730225, 1.14505, -7.449738, -4.408569, 0.7052307, 
    0.3109436, -0.4924622, -1.990082, -1.922638, -5.665863, -4.891937, 
    -0.9664001, -0.2210999, 7.648987, 1.116913, 0.0854187, -1.7117, 
    -7.775513, -3.67865, -5.888, -9.452332, -10.27188, -6.740631, -2.6026, 
    -2.300781, 14.75809, 20.00754, 15.70544, 12.57446, 7.61145, 5.788025, 
    -2.189606, -7.411713, -19.56094, -21.94507, -26.60571, -27.23724, 
    -19.91302, -14.55649, -7.380707, 1.17395, 4.721863, 3.271606, 4.059906, 
    -3.827332, 10.34766, 11.86642, -8.63385, -4.253113, -3.892456, 36.37524, 
    23.9677, -1.514862, 11.17056, 5.257019, 18.56146, 20.4138, 25.52943, 
    10.83984, -0.7593689, -6.553894, -7.618744, -6.73465, -5.329956, 
    -1.661743, 3.401306, 5.018494, 1.508057,
  3.995575, -4.761444, 5.445313, -1.252594, -2.682312, -13.87918, -13.11407, 
    -3.695038, -7.025787, 1.483856, 3.856506, -5.667175, -12.25887, 
    0.1315002, 1.265625, -2.010406, -7.299988, -8.2258, -1.720825, -3.720825, 
    -0.7098999, -7.764587, -2.148956, -0.9505005, 1.96225, 9.780487, 
    10.40936, 4.400787, -0.3135376, -4.020569, -5.317963, -5.24115, 
    -4.638275, 0.227356, 0.04846191, -2.72345, -3.623718, -3.106232, 
    -3.240631, 0.1653442, 0.9312439, 2.64035, 2.444519, -1.071625, -2.198456, 
    -1.303406, -2.121887, -6.931244, -11.51535, -11.46927, -8.867172, 
    -3.033569, -3.276047, 1.210419, 2.227325, -0.8864441, -7.443237, 
    -4.491913, -11.64481, -13.04037, -17.4328, -21.0401, -16.22159, 
    -17.16147, -15.59637, -8.740112, -6.634613, 0.8562317, 4.517975, 
    8.064819, 5.341431, 6.350525, 8.3461, 11.11353, -5.329437, -1.283325, 
    -3.360931, 22.16953, 53.30313, 12.55626, 4.397125, 15.80676, 12.49298, 
    16.1237, 28.19296, 34.1375, 0.4921875, -4.406769, -9.617432, -7.740875, 
    -6.900238, -4.335693, 0.3166809, 2.963806, 5.873444, 1.041412,
  7.643738, 8.851044, 5.634888, 4.910156, 3.964844, -3.011719, -6.943222, 
    -4.5336, 4.030731, 18.62422, 24.48619, 11.35938, 2.217194, -1.993744, 
    -0.1963501, -1.942963, -8.348419, -4.547119, -4.372406, -3.132019, 
    -0.9190063, -0.4505005, -0.2833557, 1.277588, -2.067719, 3.377594, 
    1.018219, 5.950531, 0.669281, -7.979431, -7.235138, -5.374207, -9.40625, 
    -4.072388, -4.999481, -6.367462, -4.711975, -8.000519, -10.49063, 
    -1.033569, -1.466156, -0.8453064, 0.2526245, -8.621887, -3.637238, 
    -7.851563, -6.202606, -8.845306, -9.982559, -15.84871, -21.65677, 
    -18.43463, -8.491653, -4.94635, -5.009628, -8.830719, -6.045593, 
    -6.797943, -10.40598, -15.83774, -20.70703, -18.67163, -16.97162, 
    -14.84479, -9.771362, -1.766937, 1.694794, 9.160675, 7.823441, 8.217697, 
    9.834381, 6.952332, 10.83646, 5.49765, -3.867981, -5.105988, -6.477341, 
    11.01094, 22.16068, 9.480972, 13.98749, 15.96875, 20.18437, 12.78751, 
    25.56433, 22.92499, -3.361969, -3.69165, -2.560394, -5.404694, 
    -0.05911255, 3.414063, 2.111206, 7.5289, 8.821625, 8.492706,
  11.67319, 11.3284, 5.769531, 0.7354126, 7.298691, 12.07109, 1.371094, 
    -7.259903, 6.651047, 29.37968, 15.18933, 6.68985, 10.18958, 6.091415, 
    -0.2369843, 0.3049469, -3.289581, -2.939606, -6.727844, -4.048462, 
    0.7963562, 5.894531, 0.9138184, 1.916412, 3.203125, 4.653107, 3.599243, 
    0.3976746, -3.0802, -2.859131, -6.508606, -9.027344, -5.47525, -6.336731, 
    0.1601563, -6.378632, -5.457825, -6.388794, -12.57187, -2.178894, 
    -5.644531, -13.67891, -10.89531, -24.07603, -26.49976, -17.96172, 
    -15.24895, -11.84818, -11.97266, -16.54193, -16.5237, -23.00494, 
    -16.10938, -1.905731, -7.547134, -11.05833, -7.987228, -3.974457, 
    -7.019806, -11.51953, -12.47736, -10.26379, -7.680481, -6.528412, 
    -3.941406, 0.6752625, 10.10651, 12.03151, 13.23776, 13.40288, 16.50626, 
    11.12994, 9.297668, 7.704712, -10.55444, -14.48254, 6.404686, 26.35938, 
    11.61484, 18.04141, 14.78619, 8.257034, 20.77449, 13.6198, 2.442703, 
    5.367981, 1.875, -1.535675, -0.4031372, -4.884369, -0.5135498, 1.422668, 
    5.784119, 7.54425, 9.748962, 14.31354,
  -2.191132, 0.5830994, -5.729431, -11.47003, -2.484634, 6.411972, 4.711212, 
    4.077866, -1.314575, 12.45313, -0.1927032, 3.365356, 24.37943, 26.13333, 
    9.392197, 1.516937, -5.533859, -5.382813, -0.3479156, -4.308594, 
    4.845062, 3.853638, 1.058319, -3.414581, -3.045563, -7.963287, -10.69894, 
    -15.95912, -13.38254, -4.011963, -2.555725, -6.788544, -7.115356, 
    -6.527863, -4.942444, -5.821869, -5.152863, 17.27605, 3.136719, 
    -16.49088, -24.82996, -21.38412, -18.02577, -23.16068, -29.17839, 
    -27.46719, -24.52629, -29.91068, -28.20001, -26.32733, -32.57761, 
    -38.61432, -36.13231, -33.24271, -32.20078, -32.03227, -29.13774, 
    -23.92787, -21.98619, -16.88307, -16.36069, -15.66718, -7.434113, 
    -4.551819, -1.19635, 2.02655, 2.345825, 4.130188, 7.384125, 3.256775, 
    2.195557, -0.8505249, -7.026306, -4.454956, -9.481506, 21.89401, 
    23.08775, 17.42369, 20.96277, 9.800781, 18.20886, 19.10234, 21.31511, 
    10.68306, -5.328644, -10.33151, -0.5112, -1.256531, -2.337494, -3.31485, 
    -2.868225, 1.942719, 3.701843, 2.776825, 1.499481, 1.101044,
  -6.958344, -5.619812, -6.420044, -0.5635376, 2.21875, 6.927338, 8.810936, 
    9.1138, -5.637764, -17.04921, -12.54219, 4.668488, 20.24661, 27.81093, 
    23.41901, 16.31537, -0.6244812, -3.448441, 1.105743, -2.230469, 4.35704, 
    8.664581, 5.726303, -4.279953, -5.354416, -9.104691, -6.982559, 
    -4.543762, -2.867966, -3.481247, -2.165359, -21.31693, -27.51093, 
    -15.68047, -10.67787, -7.557281, -12.78542, -4.458595, -6.921616, 
    -21.25702, -19.37994, -17.58437, -14.92213, -13.33932, -16.80208, 
    -23.80026, -26.53828, -30.60027, -27.35027, -25.07864, -25.04428, 
    -23.63829, -28.21535, -26.20573, -24.9323, -23.73669, -23.21121, 
    -22.37915, -21.08255, -18.21927, -14.94583, -14.02631, -11.05676, 
    -12.36511, -7.56015, -10.70233, -7.520599, -7.900269, -6.274994, 
    -8.678925, -5.077866, -11.99402, -12.42682, -9.592438, 11.81302, 
    18.50156, 1.702087, 5.240616, 7.120834, 6.862503, 20.22656, 15.84167, 
    9.565613, 11.56042, 4.517456, -4.936432, -2.061188, 0.2583313, -1.177338, 
    -3.433594, -5.219513, -3.465363, -1.698181, -2.578888, -3.984894, 
    -4.390106,
  -7.005981, -5.111984, 4.019272, 22.85261, 5.429169, -0.6138, -8.851303, 
    -14.66145, -20.74844, -13.95757, -11.07239, -5.481781, 8.579178, 
    10.32031, 8.855209, 10.52553, 3.945053, 8.591141, 12.33464, 9.785675, 
    11.24896, 6.948181, 5.729431, 2.526031, -6.864578, -16.3289, -19.01277, 
    10.37891, 6.030991, 7.340622, -4.413269, -12.45808, -3.407814, -11.38515, 
    -5.210678, -7.412247, -12.19453, -13.54845, -9.468491, -4.230988, 
    0.183075, 2.429947, 5.635162, 10.30495, 8.249741, -2.853394, -6.957031, 
    -7.136719, -10.94531, -11.84869, -17.12447, -13.69402, -13.58307, 
    -14.97916, -13.35886, -19.98438, -19.70209, -22.27888, -18.13411, 
    -24.12422, -16.67422, -12.18152, -11.68567, -7.899231, -8.323975, 
    -5.548431, -5.519531, -8.023697, -1.705734, -1.340881, -3.273438, 
    -2.56015, -7.574219, -26.70338, -23.69766, -3.618752, -11.19087, 
    -5.96666, -11.19063, 9.060928, 11.88022, 11.63855, 13.76849, 5.601822, 
    3.730713, 9.483597, 5.892441, 6.563019, 3.205734, 2.891403, 1.612762, 
    1.458862, 4.628113, 3.222382, -1.590103, -7.245331,
  -5.065872, -5.9487, 0.670578, -0.2585907, -10.67839, -7.795319, -9.639847, 
    -12.2039, -8.394791, -6.864075, -28.04166, -17.91223, -7.030197, 
    3.096603, 0.0921936, -6.771606, -0.3609314, 3.907288, 4.453903, 4.330475, 
    -0.4187469, -1.954681, 1.587494, 0.4252625, -1.589325, -11.45, -11.30704, 
    12.79741, 15.30025, 13.96405, 10.30495, 15.97656, 8.3461, -3.737503, 
    -1.568741, -8.335938, -13.39531, -7.576035, -2.383865, 0.7505188, 
    4.578125, 4.478912, 7.651031, 7.215622, 6.001816, 5.143753, 7.056503, 
    5.000519, 9.349213, 9.147125, 4.047134, 4.691406, 9.039581, 9.189575, 
    11.23438, 9.783585, 9.513031, 9.80574, 8.241669, 8.732559, 5.779694, 
    4.533585, 7.067184, 7.729172, 6.182297, 2.127609, 3.109375, 0.8018341, 
    1.877869, 4.733063, 10.60339, 11.22266, 3.52005, -7.803131, -13.51535, 
    -15.49974, 5.833069, 11.8474, -5.264328, 30.84427, 18.5211, 20.56198, 
    9.451035, 4.295044, 6.452072, 9.859909, 6.742462, 7.221359, 6.999741, 
    5.29921, 3.848694, 0.9200439, -0.776062, -3.720306, -6.078903, -5.896103,
  -6.970322, -8.353119, -7.003891, -9.623703, -10.86536, -7.837234, 
    -6.948959, -7.270828, -7.717178, -12.24767, -35.61093, -19.50365, 
    -10.13802, -3.141922, 4.875519, -4.346619, -0.8190155, -0.4046936, 
    0.1765594, -8.261719, -12.62917, -1.00885, 10.30598, 7.951553, 9.639069, 
    4.53801, -1.54895, 0.6018219, 6.847916, 10.77448, 18.64662, 18.14114, 
    11.16328, 17.78308, 11.09584, 0.02656555, -3.385925, 0.1187592, 2.148697, 
    1.967438, 0.4729156, -2.003387, 0.9908905, 2.762497, 3.632553, 3.599991, 
    5.039063, 7.575775, 11.98463, 10.42317, 12.35156, 14.40912, 14.07474, 
    17.85208, 21.79478, 25.94766, 29.90077, 32.50079, 30.53047, 27.36121, 
    22.20729, 18.68724, 18.15312, 9.904953, 5.630722, 5.625259, 7.177078, 
    4.847916, 4.804947, 5.207809, 12.2211, 2.182816, -1.056778, -0.8244781, 
    8.467957, 7.579956, 24.32188, 20.83751, 11.96875, 23.88879, 12.02083, 
    8.039597, 3.5914, 3.108597, 7.328384, 5.043228, 5.470581, 4.273697, 
    2.090118, -4.640884, -2.71225, -2.759109, -3.495819, -7.054169, 
    -7.705215, -8.852081,
  -8.348434, -9.271606, -10.31146, -9.880203, -7.756241, -6.129166, 
    -6.517181, -6.616928, -5.337769, -9.992706, -17.82083, -9.749741, 
    -9.381256, -2.635162, 5.138794, 1.931, 2.969009, 3.903381, -1.690369, 
    -9.321091, -10.95624, 11.82031, 10.98749, 4.558594, 14.66016, 7.21875, 
    -3.972137, -3.5802, 16.95468, 19.24036, 10.13124, 5.108856, 6.483582, 
    20.82213, 11.1302, 7.351044, 5.450516, 3.055206, 1.034637, 3.192963, 
    -0.3638, 2.835159, 5.873962, 5.970566, 7.995041, 5.7276, 4.878128, 
    3.84375, 6.334641, 6.603119, 9.832809, 10.65077, 7.756775, 10.90573, 
    11.73489, 15.51405, 14.80495, 16.88098, 12.30859, 9.066147, 10.23515, 
    9.545319, 9.266144, 8.484116, 5.431503, 1.092453, 0.8085938, 2.585938, 
    0.674469, -0.72995, 1.962509, -4.590103, -2.4375, 19.29713, 8.268494, 
    -1.746353, -0.9463501, 2.921616, 5.181519, 6.060425, 5.067184, 3.983597, 
    6.503128, -0.0158844, 0.5408936, 4.761719, 5.463013, 9.314331, 2.457809, 
    1.111206, -1.750519, -3.861191, -6.802856, -4.09166, -5.11615, -8.179947,
  -6.00885, -6.209106, -7.044281, -7.528656, -6.826035, -6.887238, -7.459122, 
    -5.515884, -5.153641, -5.821625, -11.47005, -9.039063, -8.617188, 
    -7.644012, -3.879944, -0.1908875, 1.862244, -0.1929626, -1.570572, 
    -4.889069, -10.48047, -3.176559, 0.295578, -2.271362, 6.702087, 0.97995, 
    -5.695053, -4.803391, 8.091934, 8.09375, 5.992966, 13.12552, 5.310425, 
    9.384369, 8.054169, 4.715103, 1.869537, 1.434631, 5.486725, 3.961716, 
    2.972137, 1.639069, 3.061722, 5.844788, 8.628647, 10.86823, 9.706238, 
    8.5737, 3.403656, 6.654694, 5.121872, 10.1315, 9.282806, 11.60521, 
    10.51796, 9.302856, 9.290878, 6.777878, 6.919785, 6.601044, 6.027084, 
    7.948181, 10.43333, 9.40834, 4.800781, 0.8473969, -1.377335, 2.21405, 
    -5.682281, -5.404678, 5.586716, 9.496094, 8.632034, 2.929688, -2.177612, 
    0.2367249, -0.6867218, -0.1234436, 4.5737, -3.969009, -4.976822, 
    -1.255203, -1.227356, -4.683594, -0.9848938, 5.194275, 5.019791, 
    9.302078, 6.530716, 2.239853, -4.172394, -3.130722, -4.684113, -6.365891, 
    -5.946609, -6.946365,
  -5.770569, -5.532547, -3.840118, -5.229172, -5.439316, -5.866669, 
    -8.009125, -8.205994, -4.801559, -3.353134, -7.93515, -13.23463, 
    -12.79166, -10.37474, -10.50781, -3.703384, -1.593491, -1.257034, 
    -2.064575, -4.594009, -6.552078, -8.717453, -5.910156, -5.12944, 
    -1.845306, 2.497925, -4.493484, -6.489578, -10.37213, -7.860413, 
    -4.063278, 3.632034, 5.160156, 6.909103, 5.722656, 7.494797, 6.436447, 
    2.235153, 2.424728, -0.3804626, 3.471619, 2.703125, 3.694534, 4.120056, 
    1.602341, 3.222916, 11.83723, 6.199478, 7.624481, 9.688278, 8.519272, 
    8.286209, 6.574219, 7.417969, 8.107803, 5.126816, 7.714844, 1.818756, 
    2.073181, 3.110672, 4.898956, 6.176041, 6.956253, 7.678116, 5.886459, 
    4.968231, 3.313538, 5.934906, 6.351822, 9.972137, 12.85859, 2.937241, 
    -1.774734, -4.764572, -6.531509, -5.501038, -2.868759, -0.2176971, 
    -0.2763062, -0.5838623, 2.145569, -3.68985, -1.327591, -2.284103, 
    -1.504684, -0.8033905, 4.449738, 7.913025, 6.255997, 4.529678, -1.251297, 
    -2.885162, -4.476303, -5.552353, -5.469269, -5.282547,
  -2.448685, -2.120041, -1.352859, -0.7492218, -2.888809, -4.316147, 
    -5.719788, -8.112503, -4.470047, -3.989578, -4.199997, -7.590897, 
    -12.01042, -8.630478, -7.805984, -6.316666, 3.998184, -0.5341187, 
    -3.162506, -1.957031, -4.051041, -3.816147, -1.422134, -7.226563, 
    -5.539841, -3.321106, -2.224228, -4.497406, -5.935677, -10.04115, 
    -14.51901, -4.283859, 4.476044, 6.895309, -0.7177124, 2.489578, 7.466141, 
    5.847137, 3.254944, 3.21199, 4.592972, 2.848175, -0.2406311, -1.271088, 
    -0.8825531, 1.625259, 0.8333282, 4.99556, 3.074738, 2.519531, 4.737488, 
    7.751572, 8.182297, 9.666412, 4.1651, 5.245316, 4.681244, 3.469536, 
    4.772919, 3.676292, 3.514061, 2.043747, 1.731262, 3.627594, 2.853134, 
    4.0401, 5.053909, 8.399734, 10.56693, 21.93021, 13.44218, -0.9351501, 
    -4.163017, -3.5737, -6.188538, -4.552597, 0.1377563, -0.3218689, 
    -1.008591, -1.484894, 1.944016, -0.07655334, 0.7510376, -2.4151, 
    -4.767441, -4.378387, -0.8502655, 4.27475, 6.11145, 5.442184, -1.494263, 
    -2.781509, -4.417709, -5.600006, -5.283325, -4.004684,
  -1.387238, -1.970566, 0.3661499, -0.2250061, -2.274475, -3.421356, 
    -1.526825, -5.794006, -5.04454, -4.077866, -3.736465, -2.473434, 
    -2.163544, -5.793488, -4.295319, -4.967972, 1.6875, 0.6231689, -3.150772, 
    -0.453125, 2.948166, 5.891403, 1.812759, -1.893997, -4.159637, -2.940628, 
    -4.341934, -10.62239, -3.843491, -2.540619, -9.933334, -5.382034, 
    5.082809, 7.680733, 3.494011, 3.760674, 4.273438, 5.24427, 6.841927, 
    3.048958, 5.136719, 3.729683, 4.92318, 2.876823, 4.138542, 4.04245, 
    1.539063, 5.246353, 4.628128, 4.87709, 4.294792, 3.769791, 4.776299, 
    3.276817, 1.156769, 0.08229065, -0.6679688, 0.1195297, 1.367966, 
    1.122131, -1.824219, 0.01328278, 3.659119, 4.539841, 4.068237, 
    -0.1059875, -0.5700531, 2.956512, 10.38333, 10.4026, 11.52708, 7.085419, 
    -2.544533, -3.495827, -4.66745, -1.355988, -3.989059, -2.673439, 
    -3.201828, -0.4312515, 0.2273483, -0.5408859, 0.5773468, 1.240883, 
    2.195053, -0.4510422, 0.02656555, 1.283592, 2.220314, 3.552605, 3.114319, 
    -0.08332825, -2.503906, -2.914322, -3.753906, -0.03593445,
  6.188553, 5.512238, 4.433853, 1.670311, 1.250778, 3.117973, 4.551826, 
    -0.4669266, 1.319008, 1.776825, 3.185936, 0.9802094, 0.9604034, 
    -0.8903656, -3.344528, -2.341667, -1.485413, 0.6552124, 1.284119, 
    0.9476471, 4.019791, -0.1289063, -3.129166, -4.870834, -2.898438, 
    2.79245, -2.726563, -8.553116, -4.704948, -0.7247391, -5.329681, 
    -5.804169, -1.729691, 1.607811, -2.260155, 1.40625, -0.4669266, 
    0.1023407, 0.04140472, 1.219536, 0.8861923, 1.970047, 0.1408844, 
    -0.7101593, 1.165108, 1.914322, 0.3700562, 1.418495, 1.336716, 5.419266, 
    2.486725, 1.647392, -0.2197952, -0.04557037, -1.59948, -0.02161407, 
    1.242455, 0.5393219, -0.9536438, -1.130989, 2.189323, 3.061195, 1.199486, 
    1.901566, 3.347122, 1.808594, -0.0171814, 0.8044281, 6.512497, 3.741669, 
    3.569794, 4.335411, 3.014328, 3.567444, -0.7354202, -4.471352, -5.683327, 
    0.4091187, -1.36042, -4.542442, -4.011459, -2.002083, 0.5500031, 
    -1.007813, -0.8817749, 0.2216187, -1.717705, -1.655212, -1.453125, 
    -2.711464, -0.5901031, 2.771614, 4.421875, 1.272919, 5.727089, 11.30391,
  10.9565, 13.49948, 11.21484, 3.822136, 2.958069, 6.518234, 2.519531, 
    1.357811, 4.595573, 5.418755, 5.814583, 3.550781, 2.174744, 1.142715, 
    -0.04895782, -6.598434, -5.424736, -1.81823, 0.1174469, -0.7302094, 
    -1.353119, -3.085938, -1.728645, -4.170578, -7.187241, -6.136459, 
    -4.050522, -4.070053, -5.000778, -6.496094, -5.801041, -8.128647, 
    -5.768486, -6.041405, -6.717705, -3.691666, 0.2489548, -8.501564, 
    -4.283333, 3.025002, 1.663025, -1.525002, 0.8179703, -0.8940125, 
    -0.6669235, -2.350784, -1.443489, -1.589325, -2.580467, -2.733849, 
    -2.482025, -0.5473938, 0.05806732, -1.533073, -1.508591, -4.1763, 
    -1.986198, -4.450523, -2.315628, -1.780212, -1.541664, 0.6010437, 
    1.867447, -0.6354218, 0.7401047, -0.7226563, 0.5231781, -3.106773, 
    -0.9164047, -1.639328, -1.454948, -3.008331, -3.457031, -4.87735, 
    -4.667969, -1.730209, -2.001305, 0.4802094, 2.28437, 2.261986, 1.664581, 
    3.999474, 3.189323, 2.379425, -2.115891, -1.129425, 2.768486, -1.702339, 
    -4.861977, -3.339058, -3.021614, -1.092972, 1.625778, 5.398438, 5.917969, 
    9.771873,
  2.055466, 3.862762, 7.672653, 7.23307, 1.722397, 2.768227, -0.1351585, 
    1.603127, 3.165886, 2.414322, 1.172134, -0.800518, -2.256775, -1.81823, 
    -2.629166, -3.506248, -4.462761, -6.322914, -5.225525, -3.142708, 
    -0.2903595, -3.081512, -3.035675, -2.864845, -3.794792, -5.455467, 
    -5.092705, -5.038284, -6.52005, -6.013802, -5.478386, -5.929955, 
    -6.889587, -8.136719, -8.946098, -4.375259, 0.5002594, -2.61068, 
    -3.24688, 0.8828125, 0.1656265, -0.360157, -1.366928, -1.284897, 
    1.060413, 0.3890648, -0.9036446, -3.184376, -3.310936, -2.616669, 
    -1.999741, -5.122395, -4.40234, -2.65937, -2.073177, -4.195053, 
    -3.271873, -4.607288, -2.044533, -0.7054749, -0.6518173, 0.9523392, 
    4.046356, 1.89896, 0.5080719, -1.148438, -1.870834, -2.145836, -3.596352, 
    -5.197136, -6.721092, -4.197922, -4.802086, -2.79427, -2.622398, 
    -1.902084, -2.560417, -4.003647, -3.218231, -0.9692726, 0.8872375, 
    2.30703, 1.438801, 0.9239616, 2.880726, 1.854687, 1.02552, 0.04713821, 
    -1.688023, -2.676048, -4.241142, -1.522133, -0.6869812, 4.054428, 
    6.326824, 4.486984,
  -2.46328, -0.0302124, -0.8395844, 1.47448, -1.35651, 0.1028633, -1.778385, 
    -4.258595, -3.012501, -1.857552, -3.154949, -6.110416, -5.689064, 
    -3.202343, -5.585155, -6.138283, -12.8849, -16.68359, -10.06198, 
    -7.826561, -7.646614, -6.589325, -6.823441, -6.362755, -3.922913, 
    -4.834381, -5.875786, -5.94635, -6.284897, -5.558594, -3.574478, 
    -4.598442, -3.482552, -3.069786, -5.510941, -2.341927, 0.0856781, 
    1.367188, -0.6458359, -2.082291, -4.19297, -2.99844, -2.747658, 
    -1.297398, 0.5104179, -0.499218, -1.190365, -2.094791, -0.7281227, 
    -0.4515648, -1.408855, -2.464584, -2.016926, -0.09843826, -0.1437492, 
    0.6312485, -0.297657, -1.297657, 0.4151039, 1.814323, -0.485157, 
    -0.3958321, 1.489582, -0.2880173, -1.809113, -1.624218, -1.099216, 
    -0.3372383, -3.669792, -5.505726, -6.880989, -6.023178, -4.857555, 
    -4.808071, -3.787502, -2.76432, -1.47448, -3.094532, -2.141148, 
    -0.09713364, -0.982811, 1.190624, 1.155991, 0.1385422, 1.933331, 
    -0.002605438, -0.5106773, -0.3088531, 0.001564026, -0.02526093, 
    -0.3562469, -0.07421875, -0.2778625, 1.290886, 3.153648, 0.1968765,
  0.9958324, 0.4341145, -0.6934891, -1.386457, -2.168488, -1.885157, 
    -2.272396, -1.390102, -3.670572, -3.682293, -3.318232, -4.891928, 
    -3.808332, -2.845831, -5.36198, -5.927864, -8.561459, -11.05755, 
    -10.26667, -9.135418, -9.929947, -6.415886, -5.494011, -4.872135, 
    -2.388542, -2.64922, -4.527863, -4.315624, -3.105209, -3.310417, 
    -2.653385, -2.858856, -1.679951, -1.339584, -3.923962, -3.097134, 
    -1.527084, 0.4046898, 0.8658867, 0.1541672, -1.259895, -0.6734352, 
    0.1458359, -1.183334, -1.660419, -1.916927, -2.25547, -0.02500153, 
    -0.007549286, -0.8468742, -0.8085938, -0.08880234, -0.607811, -2.04427, 
    -1.334896, -0.7807274, 0.6059914, 0.347393, 2.003906, 2.216667, 
    0.2734375, 1.719791, 2.308071, -0.4059906, -3.060156, -1.778908, 
    -2.030209, -3.334373, -5.528648, -5.094013, -5.162498, -5.966408, 
    -2.780991, -0.6390648, -2.140364, -4.006248, -2.529428, -2.666405, 
    -2.477341, -0.2955742, 0.3213539, -0.8994789, 0.794529, 1.523178, 
    -0.3442726, 1.134117, 1.090363, -0.6901016, -1.391926, -1.689842, 
    -0.35495, -0.6046867, -2.420052, 0.2619781, 1.283073, 0.4692707,
  2.233072, 0.03645897, -0.4752617, -0.4036465, -1.226042, -2.099739, 
    -0.9588547, -0.1033859, -1.608854, -1.752342, -1.144531, -2.115364, 
    -3.469791, -1.919792, -3.821095, -6.347918, -5.968229, -5.363281, 
    -5.7875, -5.404688, -3.329947, -2.97578, -3.393488, -3.857813, -1.646357, 
    -1.943489, -2.929169, -1.845314, -3.076305, -3.171616, -1.289845, 
    -1.202866, -1.468491, -1.572132, -1.610157, -2.200001, -2.214844, 
    -1.874741, -0.2528629, 0.5101566, -0.7625008, -0.557291, 0.2281246, 
    0.3424473, 0.3942719, 0.5187492, -0.4013023, 0.00104332, -1.063282, 
    -0.8416672, 0.04036522, 0.8151054, 0.3554688, -0.198698, -0.1658859, 
    -0.6463528, 0.6744785, 1.164583, 0.916666, 0.4598961, 0.6442719, 
    0.4937496, 0.0901041, 0.276042, -0.3531246, -1.951302, -3.004948, 
    -2.120314, -2.988802, -2.91198, -2.159115, -1.653387, -1.271355, 
    -2.35651, -3.428646, -2.813021, -2.007813, -2.232553, -1.163801, 
    0.3059902, 2.367447, 1.31875, 2.245832, 1.871094, 0.4166679, 0.3854179, 
    1.202084, 0.5731754, -0.004688263, -0.1132813, -1.040886, -1.830469, 
    -1.062759, -1.077604, -1.584896, 0.7661457,
  0.1531248, 0.2226563, -0.9507809, -1.722136, -1.600521, -1.012239, 
    -0.296093, -0.5289059, -1.528646, -1.696355, -1.835677, -1.998697, 
    -2.180469, -2.460418, -2.011458, -2.609114, -2.346615, -2.439583, 
    -2.386459, -1.71276, -1.142189, -1.46875, -1.286459, -0.7062492, 
    -0.4932289, 0.04583359, -0.4593754, -0.4182281, -0.5372391, -1.101824, 
    -1.53047, -1.166147, -1.391146, -1.144011, -1.563282, -1.788801, 
    -1.282291, -1.915104, -0.3195305, -0.7184896, -0.3747396, -0.656251, 
    -0.6744795, -0.2278652, 0.3098965, -0.2229166, -0.6617184, 0.02838516, 
    0.05182362, 0.4986973, 0.3231773, -0.3830738, -0.244791, 0.09062481, 
    0.3734379, 0.008853912, 0.2234383, 0.3289061, 0.8343744, 1.275261, 
    0.9203129, -0.109375, 0.01822948, 0.9661465, 0.7539063, -1.234375, 
    -1.105207, -1.311979, -0.9919281, -0.5429688, -0.2361975, -1.63776, 
    -1.989583, -2.496875, -1.964323, -1.823698, -1.539063, -1.773958, 
    -1.726563, -0.5872402, 0.8682289, 1.797657, 1.795833, 0.817709, 
    0.2458334, 0.5835943, 1.046615, 0.776042, 0.6903648, 1.218229, 0.7703123, 
    0.1786461, 0.02682304, -0.6742182, -1.486458, -1.14375,
  -0.2263021, -0.2507815, -0.2328129, -0.2867188, -0.5088539, -0.2104168, 
    0.1429691, -0.08984375, -0.3153644, -0.3268228, 0.1604166, -0.4124999, 
    -0.794271, -0.9518228, -0.6229167, -0.6302085, -0.953125, -1.354948, 
    -1.345313, -1.503386, -1.699739, -1.153125, -0.6328125, -0.2830725, 
    -0.1367188, -0.200521, -0.1114583, -0.2627602, -0.1653652, -0.4601564, 
    -0.9466143, -1.058854, -1.040365, -1.310156, -1.592968, -1.716928, 
    -1.404427, -1.257552, -0.3468752, -0.01484394, 0.2158852, -0.4388027, 
    -0.796875, -0.5703125, -0.04635382, 0.4968753, 0.2315102, 0.06145859, 
    0.1526041, 0.3286457, 0.3125, 0.3994799, 0.8877602, 1.001302, 
    -0.09557295, -0.0546875, -0.2476559, -0.2028642, 0.2518229, 0.04140615, 
    -0.2671876, -0.2437501, -0.2104168, -0.1088543, -0.2776036, -0.05234337, 
    0.0817709, -0.09479141, -0.05755234, -0.4005208, -0.8325524, -1.265364, 
    -1.33776, -1.058333, -1.503125, -1.908593, -1.182032, -1.115625, 
    -1.108854, -0.7401042, -0.1395836, 0.4132814, 0.2598958, 0.1994791, 
    -0.04296875, 0.1726561, 0.1312499, -0.08359432, 0.2210937, 0.6333332, 
    0.3901043, -0.3390622, -0.3669271, -0.09505177, -0.5122395, -0.5052085,
  -0.05989599, -0.2445312, -0.3111979, -0.2601563, -0.1513021, 0.03723955, 
    0.006510496, -0.08411479, -0.3007811, -0.3893229, -0.2651043, -0.1875001, 
    -0.248698, -0.2778646, -0.3302084, -0.4919271, -0.4591146, -0.4153645, 
    -0.335677, -0.2955728, -0.3388021, -0.340625, -0.3502603, -0.3200521, 
    -0.3041666, -0.2447917, -0.1604167, -0.0617187, -0.06640625, -0.1914063, 
    -0.2640624, -0.463021, -0.3372397, -0.4710937, -0.5979168, -0.7718749, 
    -0.5710936, -0.5273435, -0.4885418, -0.4908855, -0.5783854, -0.5856771, 
    -0.6098957, -0.6158855, -0.58125, -0.46875, -0.1742188, 0.0005209446, 
    0.04791665, 0.08411455, -0.001822948, -0.1591146, -0.2427084, -0.5515623, 
    -0.7291667, -0.6299479, -0.3164063, -0.1367188, -0.03593743, -0.0979166, 
    -0.1078125, -0.1864583, -0.1302083, -0.008072853, -0.04140615, 0.015625, 
    -0.2101562, -0.1807292, -0.06354165, -0.2111979, -0.3768229, -0.8203125, 
    -1.030469, -1.202865, -1.146354, -0.8528647, -0.6781249, -0.9169272, 
    -1.053906, -0.6520832, -0.4953125, -0.4132814, -0.4242189, -0.4200521, 
    -0.1231771, 0.07500005, 0.1903646, 0.2119792, 0.1679688, 0.2190104, 
    0.1369791, -0.08333325, 0.0270834, 0.201823, 0.1697917, 0.03072906,
  0.001041681, -0.01406249, -0.01927084, -0.05078124, -0.04140624, 
    -0.002343744, 0.002083331, -0.02005209, -0.03567708, -0.05416667, 
    -0.05260417, -0.03229167, -0.02890626, -0.03411458, -0.03541668, 
    -0.03333333, -0.02473958, -0.04348958, -0.05026042, -0.08697917, 
    -0.07187502, -0.03880207, -0.02005209, -0.04374999, -0.03437501, 
    -0.02187499, -0.01901041, -0.04739583, -0.07161459, -0.1122396, 
    -0.1049479, -0.09739584, -0.1166667, -0.1184896, -0.1088542, -0.08203125, 
    -0.07447916, -0.09791669, -0.09713542, -0.1109375, -0.06927085, 
    -0.06276041, -0.05104166, -0.06536457, -0.07604167, -0.07057291, 
    -0.06276041, -0.07343748, -0.09869793, -0.1140625, -0.1171875, -0.1625, 
    -0.1223958, -0.1114583, -0.08307293, -0.08802083, -0.09713542, 
    -0.08906251, -0.06354165, -0.04401043, -0.02812502, -0.01640627, 
    -0.01406249, -0.0127604, -0.004166663, 0.02291664, 0.001041651, 
    -0.01692709, -0.0341146, -0.008333325, -0.007552058, -0.03932291, 
    -0.07447916, -0.07838541, -0.07682294, -0.04609373, -0.06588542, 
    -0.1247396, -0.1723958, -0.1544271, -0.1744792, -0.1677083, -0.1481771, 
    -0.1481771, -0.1018229, -0.06197917, -0.04062501, -0.02526042, 0.0078125, 
    0.02083334, 0.03203124, 0.02317709, 0.03463539, 0.008854151, -0.01640624, 
    -0.02135417,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0,
  0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0 ;
}
