netcdf CGMR_SRA1B_1_vas-change_2070-2099 {
dimensions:
	time = 12 ;
	latitude = 48 ;
	longitude = 96 ;
	bounds = 2 ;
Data:
 northward_wind_anomaly =
  -0.127372, -0.1206014, -0.1133585, -0.1065063, -0.1008584, -0.09682202, 
    -0.09457612, -0.09394145, -0.09340429, -0.09355044, -0.09504771, 
    -0.09674048, -0.09799385, -0.09918189, -0.09804273, -0.09612203, 
    -0.09384334, -0.09193933, -0.09125578, -0.09250915, -0.09652922, 
    -0.1025839, -0.1119915, -0.1238242, -0.1386517, -0.1548626, -0.1745405, 
    -0.1974566, -0.2215781, -0.2475543, -0.2759724, -0.3065388, -0.336731, 
    -0.366744, -0.3967893, -0.4246867, -0.4479132, -0.4667282, -0.4796515, 
    -0.4883752, -0.4930143, -0.4953413, -0.4935348, -0.4875774, -0.4807739, 
    -0.4716756, -0.4576132, -0.439384, -0.4168251, -0.3874631, -0.3614049, 
    -0.3183064, -0.297701, -0.27677, -0.2271607, -0.1996378, -0.1475058, 
    -0.1063602, -0.06915301, -0.0340293, -0.01148701, 0.04905987, 0.08753645, 
    0.1160032, 0.145235, 0.1721393, 0.1950885, 0.2127155, 0.229317, 
    0.2424355, 0.2514036, 0.2550331, 0.2499063, 0.2190631, 0.2270384, 
    0.2187052, 0.1933144, 0.169942, 0.1605996, 0.1380736, 0.1123411, 
    0.08597404, 0.05924878, 0.03314199, 0.007979229, -0.01716724, 
    -0.03990501, -0.06060809, -0.07891858, -0.09416926, -0.107564, 
    -0.1174599, -0.1253541, -0.1302533, -0.131978, -0.1308386,
  -0.2141399, -0.1825645, -0.1415486, -0.08804941, -0.03328061, 0.01849413, 
    0.06221151, 0.09593511, 0.1197146, 0.1276571, 0.1148803, 0.08971739, 
    0.05648184, 0.02218822, -0.01039642, -0.03948173, -0.06428638, 
    -0.08212492, -0.09333912, -0.09853119, -0.09854746, -0.0968222, 
    -0.09193938, -0.08464772, -0.07733977, -0.06833923, -0.06322861, 
    -0.07234323, -0.09039271, -0.1258259, -0.1704221, -0.2185669, -0.2574341, 
    -0.2841756, -0.2955532, -0.2957001, -0.2844372, -0.2716932, -0.2649217, 
    -0.2638636, -0.2714317, -0.2725055, -0.2624307, -0.2642701, -0.2765906, 
    -0.2624958, -0.2940385, -0.300891, -0.3068482, -0.3031372, -0.2992961, 
    -0.3104128, -0.2856243, -0.2663698, -0.194511, -0.1959921, -0.1380331, 
    -0.08469653, -0.0428347, 0.01370829, 0.07472718, 0.1238972, 0.1583862, 
    0.1745481, 0.1914752, 0.2211465, 0.2399616, 0.2522175, 0.2777058, 
    0.3099324, 0.3440306, 0.3535032, 0.3517944, 0.3454145, 0.2940632, 
    0.2431195, 0.1929568, 0.1541384, 0.1027546, 0.0756712, 0.05438215, 
    0.02663156, 0.01265046, -0.02382415, -0.05338144, -0.09050712, 
    -0.1279909, -0.159013, -0.1850547, -0.205367, -0.2225542, -0.230204, 
    -0.2377889, -0.2489705, -0.2507606, -0.2369914,
  -0.4665649, -0.3981729, -0.2935345, -0.1701131, -0.0470171, 0.0733602, 
    0.1831746, 0.2472207, 0.2612833, 0.2594603, 0.2562702, 0.2573119, 
    0.2477579, 0.2265338, 0.1994668, 0.1814004, 0.1628621, 0.133728, 
    0.09294017, 0.03851309, -0.01659769, -0.05619729, -0.07419848, 
    -0.05950135, -0.02491474, 0.01095775, 0.03584382, 0.0510945, 0.04881579, 
    0.01738703, -0.04187417, -0.127063, -0.2162716, -0.2884884, -0.3299601, 
    -0.3372843, -0.3087687, -0.2751751, -0.2421346, -0.2149374, -0.2153115, 
    -0.1831822, -0.1305618, -0.1328247, -0.1262164, -0.1160765, -0.105839, 
    -0.1257609, -0.1591108, -0.1898073, -0.2123171, -0.2343385, -0.243746, 
    -0.2308554, -0.1819786, -0.09693617, -0.0084759, 0.05553794, 0.1249229, 
    0.1967815, 0.2529336, 0.2815796, 0.2822306, 0.2634158, 0.2531617, 
    0.2464719, 0.2716511, 0.311267, 0.3603554, 0.3789102, 0.3636436, 
    0.3213745, 0.2541218, 0.1765342, 0.1134646, 0.08192134, 0.07168376, 
    0.09617937, 0.1153197, 0.1340533, 0.1408567, 0.1312377, 0.1163288, 
    0.09194733, 0.05203849, 0.0107787, -0.04057229, -0.09713155, -0.1587852, 
    -0.205416, -0.2905395, -0.3397094, -0.4007608, -0.4647907, -0.5049114, 
    -0.504781,
  -0.1218547, -0.02187085, 0.09012425, 0.2081907, 0.3132527, 0.3901895, 
    0.4451863, 0.4683959, 0.4307495, 0.3484417, 0.2452679, 0.142224, 
    0.07632226, 0.04277736, 0.0472858, 0.07067454, 0.07047927, 0.04300559, 
    -0.007645845, -0.05388603, -0.09477141, -0.1446897, -0.176363, -0.162528, 
    -0.1025677, -0.02330339, 0.06903067, 0.1402221, 0.1569863, 0.1229695, 
    0.05034578, -0.03443623, -0.1018516, -0.1471803, -0.1539024, -0.1163861, 
    -0.0618124, -0.04534078, -0.08371973, -0.1524212, -0.2218053, -0.2758093, 
    -0.2028606, -0.1012816, -0.02289629, 0.005603075, -0.04875875, -0.172245, 
    -0.2299441, -0.3278282, -0.3624147, -0.3880494, -0.3543417, -0.269446, 
    -0.1788372, -0.07869083, -0.004341841, 0.1066122, 0.1368366, 0.1186888, 
    0.0907917, 0.02446684, -0.03326426, -0.0551067, -0.04906827, -0.02082944, 
    0.02438533, 0.05988371, 0.0751996, 0.05308056, -0.01052666, -0.09276938, 
    -0.1744425, -0.2191855, -0.2198853, -0.1580685, -0.07502854, 0.03748775, 
    0.1537636, 0.2207233, 0.2233601, 0.2044148, 0.1451863, 0.08937572, 
    0.02052806, -0.04991466, -0.1126588, -0.184778, -0.2398562, -0.2564577, 
    -0.2854291, -0.3119752, -0.3015097, -0.2872028, -0.2513793, -0.1845171,
  0.05439851, 0.1317748, 0.2071654, 0.249597, 0.2398802, 0.2222695, 
    0.1403849, 0.04313588, -0.05828047, -0.1504681, -0.2064247, -0.2060997, 
    -0.1662883, -0.1268189, -0.1038861, -0.1153768, -0.1334105, -0.169934, 
    -0.1662395, -0.1205198, -0.06527923, -0.008573651, 0.05065536, 0.134656, 
    0.2127479, 0.2675984, 0.3108602, 0.3306195, 0.2933633, 0.1967, 
    0.06850994, -0.03806579, -0.1092572, -0.1360314, -0.09602451, 
    -0.03282475, -0.001964808, -0.04221606, -0.1601033, -0.3044069, 
    -0.4072387, -0.3940878, -0.2469361, -0.03433847, 0.1202679, 0.1854858, 
    0.09014106, -0.0445106, -0.1727498, -0.2290977, -0.2497193, -0.2340129, 
    -0.1609173, -0.06308196, -0.01965748, -0.0432903, -0.06881113, 
    -0.0898886, -0.09075124, -0.08287363, -0.1130168, -0.2059531, -0.298287, 
    -0.381604, -0.4105592, -0.3906701, -0.3273237, -0.2333946, -0.1610473, 
    -0.1193973, -0.05920815, -0.079, -0.08127868, -0.1144493, -0.1368776, 
    -0.1146445, -0.07397065, 0.01042064, 0.08198639, 0.1425984, 0.09839265, 
    0.01045318, -0.04530852, -0.03809823, -0.0003866553, 0.03750397, 
    0.0537963, 0.01382233, -0.0609498, -0.1351523, -0.1976848, -0.1390748, 
    -0.1431763, -0.124817, -0.09094656, -0.0246054,
  -0.06039643, 0.01248771, 0.03312573, 0.007425845, -0.02836525, -0.07948828, 
    -0.1201621, -0.08572209, -0.08328044, -0.1090454, -0.1055625, -0.1294557, 
    -0.1392701, -0.09062102, -0.07846284, -0.1476682, -0.3002396, -0.3909791, 
    -0.4369588, -0.3311645, -0.1421836, -0.00829681, 0.09290762, 0.1354206, 
    0.1622924, 0.1503947, 0.1087122, 0.02770615, -0.07873917, -0.1818806, 
    -0.2563925, -0.2882935, -0.3226521, -0.3556112, -0.3863075, -0.3815062, 
    -0.3710079, -0.3707962, -0.4486935, -0.4939899, -0.4915974, -0.3689735, 
    -0.1387649, 0.09198046, 0.1725953, 0.1508503, -0.02135015, -0.1043251, 
    -0.1154746, -0.05190033, 0.06043692, 0.2207071, 0.2668822, 0.2012735, 
    0.09780669, -0.09394133, -0.2355755, -0.2985312, -0.2691692, -0.257483, 
    -0.3147421, -0.3676393, -0.450403, -0.5101361, -0.5108034, -0.4567508, 
    -0.2970665, -0.1523889, -0.006587863, 0.1885293, 0.2175494, 0.2091022, 
    0.1528848, 0.07842195, 0.01611725, -0.04761972, -0.06257741, -0.1112591, 
    0.03044017, 0.04702546, 0.02226961, -0.04706635, -0.06710215, 
    -0.06112884, -0.01763926, -0.01995045, -0.03479421, -0.1079225, 
    -0.2106243, -0.2603964, -0.2449504, -0.1766236, -0.1144167, -0.1001425, 
    -0.1309531, -0.1162884,
  -0.1947877, -0.1366334, -0.08671486, -0.06982017, -0.01890862, 0.02018631, 
    0.02340901, -0.003837228, -0.06304932, -0.1676067, -0.2993287, -0.412789, 
    -0.476819, -0.4861938, -0.4328735, -0.3850706, -0.3357217, -0.2795043, 
    -0.2268186, -0.1366981, -0.08209252, -0.05286068, 0.00181067, 
    -0.005513728, -0.0399375, -0.0180788, 0.01362693, 0.02301848, 
    -0.01534414, -0.09726167, -0.159013, -0.1592246, -0.1518191, -0.1093061, 
    -0.2825643, -0.4458455, -0.4004028, -0.2952267, -0.4249793, -0.5342405, 
    -0.492704, -0.2758095, 0.0678103, 0.3785354, 0.4610716, 0.2831583, 
    0.1055377, 0.07254621, 0.1303751, 0.1797891, 0.1718464, 0.03651112, 
    -0.1312135, -0.2556275, -0.356246, -0.412024, -0.4699179, -0.6084107, 
    -0.7193808, -0.8128867, -0.8925905, -0.9794719, -1.096953, -1.219625, 
    -1.212675, -1.032581, -0.7258427, -0.4255332, -0.1630006, -0.03528261, 
    -0.01394463, -0.03358984, -0.07683533, -0.05740166, 0.007507235, 
    0.03444408, 0.09647207, 0.09858796, 0.07209057, 0.03789461, -0.056539, 
    -0.03482676, 0.1130574, 0.2752156, 0.3810587, 0.2859089, 0.1269245, 
    -0.02779555, -0.182776, -0.270276, -0.2447064, -0.1084108, 0.04368877, 
    0.0473997, -0.02533787, -0.1471315,
  -0.5909791, -0.5268191, -0.4802045, -0.458411, -0.5011518, -0.5719852, 
    -0.6573856, -0.7950158, -0.8411909, -0.8597131, -0.9470013, -1.095894, 
    -1.168697, -1.162692, -1.12179, -1.007531, -0.8431597, -0.5740356, 
    -0.3415002, -0.204163, -0.1492474, -0.07167584, 0.01868874, 0.08361387, 
    0.1274615, 0.1495808, 0.1882689, 0.2234577, 0.1405313, -0.02359641, 
    -0.1458619, -0.2310996, -0.3243288, -0.5277141, -0.7841268, -0.9449015, 
    -0.9587687, -0.8741173, -0.7534955, -0.6355593, -0.444674, -0.1665163, 
    0.1313515, 0.3111042, 0.2300006, 0.08166088, -0.003381443, 0.03044017, 
    0.05641672, 0.0006224513, -0.194983, -0.4110312, -0.6450319, -0.7424601, 
    -0.7889772, -0.757304, -0.8298789, -1.055839, -1.368079, -1.634387, 
    -1.730237, -1.715833, -1.725045, -1.821171, -1.824508, -1.544121, 
    -1.056148, -0.5907837, -0.3044396, -0.2619752, -0.2581667, -0.2635866, 
    -0.2315065, -0.1628216, -0.07979746, -0.02595632, -0.06635347, 
    -0.1562786, -0.2240031, -0.2456178, -0.2229941, -0.09114186, 0.1433633, 
    0.3626179, 0.3915078, 0.2447631, 0.0989134, -0.03819603, -0.2318483, 
    -0.5082318, -0.6477662, -0.5346152, -0.3970826, -0.374931, -0.4642048, 
    -0.5701782,
  -1.052177, -0.9565878, -0.8221477, -0.8149537, -0.9485473, -1.080432, 
    -1.201152, -1.231344, -1.283639, -1.379097, -1.561552, -1.655139, 
    -1.632597, -1.551559, -1.434322, -1.264026, -1.016532, -0.7973105, 
    -0.6880168, -0.685787, -0.6549603, -0.4938599, -0.3244589, -0.1564251, 
    0.01942129, 0.1215046, 0.02666412, -0.1779095, -0.3915977, -0.5208131, 
    -0.6303183, -0.7256471, -0.8746217, -1.038456, -1.158964, -1.209908, 
    -1.194723, -1.197115, -1.133997, -0.9917278, -0.8465618, -0.6725546, 
    -0.6141399, -0.5853964, -0.6089153, -0.6007122, -0.4750611, -0.3193483, 
    -0.3537722, -0.3961225, -0.470878, -0.6222776, -0.7958617, -0.9055134, 
    -1.020552, -1.103121, -1.310006, -1.592639, -1.902258, -2.135869, 
    -2.222099, -2.221627, -2.173483, -2.116451, -1.926933, -1.51204, 
    -1.007402, -0.5810344, -0.3864218, -0.3291139, -0.2293417, -0.1406537, 
    -0.1631633, -0.1676882, -0.06687438, -0.05738544, -0.22594, -0.4331666, 
    -0.3982383, -0.2410768, -0.1917603, -0.2744752, -0.2086223, -0.05992441, 
    0.009362698, -0.06243092, -0.1488404, -0.3033815, -0.6722943, -1.10636, 
    -1.353642, -1.267086, -1.064205, -0.9739543, -1.006148, -1.060038,
  -1.30343, -1.224427, -1.22096, -1.312203, -1.460152, -1.505611, -1.42205, 
    -1.331181, -1.468453, -1.732353, -1.813815, -1.730286, -1.644902, 
    -1.546204, -1.439433, -1.276347, -1.005465, -0.802763, -0.8585244, 
    -0.9253213, -0.831197, -0.648238, -0.5856402, -0.5424926, -0.4072715, 
    -0.4719688, -0.7503378, -0.9882285, -1.068144, -1.028056, -1.054065, 
    -1.186145, -1.329439, -1.401786, -1.32703, -1.251509, -1.338391, 
    -1.511633, -1.539172, -1.427258, -1.361845, -1.441142, -1.429635, 
    -1.365507, -1.186894, -0.976005, -0.8378052, -0.69884, -0.6215291, 
    -0.525175, -0.4771281, -0.553707, -0.6577595, -0.8288047, -1.041272, 
    -1.277258, -1.583574, -1.880595, -2.024296, -2.098238, -2.214742, 
    -2.308915, -2.203642, -1.890247, -1.507125, -1.251884, -1.020699, 
    -0.7586875, -0.4941855, -0.3117636, -0.2269003, -0.267216, -0.3292439, 
    -0.2708781, -0.1084105, -0.1330528, -0.4450157, -0.6632121, -0.5413858, 
    -0.3561646, -0.4977337, -0.7727174, -0.800289, -0.7018189, -0.6666139, 
    -0.6440879, -0.5983847, -0.7519817, -1.178398, -1.460673, -1.47013, 
    -1.392346, -1.362154, -1.353902, -1.348238, -1.355986,
  -1.177746, -1.130204, -1.229781, -1.41051, -1.488245, -1.447473, -1.429667, 
    -1.409566, -1.509957, -1.618876, -1.572587, -1.428251, -1.313391, 
    -1.255367, -1.186194, -1.061991, -0.8559368, -0.6201458, -0.5921998, 
    -0.6568317, -0.5655069, -0.4550741, -0.525419, -0.6344526, -0.6984985, 
    -0.8624471, -1.075273, -1.145699, -1.149117, -1.184094, -1.179944, 
    -1.1283, -1.058069, -1.06414, -1.139335, -1.296741, -1.469348, -1.56982, 
    -1.570683, -1.514953, -1.522571, -1.660217, -1.824784, -1.821887, 
    -1.583443, -1.254146, -0.9456501, -0.7317016, -0.5738406, -0.4436324, 
    -0.3747029, -0.369169, -0.3338501, -0.523108, -0.9218873, -1.358085, 
    -1.659713, -1.845439, -1.970895, -2.067688, -2.176656, -2.158166, 
    -1.849166, -1.375159, -1.052339, -0.9118282, -0.7409787, -0.4954058, 
    -0.2134726, -0.07641196, -0.112561, -0.1344361, -0.04042578, 0.1092813, 
    0.1300983, -0.1646771, -0.5854292, -0.5609663, -0.2804811, -0.2676556, 
    -0.6526165, -1.024752, -1.126412, -1.121545, -1.031116, -0.8636679, 
    -0.7336875, -0.8397906, -1.092753, -1.159045, -1.123466, -1.252291, 
    -1.43595, -1.464449, -1.391402, -1.286861,
  -0.6802368, -0.7800415, -0.8824992, -0.9770956, -0.9850057, -0.9812294, 
    -0.9788535, -0.9322224, -0.8732053, -0.8170205, -0.6989055, -0.595422, 
    -0.5416625, -0.4753861, -0.3746214, -0.2796671, -0.2259235, -0.1725221, 
    -0.1469362, -0.1944947, -0.2781534, -0.3804972, -0.5007281, -0.5576291, 
    -0.6046669, -0.702014, -0.7588825, -0.7864866, -0.8636842, -0.8738403, 
    -0.726721, -0.5837684, -0.5756795, -0.6308391, -0.7559204, -0.9134886, 
    -1.003397, -1.086682, -1.237854, -1.370471, -1.525728, -1.691826, 
    -1.76344, -1.724964, -1.487561, -1.012235, -0.5942013, -0.3343387, 
    -0.1676068, 0.02244902, 0.1645062, 0.2228072, 0.1024783, -0.2710087, 
    -0.8436158, -1.266777, -1.412447, -1.499199, -1.6811, -1.851103, 
    -1.836601, -1.589498, -1.189254, -0.8732706, -0.7443318, -0.6151001, 
    -0.4128375, -0.1295366, 0.11449, 0.2928269, 0.4296267, 0.5583048, 
    0.6333699, 0.6288128, 0.491101, 0.2092164, -0.04721284, -0.06830645, 
    -0.01679254, -0.2987754, -0.6610472, -0.7991496, -0.8977172, -0.9174111, 
    -0.647652, -0.3031696, -0.2287391, -0.4077759, -0.5863078, -0.6127726, 
    -0.7262166, -0.8936808, -0.9169068, -0.8431926, -0.749475, -0.6602662,
  -0.1747682, -0.2415648, -0.1933224, -0.2548623, -0.3031857, -0.2759725, 
    -0.2064573, -0.07906497, 0.00078547, 0.06336701, 0.0950886, 0.03726006, 
    -0.006945372, -0.04429889, -0.03261304, 0.02995205, 0.03491616, 
    0.02736402, 0.03130293, -0.04325771, -0.1151326, -0.1359823, -0.1695597, 
    -0.2367799, -0.3346801, -0.4107218, -0.4185343, -0.3974078, -0.2827919, 
    -0.07781172, 0.1024942, 0.1582401, 0.1021693, 0.06545043, -0.02076387, 
    -0.1829872, -0.3040161, -0.4906373, -0.5784304, -0.5444943, -0.8717407, 
    -1.214937, -1.106279, -0.9826295, -0.9201617, -0.5236287, -0.1438923, 
    0.09417748, 0.3074098, 0.6022503, 0.8109906, 0.6681843, 0.2421429, 
    -0.1489871, -0.3939252, -0.5625613, -0.6926069, -0.8928671, -1.174101, 
    -1.283769, -1.120064, -0.8266238, -0.537138, -0.3216758, -0.1938598, 
    -0.04482007, 0.2860394, 0.5770226, 0.7881067, 0.9741743, 1.037993, 
    1.004318, 1.00212, 0.8882532, 0.7465374, 0.7312216, 0.7168664, 0.5701214, 
    0.3165892, -0.2129518, -0.6045859, -0.481604, -0.2852825, -0.1864706, 
    -0.02926052, 0.01388752, -0.09635007, -0.2157184, -0.2291789, -0.1401162, 
    -0.1517699, -0.1485469, -0.02470255, -0.05302334, -0.09569883, -0.05066323,
  0.2243209, 0.207068, 0.2231815, 0.1929562, 0.3168983, 0.3695678, 0.3593301, 
    0.4578815, 0.3777872, 0.1268268, -0.1130493, -0.2700968, -0.2025836, 
    -0.03594947, 0.08613753, 0.1847372, 0.2036173, 0.2529502, 0.3578491, 
    0.3843789, 0.3466187, 0.3026083, 0.1980672, 0.07368565, 0.01691484, 
    0.1339073, 0.2969282, 0.488204, 0.807426, 0.9687216, 0.9243203, 0.905717, 
    0.7960815, 0.62087, 0.4548055, 0.3307823, 0.3472369, 0.4317096, 
    0.6331908, 0.5530475, -0.2873333, -1.019153, -0.7847286, -0.5515418, 
    -0.4776654, 0.05067134, 0.457345, 0.5654669, 0.7738488, 0.9482787, 
    0.948751, 0.7366905, 0.410697, 0.205261, 0.1347857, -0.03694272, 
    -0.2617962, -0.5361617, -0.6968061, -0.657076, -0.4568158, -0.225468, 
    -0.01483989, 0.1288617, 0.2193401, 0.4086633, 0.7103887, 0.8833541, 
    0.9339232, 1.041671, 1.069373, 1.064083, 1.104122, 0.974955, 0.7515827, 
    0.868445, 1.040906, 0.6369182, 0.1196166, -0.4544231, -0.5418417, 
    -0.1840944, 0.0664264, 0.1666217, 0.1747437, 0.02142334, -0.1052531, 
    -0.07821834, -0.07885313, 0.07031655, 0.2761924, 0.2756553, 0.3464558, 
    0.3537474, 0.3021526, 0.3091512,
  0.4735065, 0.4774455, 0.619877, 0.813985, 1.073376, 1.035307, 0.8521528, 
    0.5353559, -0.2095499, -0.7330365, -0.4252723, 0.1504925, 0.4273969, 
    0.4164916, 0.3427613, 0.4353559, 0.6117067, 0.7221236, 0.8225467, 
    0.8658085, 0.7566452, 0.6082892, 0.5575564, 0.5532755, 0.5844768, 
    0.7545936, 1.00059, 1.165743, 1.309753, 1.505685, 1.665531, 1.380131, 
    0.8109579, 0.5714723, 0.7189329, 0.8848022, 0.9797894, 1.146358, 
    1.093266, 0.6301146, -0.4031862, -1.057841, -0.8155069, -0.4705036, 
    -0.1599729, 0.4582722, 0.8341346, 0.8423055, 1.026811, 1.155815, 
    1.083858, 0.9805056, 0.8134156, 0.578406, 0.3534871, 0.1973996, 
    0.03962004, -0.1661904, -0.2384233, -0.1678345, -0.0964638, 
    -0.0008420944, 0.1898482, 0.2619669, 0.3378296, 0.5526897, 0.7676147, 
    0.8274782, 0.7985066, 0.8750363, 0.9891314, 0.9829953, 0.8592813, 
    0.7659222, 0.6817588, 0.8474979, 0.7873411, 0.2677937, -0.3712363, 
    -0.4912559, -0.04989837, 0.315629, 0.3254922, 0.06317127, -0.188912, 
    -0.4513795, -0.6525999, -0.4731894, -0.1652954, 0.1429079, 0.4900599, 
    0.4951539, 0.4958537, 0.6049032, 0.5722377, 0.5549523,
  0.4596719, 0.553894, 0.8323932, 1.141883, 1.079594, 0.8597202, 0.3957398, 
    -0.09820557, -0.5701783, -0.5429971, 0.1760456, 0.6357136, 0.4161173, 
    0.05404043, 0.05706769, 0.3984575, 0.7544799, 0.9776894, 1.031954, 
    1.044031, 0.9594604, 0.898409, 0.9229695, 0.9105834, 0.8833047, 
    0.9586303, 1.185991, 1.340173, 1.45168, 2.072237, 2.23407, 1.24421, 
    0.4559939, 0.7375041, 0.9776735, 0.9856976, 1.014604, 0.9178097, 
    0.5389692, -0.1924765, -0.7611448, -0.6194131, -0.112577, 0.2735877, 
    0.476957, 0.7891967, 1.022367, 1.132556, 1.366345, 1.425557, 1.247058, 
    1.04172, 0.8174193, 0.5968464, 0.4243204, 0.1779825, 0.02239981, 
    -0.1037721, -0.1480592, -0.03308535, 0.04201239, 0.0991087, 0.1889686, 
    0.2534382, 0.4397986, 0.6108761, 0.7110229, 0.7701211, 0.7636433, 
    0.7242715, 0.7851927, 0.8972045, 0.791801, 0.7175331, 0.6083207, 
    0.3670292, -0.07149601, -0.181376, 0.05814183, 0.2827187, 0.2496459, 
    0.04731843, -0.05017507, -0.07289642, -0.6463011, -0.8446898, -0.5025673, 
    0.03726029, 0.494308, 0.5461469, 0.5929897, 0.5932333, 0.5583378, 
    0.548816, 0.52253, 0.5368855,
  0.4536335, 0.497139, 0.4511747, 0.4490433, 0.1267457, -0.4381957, 
    -1.109062, -0.7648884, 0.006742358, 0.4743041, 0.8391644, 0.8780313, 
    0.06846082, -0.7377076, -0.5205687, 0.3157916, 0.807149, 1.032849, 
    1.041247, 0.9168497, 0.8426797, 0.7951699, 0.7127156, 0.6292686, 
    0.667973, 0.7623086, 0.9553428, 1.097366, 1.300214, 1.783125, 1.039327, 
    -0.09680581, 0.02620828, 0.7176797, 0.6835814, 0.715385, 0.8027706, 
    0.6363157, 0.06050229, -0.6880332, -0.3464476, 0.8453002, 1.334867, 
    1.240792, 1.079773, 1.004269, 1.019324, 1.072302, 1.168803, 1.128438, 
    0.8288126, 0.6226764, 0.4536822, 0.2618365, 0.1247597, -0.03160417, 
    -0.0590944, -0.02611907, -0.1015585, -0.09078379, 0.01473385, 0.07002352, 
    0.1698119, 0.3434773, 0.5865274, 0.790808, 0.8220417, 0.8020222, 
    0.8366739, 0.8090208, 0.7259808, 0.7558311, 0.6821332, 0.461463, 
    0.2289262, 0.1886759, -0.101932, -0.04763579, 0.2487669, -0.05435807, 
    -0.4274212, -0.3679647, -0.1280235, -0.1034303, -0.7471478, -0.9779416, 
    -0.1311646, 0.4962606, 0.5472212, 0.4250858, 0.3817589, 0.388692, 
    0.4171101, 0.4112833, 0.4590535, 0.4883015,
  0.1772985, 0.04316711, -0.2830038, -0.3765249, -0.5921841, -0.9905072, 
    -0.9369101, -0.1456342, 0.3474975, 0.3892784, 0.8450075, 0.7802451, 
    -0.1785276, -1.071985, -0.8618938, 0.3406453, 0.9946166, 1.100346, 
    0.9955118, 0.7870807, 0.7590863, 0.6592164, 0.5518109, 0.5269735, 
    0.5548055, 0.6164749, 0.7164426, 0.5519571, 0.4586959, 0.373148, 
    -0.618566, -0.7007606, 0.005684301, 0.4191933, 0.3523967, 0.5610553, 
    0.6197143, 0.106401, -0.5003216, -0.5067992, 0.8216836, 1.943396, 
    1.684428, 1.108777, 0.8228071, 0.6985555, 0.6441121, 0.8394899, 
    0.7505251, 0.5434124, 0.3755252, 0.1355183, 0.0297401, -0.003593087, 
    0.05198944, 0.118233, 0.06681705, -0.04312754, -0.1071412, -0.03699146, 
    0.2780964, 0.5183308, 0.7013386, 0.8487671, 0.9112344, 0.984086, 
    0.8797403, 0.7655963, 0.7394574, 0.6897992, 0.6020715, 0.4719119, 
    0.5050817, 0.4262071, 0.3175492, 0.3903689, 0.0366888, 0.01486397, 
    0.2127156, -0.267151, -0.5705689, -0.1995729, 0.02132559, -0.09801035, 
    -0.4108197, -0.4853148, 0.255033, 0.6955123, 0.5356162, 0.3945515, 
    0.2580931, 0.2307494, 0.3036661, 0.2864788, 0.315922, 0.2406943,
  -0.08022118, -0.2270312, -0.3537073, -0.315588, -0.4771933, -0.3641887, 
    0.2133502, 0.4649942, 0.4165241, 0.3558308, 0.7213256, 0.520463, 
    -0.1786419, -0.4806926, -0.5670208, 0.340515, 1.082475, 1.149499, 
    1.003194, 0.8310588, 0.7069051, 0.5358276, 0.3992391, 0.3014364, 
    0.3332236, 0.2930703, 0.1002312, -0.253643, -0.441875, -0.6572561, 
    -1.043813, -0.8074831, -0.3028118, 0.01243889, 0.1001183, 0.1053914, 
    0.07978904, -0.1370403, -0.1077598, 0.4785848, 1.382572, 1.532752, 
    1.020186, 0.5608602, 0.2341354, 0.328064, 0.4883016, 0.4756389, 
    -0.02082896, -0.3401651, -0.252714, -0.3328576, -0.2598755, -0.09708267, 
    0.01055074, 0.1418984, 0.1112506, 0.1192259, 0.2655638, 0.3617715, 
    0.6635944, 0.8530965, 0.850362, 0.9279176, 0.9265504, 0.9211142, 
    0.8237997, 0.8108443, 0.7135782, 0.581254, 0.5158243, 0.3884475, 
    0.4306355, 0.2907104, 0.2576852, 0.3207712, 0.3484745, 0.2399452, 
    -0.09737557, -0.1151165, -0.2251915, -0.1017373, 0.03486717, -0.08910745, 
    -0.008134127, 0.1220418, 0.6713741, 0.8367395, 0.4908407, 0.3270873, 
    0.2078653, 0.253194, 0.2459675, 0.1472862, 0.1296427, -0.03463173,
  -0.1102347, -0.1362114, -0.05426025, 0.1277547, 0.0415892, 0.2264199, 
    0.4145872, 0.2370645, 0.2575235, 0.1170123, 0.3769733, 0.5530804, 
    0.0903852, 0.05470775, 0.167289, 0.6945677, 1.168428, 0.9787638, 
    0.6932496, 0.4354533, 0.2723026, 0.1918173, 0.04072666, -0.06295156, 
    0.005846977, -0.07506227, -0.3084774, -0.5087214, -0.746563, -1.003821, 
    -1.084322, -0.9412723, -0.6395469, -0.2384563, -0.2173787, -0.2596967, 
    -0.05028901, -0.119625, -0.04335535, 0.3279988, 0.4283736, 0.2251997, 
    0.01380658, -0.08746314, -0.2472124, 0.142045, 0.07059312, -0.6136842, 
    -0.9450646, -0.8401655, -0.6440063, -0.4610638, -0.3088177, -0.1831992, 
    0.08227935, 0.2621621, 0.4088256, 0.4940957, 0.5395872, 0.5818073, 
    0.7766153, 0.8965209, 0.8834351, 0.8979859, 0.818103, 0.7490603, 
    0.6445839, 0.556124, 0.4469118, 0.3971395, 0.3517456, 0.3397176, 
    0.3519244, 0.1820016, 0.3531442, 0.2330432, 0.4552778, 0.3227252, 
    -0.3301878, -0.1774045, -0.07766497, -0.03209186, 0.08569729, 0.1253134, 
    0.245772, 0.3298057, 0.7359092, 0.5420773, 0.2211954, 0.1829303, 
    0.1470578, 0.1520059, 0.03550243, -0.02258706, -0.04880762, -0.1816854,
  0.003535986, -0.001151562, -0.001346827, -0.0719524, -0.04447845, 0.109265, 
    0.293591, 0.08675516, 0.1070677, 0.07894278, 0.3018106, 0.7104859, 
    0.1235069, 0.3928425, 0.6775429, 0.7497599, 0.8269733, 0.5687864, 
    0.4036986, 0.1197954, -0.09112525, -0.2126424, -0.4098425, -0.3732054, 
    -0.4416625, -0.4425738, -0.5611777, -0.8926878, -1.001379, -0.9403446, 
    -0.8444134, -0.5673138, 0.08714592, 0.3861535, 0.1596072, -0.01918507, 
    -0.1287229, -0.4136028, -0.220569, -0.02761647, -0.02354741, -0.1207968, 
    -0.3127402, -0.1876588, -0.2529745, -0.2109498, -0.5939902, -1.113163, 
    -0.8149211, -0.452649, -0.466386, -0.2001751, 0.01823315, 0.06354564, 
    0.3555378, 0.3614135, 0.4141153, 0.474597, 0.4580443, 0.6042032, 
    0.7279499, 0.7162802, 0.699337, 0.6125857, 0.4557986, 0.4048543, 
    0.4376669, 0.3963583, 0.3464398, 0.355896, 0.3281615, 0.3434122, 
    0.2788291, 0.1538768, 0.1331096, 0.07674587, -0.09656185, 0.1853068, 
    0.007165551, 0.232621, 0.08320701, 0.0971067, 0.1993365, 0.2301309, 
    0.1577513, 0.1241901, 0.4253132, 0.244112, 0.1160032, 0.02143955, 
    -0.0508585, -0.06933165, -0.06908727, -0.05050039, -0.1239705, -0.09267163,
  0.0291872, -0.003462791, -0.01301694, -0.1861451, -0.08800057, 0.03781313, 
    0.107475, 0.07742953, 0.1028849, 0.1060586, 0.2800986, 0.9487181, 
    0.525769, 0.6365762, 0.5204792, 0.1022663, 0.1919311, 0.1522175, 
    0.1130248, -0.08661705, -0.3105593, -0.3804159, -0.2443811, -0.129114, 
    -0.3541955, -0.4036092, -0.6741988, -1.061357, -0.9429811, -0.8177533, 
    -0.5386354, -0.1209108, 0.2963742, 0.2732303, 0.01237404, -0.226249, 
    -0.5331826, -0.6093708, -0.192265, -0.1439413, -0.3221804, -0.3739218, 
    -0.3523235, -0.1973919, -0.4725547, -0.5862103, -0.6366009, -0.5951295, 
    -0.3241823, -0.0793255, -0.04680604, 0.1907592, 0.3711628, 0.3471231, 
    0.4414753, 0.4521036, 0.4831583, 0.4321492, 0.3689004, 0.3883339, 
    0.4530964, 0.4830608, 0.5105675, 0.5124718, 0.5181358, 0.4958534, 
    0.4349976, 0.4052453, 0.3968632, 0.3857787, 0.3269572, 0.2576048, 
    0.1461792, 0.0649457, -0.0372839, 0.04287507, 0.1930704, 0.1076536, 
    0.1381387, 0.1702188, 0.1040241, 0.1765502, 0.1859578, 0.1437051, 
    -0.04937768, 0.1054239, 0.2029174, 0.06387116, 0.09855533, 0.04792047, 
    0.1075401, 0.02664816, 0.01141357, -0.0051229, -0.07120371, 0.04502392,
  -0.0004193783, -0.1260211, -0.2449505, -0.2307903, 0.01476622, 0.06478262, 
    0.009085894, -0.04595965, -0.007076144, 0.04282618, 0.4684285, 1.154692, 
    0.7308962, 0.4602418, 0.2145221, -0.01348895, 0.1375365, 0.2165893, 
    0.07908927, 0.05697012, -0.05562755, -0.09701751, 0.0386433, -0.1719687, 
    -0.4224244, -0.3910605, -0.5711875, -0.3699667, -0.1818645, -0.5766074, 
    -0.1918743, 0.3137572, 0.2584024, -0.05074477, -0.3637004, -0.2467083, 
    -0.1584433, -0.04778248, 0.01966545, -0.105058, -0.5042925, -0.4852659, 
    -0.2617799, -0.2636516, -0.6727172, -0.7248333, -0.7544228, -0.8228476, 
    -0.8248656, -0.6382446, -0.5010048, -0.2693807, -0.04317629, 0.1140665, 
    0.2853391, 0.3972858, 0.4515339, 0.3549031, 0.3618692, 0.2966837, 
    0.2241413, 0.1369343, 0.1248412, 0.1925983, 0.215336, 0.2406288, 
    0.1805542, 0.1692101, 0.1654174, 0.1652548, 0.139246, 0.03652787, 
    -0.07043839, -0.2345004, -0.2541461, 0.03620188, 0.008841813, 0.03708079, 
    0.09502351, 0.09839265, 0.192045, 0.1316934, 0.1052937, 0.1418497, 
    -0.04540628, -0.003934622, -0.03079045, -0.06970632, 0.006612062, 
    0.05638418, 0.1118529, 0.02573627, 0.06626368, 0.1118855, 0.06525505, 
    0.05631936,
  -0.05927342, -0.1748008, -0.2576946, -0.03121346, 0.0519082, -0.009875584, 
    -0.04628509, -0.06868093, 0.09556061, 0.2835489, 0.3813841, 0.442143, 
    0.5157106, 0.6177921, 0.595561, 0.6079307, 0.5327186, 0.3547727, 
    0.02448308, -0.04216725, -0.01414001, -0.07927674, -0.03059494, 
    -0.08747971, -0.08580345, -0.09706633, -0.2868775, -0.04566659, 
    -0.1329547, -0.5426228, -0.1177695, 0.001045614, -0.01479095, 0.1005411, 
    -0.2908494, -0.1554974, -0.06547457, -0.02735603, -0.04242754, 
    -0.5696735, -0.7836385, -0.6674759, -0.5354774, -0.4910111, -0.678267, 
    -0.6984658, -0.7264607, -0.8273234, -0.7797482, -0.7322547, -0.7342732, 
    -0.63761, -0.6554481, -0.5777301, -0.3985634, -0.2772906, -0.1465942, 
    -0.1203737, -0.1340944, -0.1717246, -0.2190228, -0.2652793, -0.3204225, 
    -0.3014609, -0.2654257, -0.2177206, -0.2352174, -0.1026978, -0.01991791, 
    -0.05754811, -0.1456504, -0.1715782, -0.04355085, -0.1552696, -0.2322388, 
    -0.05886647, 0.08634837, 0.2038614, 0.1828002, 0.1804076, 0.1332885, 
    0.09463274, -0.08570576, -0.3271767, -0.1355917, -0.2302043, -0.2385705, 
    -0.2290488, -0.1727826, -0.06449798, -0.03105071, 0.02209055, 
    0.006725907, -0.06612569, -0.06887633, -0.05816656,
  0.2541544, 0.1609907, 0.02866638, 0.06950268, 0.02016999, -0.01125905, 
    0.02049551, 0.09586985, 0.3765177, 0.2832884, -0.05670175, -0.07877219, 
    0.3458536, 0.6356816, 0.6055856, 0.7907267, 0.8027062, 0.5909224, 
    0.3656781, 0.1903363, 0.1454145, 0.05631924, -0.04547119, -0.03059483, 
    0.08213317, 0.1106648, 0.00618881, -0.08515233, -0.2391562, -0.3194799, 
    -0.1173134, -0.0012981, 0.002542913, 0.1524456, -0.1127563, -0.2820923, 
    -0.3087037, -0.1915483, -0.09597588, -0.2532349, -0.3277147, -0.3445597, 
    -0.4994915, -0.5664184, -0.6090128, -0.5876098, -0.5201619, -0.5100384, 
    -0.3487427, -0.149231, -0.05608273, -0.02613521, -0.1058064, -0.312691, 
    -0.5083617, -0.6158815, -0.7064576, -0.7414675, -0.7665, -0.7886841, 
    -0.8467571, -0.7664348, -0.7517376, -0.7669719, -0.7044556, -0.5701946, 
    -0.4218385, -0.2414348, -0.08689383, 0.00698638, 0.02664787, -0.02397072, 
    0.009313866, 0.1314492, 0.3007201, 0.04787182, 0.3718138, 0.7385782, 
    0.4116899, 0.3033243, 0.2267456, -0.03122938, -0.2029579, -0.1047173, 
    0.03356504, -0.1668904, -0.1935341, -0.2727988, -0.2939086, -0.2673625, 
    -0.2386354, -0.1710735, -0.1145305, 0.1089883, 0.2779502, 0.3511109,
  0.1758666, 0.1404988, 0.0656127, -0.01415618, 0.009623051, 0.1091837, 
    0.1111203, 0.1426475, 0.05586362, 0.02357167, 0.1535358, 0.2638711, 
    0.3426311, 0.490027, 0.4557495, 0.6073761, 0.9476266, 1.066866, 
    0.8542035, 0.5696819, 0.4667363, 0.423995, 0.2467816, 0.08188868, 
    0.05791426, 0.1017292, 0.05693752, 0.08532286, -0.01243067, -0.2842402, 
    -0.374249, -0.1139605, -0.01695549, 0.2357626, 0.2966018, 0.1488309, 
    0.1521037, 0.1678588, 0.1764848, 0.2096553, 0.1220093, 0.05132151, 
    -0.06977272, -0.3070111, -0.3764935, -0.3500133, -0.3013473, -0.2969041, 
    -0.2229786, -0.08638954, 0.03159571, 0.1193888, 0.2441936, 0.2788942, 
    0.1003296, -0.09175992, -0.4043255, -0.6194458, -0.799003, -0.8631632, 
    -0.9498495, -0.9882607, -0.9435831, -0.8281859, -0.8380494, -0.7623495, 
    -0.6344362, -0.5023562, -0.2239056, 0.01803774, 0.2505738, 0.5138386, 
    0.4695027, 0.3415406, 0.8866091, 0.1808145, 0.1461635, 0.4428921, 
    0.3087118, -0.135103, -0.1660767, 0.01007891, 0.654496, 0.4722204, 
    0.2901568, 0.1904826, 0.1318886, 0.05630302, 0.07808018, 0.02189517, 
    0.06649184, -0.03105032, -0.009924471, 0.2464395, 0.1959187, 0.1852904,
  0.3694052, 0.147579, -0.07486558, -0.1189737, -0.2119915, -0.1785767, 
    -0.1035112, -0.1056924, -0.1764607, 0.04460073, 0.1827188, 0.3207071, 
    0.2793985, 0.2796102, 0.2184615, 0.2194386, 0.4717803, 0.7372427, 
    0.7639847, 0.6281619, 0.6249387, 0.4816611, 0.4854853, 0.3010457, 
    0.1091349, -0.2472463, -0.1784139, 0.07301807, 0.1590209, -0.1099892, 
    -0.3167763, -0.1035457, -0.1257935, 0.1392784, 0.2182159, 0.0229373, 
    0.05348706, 0.1297231, 0.2568882, 0.2165885, 0.1674509, 0.1718454, 
    0.1834836, 0.0775094, -0.009892464, -0.05528641, -0.07361317, 
    -0.08380222, -0.05997419, -0.03572273, 0.0233593, 0.09258127, 0.1257529, 
    0.3229527, 0.4480181, 0.475915, 0.3354039, 0.08514357, -0.1919885, 
    -0.3185186, -0.38027, -0.5146122, -0.5926561, -0.5822387, -0.7193806, 
    -0.7691205, -0.8299111, -0.7070597, -0.3286581, 0.03159571, 0.2231324, 
    0.5801148, 1.188545, 0.6003938, 0.04997134, -0.11746, -0.5032022, 
    -0.4715779, -0.2747355, -0.0616982, 0.2603719, 0.3871624, 0.4392285, 
    0.2775431, 0.1768746, 0.07726574, 0.009931564, -0.02078152, -0.007321358, 
    0.005553246, 0.2015982, 0.3513224, 0.4554888, 0.3862995, 0.3703492, 
    0.3817754,
  0.2940795, 0.2775109, 0.1699259, 0.05827236, -0.170228, -0.2655077, 
    -0.2631958, -0.1594043, -0.100142, -0.2525511, -0.1546674, 0.07581778, 
    0.127071, 0.01696336, 0.1713252, 0.0847044, 0.07610989, 0.3066435, 
    0.5634155, 0.4325073, 0.3074095, 0.538285, 0.8425815, 0.4843466, 
    0.4314008, 0.1026406, -0.177942, -0.1785113, -0.1763303, -0.4255977, 
    -0.5301719, -0.2307267, -0.4048948, -0.1329386, 0.0372107, -0.1413054, 
    -0.1068983, -0.06134129, 0.0791707, 0.07842112, 0.1818726, 0.1670117, 
    0.1486857, 0.1032593, 0.01728916, -0.01811075, -0.04392505, -0.04202032, 
    -0.02455616, 0.05773497, 0.07905674, 0.09163809, 0.1305542, 0.2522011, 
    0.32393, 0.4147012, 0.4326539, 0.3261435, 0.1704957, 0.03719425, 
    -0.1433239, -0.2810669, -0.3257608, -0.375061, -0.5587211, -0.7069788, 
    -0.8601522, -0.8694131, -0.6578084, 0.1528358, 0.7111862, 0.3654661, 
    0.4862018, -0.0251112, -0.6783004, -0.4128537, -0.2850705, -0.1373004, 
    0.2518272, 0.7021853, 0.841378, 0.6021528, 0.3723187, 0.2411175, 
    0.1214073, -0.0960896, -0.1939569, -0.2653599, -0.3371701, -0.2953897, 
    -0.2468395, 0.05312824, 0.3038619, 0.225704, 0.2499228, 0.3019738,
  0.2646363, 0.2471724, 0.29338, 0.4136758, 0.2496624, -0.1083941, 
    -0.3025513, -0.2642701, -0.1753712, -0.2251606, -0.4441202, -0.07327086, 
    0.01475006, -0.1062298, 0.08503032, 0.1158569, -0.0563283, -0.1509409, 
    0.1927114, 0.2540398, 0.1566446, 0.5338745, 0.8818567, 0.5031946, 
    0.6678104, 0.3798379, -0.09592703, -0.2953571, -0.52301, -0.7972794, 
    -0.8630004, -0.434453, -0.5861778, -0.5129027, -0.2962861, -0.4856737, 
    -0.4577928, -0.3811977, -0.2711551, -0.2116008, -0.1541951, -0.09910083, 
    0.03532314, -0.04620361, -0.2187297, -0.268518, -0.2603149, -0.2470987, 
    -0.3015585, -0.1853964, -0.04719663, 0.03932714, 0.1769083, 0.3315473, 
    0.4467816, 0.5829308, 0.7405479, 0.7170942, 0.4813192, 0.2629108, 
    0.1229043, 0.03188801, -0.04042578, -0.05673504, -0.1332645, -0.3452106, 
    -0.6181281, -0.9066694, -0.7150836, -0.007076144, 0.3923542, 0.0884645, 
    -0.1535927, -0.5193319, -0.550159, -0.2411744, 0.07873119, 0.5326049, 
    0.7374876, 0.7047241, 0.6051149, 0.618901, 0.578048, 0.2758832, 
    -0.02156162, -0.2066855, -0.4409628, -0.6114542, -0.6807904, -0.6860313, 
    -0.6828265, -0.4455209, -0.04372978, 0.2123086, 0.3554077, 0.3611856,
  0.5198607, 0.3508503, 0.149158, 0.1408405, 0.1915734, -0.01815975, 
    -0.2369423, -0.2719359, -0.2035112, -0.1920547, -0.3508601, -0.04727757, 
    0.01164134, -0.2348757, -0.07803988, 0.1164591, -0.1844683, -0.5227985, 
    -0.03191328, 0.2876496, 0.07402778, 0.1211953, 0.2107298, 0.2957396, 
    0.4138061, 0.0383015, 0.07179759, 0.06367588, -0.2173463, -0.5948696, 
    -0.7042766, -0.394804, -0.463604, -0.7002723, -0.7015095, -0.7958779, 
    -0.7759073, -0.7331829, -0.6408486, -0.5006309, -0.4018025, -0.3104451, 
    -0.2023885, -0.1747518, -0.2058389, -0.285917, -0.3394165, -0.4584761, 
    -0.5564574, -0.4412556, -0.2587035, -0.103056, 0.03898525, 0.2380574, 
    0.4709516, 0.6005249, 0.7410357, 0.8924682, 0.8534713, 0.7373741, 
    0.5439656, 0.3218465, 0.1255898, 0.1096549, 0.04904318, -0.0648241, 
    -0.1057916, -0.3146443, -0.02971619, 0.05770254, 0.05509877, 0.2795128, 
    -0.020455, -0.5477986, -0.480546, -0.3026813, -0.02040631, 0.4414753, 
    0.6044636, 0.8224487, 1.049955, 0.9256874, 0.7389363, 0.6260946, 
    0.4128298, 0.1367556, -0.3528115, -0.6062462, -0.6936157, -0.8888142, 
    -0.8873, -0.6250448, -0.07917881, 0.2038778, 0.2113488, 0.4297891,
  0.1320355, 0.38197, 0.3778523, 0.1695356, 0.09058046, -0.07291281, 
    -0.3621706, -0.4071734, -0.4410276, -0.3153932, -0.2931447, -0.2000775, 
    -0.08969329, -0.2278932, -0.1416135, 0.002640545, -0.1863568, -0.3580527, 
    -0.1533163, -0.02117085, 0.1437056, 0.2276407, 0.2242391, 0.3347859, 
    -0.09359962, -0.3526979, -0.1111125, -0.2885702, -0.252063, 0.0173707, 
    -0.1639605, -0.2690077, -0.1127086, -0.2376437, -0.4124634, -0.4486775, 
    -0.4398723, -0.4729779, -0.544543, -0.5689905, -0.5303832, -0.442997, 
    -0.419413, -0.3808552, -0.3874147, -0.3634887, -0.2936647, -0.5075316, 
    -0.7546182, -0.8353474, -0.7528604, -0.4755981, -0.2364218, 0.004723966, 
    0.3430378, 0.621586, 0.8018594, 0.8788288, 0.8161824, 0.7524126, 
    0.6498737, 0.5601118, 0.4208374, 0.3259802, 0.04928684, -0.1487112, 
    0.002542973, 0.02417397, 0.1278686, 0.09910893, 0.1867715, 0.4697306, 
    0.06761456, -0.1640911, -0.1106079, -0.2237103, -0.1403443, 0.1144083, 
    0.3868041, 0.6235065, 0.8447468, 0.8851601, 0.8217813, 0.652836, 
    0.3710326, 0.1571654, -0.243502, -0.6161419, -0.8368285, -1.03219, 
    -0.9869425, -0.7879841, -0.2720337, 0.124369, 0.08929467, 0.001582861,
  -0.05759668, 0.03463972, 0.2464883, 0.1783894, 0.1130248, -0.0785442, 
    -0.4404583, -0.5183555, -0.5679649, -0.4126422, -0.2694786, -0.3431764, 
    -0.2251263, -0.05717397, -0.1527956, -0.2826783, -0.2138959, -0.1563108, 
    -0.2303672, -0.1272907, 0.2315793, -0.01254475, -0.2477336, -0.2693808, 
    -0.3119588, -0.3314251, -0.02834892, -0.2878385, -0.2463665, 0.2142773, 
    0.1647177, 0.1239624, 0.3204293, 0.3383341, 0.1025257, -0.0326457, 
    -0.05727124, -0.05046773, -0.06173074, -0.07608664, -0.1339478, 
    -0.2161744, -0.366679, -0.4147584, -0.4436321, -0.4396282, -0.3179322, 
    -0.2780885, -0.3653769, -0.635429, -0.7703086, -0.6456178, -0.535136, 
    -0.2223756, 0.1600626, 0.3890668, 0.5823611, 0.7311893, 0.7320518, 
    0.6862832, 0.6150104, 0.526469, 0.39644, 0.2631063, 0.09364033, 
    0.09915733, 0.1215701, 0.08338612, 0.05856517, -0.1582154, -0.09879172, 
    -0.02891827, -0.3772744, -0.2078412, 0.1492064, 0.1513874, 0.1543985, 
    0.2457884, 0.4548541, 0.4984415, 0.5117389, 0.6680704, 0.6607949, 
    0.4002318, 0.1493204, 0.08210033, -0.2277791, -0.7104616, -0.8326132, 
    -0.8192343, -0.7951783, -0.6822712, -0.3587036, 0.07900786, 0.2285359, 
    0.1356652,
  0.5120158, 0.2955933, 0.08060288, -0.108427, -0.05487884, -0.2307579, 
    -0.6972616, -0.8677369, -1.002389, -0.6325481, -0.3512493, -0.3776653, 
    -0.3795696, -0.1012656, -0.07445902, -0.2962689, -0.2732545, -0.06783457, 
    -0.2470501, -0.3538375, -0.02654219, -0.2936808, -0.5931118, -0.6020792, 
    -0.7391236, -0.8845339, -0.6769328, -0.2912068, 0.007409573, 0.09946728, 
    0.1386598, 0.04940224, 0.2510452, 0.527739, 0.4098997, 0.4281607, 
    0.3798699, 0.2937865, 0.2676148, 0.2050985, 0.1611205, 0.113383, 
    -0.06293559, -0.1675906, -0.1956666, -0.299426, -0.3474407, -0.2182413, 
    -0.09820557, -0.2122358, -0.28442, -0.3888471, -0.567265, -0.3091433, 
    0.08659267, 0.2560589, 0.4419639, 0.5521362, 0.5238814, 0.5138716, 
    0.4824748, 0.4931843, 0.515092, 0.4036827, 0.1205447, -0.06028247, 
    -0.1231732, -0.1998984, -0.203121, -0.2694784, -0.2592246, -0.05523688, 
    -0.1566203, -0.1532187, 0.03089589, 0.2676634, 0.3922566, 0.3949421, 
    0.5293498, 0.7338583, 0.7972697, 0.6915568, 0.5838747, 0.3420614, 
    -0.005448222, -0.1425741, -0.4040811, -0.9728963, -1.132792, -0.8449992, 
    -0.5464154, -0.3233847, -0.1382935, 0.09674877, 0.2581258, 0.4317911,
  0.6244017, 0.8580606, 0.5899615, 0.3629273, 0.3828328, 0.1905801, 
    -0.4979452, -0.7143677, -0.7690715, -0.8334755, -0.3805135, -0.1965943, 
    -0.2880006, -0.06679285, 0.1857949, 0.05425203, -0.03782165, 0.0943886, 
    0.03778064, -0.09143482, 0.0275104, 0.09971094, 0.01566195, 0.04984128, 
    -0.07745373, -0.3374957, -0.2831342, -0.1218385, 0.07091868, 0.2601763, 
    0.3838094, 0.2390018, 0.3661013, 0.5882678, 0.4957061, 0.4168005, 
    0.2113646, 0.2051146, 0.4639854, 0.2934287, 0.0893594, 0.1533895, 
    0.157263, 0.070333, -0.005708933, -0.07799053, -0.1354284, -0.1319621, 
    -0.08608007, -0.02797413, 0.1202517, 0.1472051, -0.05847526, -0.0210731, 
    0.1902058, 0.3996136, 0.6391315, 0.6842155, 0.5749388, 0.4210653, 
    0.2827842, 0.3809451, 0.5346069, 0.3985553, 0.112097, 0.04204506, 
    -0.06109625, -0.1454387, -0.2299602, -0.555009, -0.6088827, -0.143567, 
    0.08839905, -0.06921792, -0.1265261, -0.008052677, 0.3159219, 0.621586, 
    0.7131224, 0.8645387, 1.023897, 0.9777386, 0.8071003, 0.4967163, 
    0.08146572, -0.03181553, -0.09073472, -0.6143839, -1.117167, -1.032499, 
    -0.5962195, -0.1337687, 0.2951374, 0.5799681, 0.5598021, 0.4365436,
  0.7803099, 1.302543, 1.136723, 0.8457069, 0.9704468, 0.7006224, 0.04082429, 
    0.07725006, -0.1225709, -0.6246379, -0.4746054, -0.1254188, -0.05767822, 
    0.06894928, 0.2482625, 0.2157591, 0.09575588, 0.06312251, 0.1292684, 
    0.4055054, 0.314425, -0.03163671, -0.08171809, 0.02057678, 0.2742065, 
    0.2977415, 0.2231811, -0.05927339, -0.2638307, -0.1201947, 0.1704311, 
    0.1694214, 0.1326213, 0.08354902, 0.1128783, 0.6151886, 0.4204142, 
    0.2111368, 0.5035033, 0.6150267, 0.4502647, 0.3482299, 0.24753, 
    0.03613679, -0.1115847, -0.1356893, -0.2094197, -0.2610469, -0.1542115, 
    -0.00902915, 0.2045777, 0.4746134, 0.509721, 0.4815633, 0.6007853, 
    0.7165899, 0.6753616, 0.604496, 0.6218295, 0.450932, 0.1774292, 
    0.2095096, 0.3028038, 0.1378621, -0.04346931, -0.2027141, -0.3247194, 
    -0.3050741, -0.3111777, -0.6018838, -0.736259, -0.3953899, 0.04466534, 
    0.1387576, 0.08304477, 0.07440168, 0.2723184, 0.4889038, 0.5716186, 
    0.6566283, 0.8541869, 0.8980672, 0.7467488, 0.5455122, 0.3112342, 
    0.07409263, -0.1411254, -0.4025683, -0.7583134, -0.9293096, -0.7627892, 
    -0.3655396, 0.1804893, 0.7265668, 0.8197308, 0.6737345,
  1.068428, 1.458728, 1.2467, 1.084281, 1.386642, 1.028455, 0.3105346, 
    0.2975788, 0.2828002, -0.04649627, -0.009159088, -0.003951073, 
    -0.09005141, 0.05687246, 0.2561889, 0.228601, 0.3008178, 0.2536173, 
    0.1147016, 0.2217815, -0.03995371, 0.02405977, 0.02272534, -0.08363867, 
    -0.09193939, 0.06554759, 0.05796289, -0.1568157, -0.2603801, -0.1744915, 
    0.02386463, 0.07604575, 0.02456474, 0.04201281, 0.1138223, 0.2556844, 
    0.3032594, -0.01003838, -0.06347257, 0.2831582, 0.3353722, 0.3897012, 
    0.4921426, 0.2854694, -0.007857352, -0.0006797314, 0.01929116, 
    -0.1266396, -0.1381142, -0.05826402, 0.2095098, 0.6678753, 0.9242067, 
    0.8909872, 1.002299, 1.221879, 1.231189, 1.080897, 0.9902544, 0.8517776, 
    0.6422899, 0.4201701, 0.1349001, -0.140686, 0.0983603, -0.06394434, 
    -0.4223914, -0.486422, -0.3143679, -0.3457316, -0.4961224, -0.5221314, 
    -0.3471152, -0.1037071, 0.1286497, 0.1829792, 0.2297565, 0.3983438, 
    0.7118853, 0.8336629, 0.8408895, 0.8102904, 0.6893108, 0.5056031, 
    0.3587928, 0.2363319, 0.1201701, -0.03988886, -0.3537078, -0.6336231, 
    -0.6763477, -0.4610643, -0.06130791, 0.6310759, 1.159265, 1.076567,
  1.017143, 1.226127, 0.9095905, 0.7055704, 1.144177, 1.07904, 0.6323769, 
    0.5507201, 0.5314655, 0.2287964, 0.07952905, 0.03616977, -0.02929258, 
    0.001403511, 0.1622436, 0.2114952, 0.3267128, 0.3691446, 0.148002, 
    -0.1408648, -0.1803019, 0.05171371, 0.09126425, -0.0384239, -0.05536713, 
    0.1018757, 0.1043171, -0.06786704, -0.1339966, -0.0271771, 0.03350008, 
    -0.05717349, -0.03137589, 0.02113068, 0.01824942, 0.02913809, 0.08859468, 
    0.144567, 0.06531858, 0.115449, 0.2199426, 0.4046427, 0.6680376, 
    0.6245807, 0.255668, -0.02566335, -0.1458945, -0.2462363, -0.2942992, 
    -0.224996, 0.02292097, 0.5286664, 0.9898156, 1.105522, 1.066378, 
    1.146945, 1.259673, 1.212684, 1.088546, 1.009103, 0.9539752, 0.6404328, 
    0.1520386, -0.1162231, 0.2206094, -0.09965396, -0.1719358, -0.188977, 
    -0.2290977, -0.2624471, -0.1369265, -0.0636679, -0.1101197, -0.1874635, 
    0.06577544, 0.2555541, 0.2077839, 0.1544962, 0.2797077, 0.4563355, 
    0.727478, 0.8716022, 0.8380572, 0.5132202, 0.1754601, 0.05882549, 
    -0.0216918, -0.293828, -0.6099415, -0.7717748, -0.8213835, -0.8262162, 
    -0.595016, -0.01993418, 0.5253119, 0.7342491,
  0.5637741, 0.6925502, 0.6239948, 0.4849162, 0.7183799, 0.8683962, 
    0.7821006, 0.7655153, 0.6154338, 0.1914918, -0.03508687, -0.04101133, 
    -0.02836537, -0.009598732, 0.1685586, 0.272563, 0.1427615, 0.01221156, 
    -0.08673096, -0.2016889, -0.2748657, -0.1756792, -0.08135986, 
    -0.05709243, 0.06271601, -0.06158423, -0.1284624, -0.1855104, -0.1901328, 
    -0.1289349, -0.1243447, -0.08852148, -0.06851816, -0.1422, -0.2638309, 
    -0.1206992, 0.02978912, -0.09913301, -0.9440241, -0.546041, 0.1206083, 
    0.1268437, -0.006847858, 0.1316612, 0.3022174, 0.1573118, -0.1591269, 
    -0.4038372, -0.5302043, -0.5596152, -0.2995241, 0.2521849, 0.8731487, 
    1.272791, 1.387439, 1.3453, 1.317582, 1.266475, 1.230083, 1.280148, 
    1.14548, 0.6508183, 0.04328275, -0.2004678, -0.2812781, -0.285445, 
    -0.1486776, 0.01434314, 0.01281321, -0.08757743, -0.03835866, 0.09071034, 
    0.1072305, 0.159379, 0.313741, 0.4212605, 0.3192748, 0.2062214, 
    0.1648803, 0.2676959, 0.6928266, 0.6977092, 0.8729044, 0.5360066, 
    0.1890664, 0.1709841, 0.209851, -0.1029906, -0.5031214, -0.6313605, 
    -0.6643529, -0.7998338, -0.8020968, -0.4390264, -0.07104111, 0.206759,
  0.2104697, 0.3147337, 0.2504272, 0.2013714, 0.3734251, 0.4611044, 
    0.4805541, 0.5280477, 0.3505738, 0.07835686, -0.09727764, -0.1471636, 
    -0.2036252, -0.2225378, 0.007865191, 0.1907759, 0.2298219, 0.2017622, 
    0.1186891, -0.0806272, -0.3827267, -0.481425, -0.3129692, -0.01101494, 
    -0.002697468, -0.1854124, -0.2161739, -0.1193316, -0.164905, -0.1659628, 
    -0.1203737, -0.004097462, -0.1131308, -0.3514769, -0.49915, -0.2849245, 
    -0.2069948, -0.6510372, -1.20509, -0.6800594, 0.4384146, 0.4019737, 
    -0.2500281, -0.5676391, -0.4561968, -0.3673947, -0.4182576, -0.4713992, 
    -0.5647421, -0.6413372, -0.384957, 0.2838581, 1.072823, 1.672774, 
    1.997595, 1.976208, 1.588318, 1.167061, 1.011804, 1.17406, 1.163595, 
    0.7748253, 0.2089071, 0.03276777, 0.07562256, 0.1126182, -0.03044862, 
    -0.1703574, -0.09075124, 0.1312051, 0.2742878, 0.3068562, 0.3718301, 
    0.4945351, 0.3850463, 0.3891641, 0.1471719, 0.282019, 0.3375528, 
    0.2150105, 0.3295128, 0.5944867, 0.9852419, 0.5891151, 0.1061726, 
    0.05916727, 0.1705935, 0.0300982, -0.3175089, -0.4706671, -0.5417767, 
    -0.7234173, -0.808835, -0.590508, -0.2467895, 0.01269937,
  -0.1010213, 0.09416103, 0.06190205, 0.01603591, 0.0475136, 0.1941609, 
    0.1488321, 0.1314007, -0.1392051, -0.1711876, -0.09776628, -0.07532179, 
    -0.0906049, -0.1222613, -0.07139874, 0.03932714, 0.1409383, 0.1359093, 
    0.09753013, -0.07982969, -0.238049, -0.3146603, -0.22052, -0.09623623, 
    -0.1014602, -0.2260861, -0.2438598, -0.2807411, -0.2752236, -0.2587035, 
    -0.2874309, -0.2635377, -0.2779582, -0.3079222, -0.2810344, -0.3137814, 
    -0.6112914, -1.100044, -1.567688, -1.970764, -1.514678, -1.255008, 
    -0.8077273, -0.9296997, -1.248564, -0.9923959, -0.6392207, -0.1629674, 
    0.1182172, 0.22157, 0.4698124, 1.042794, 1.64377, 2.02017, 1.881531, 
    2.108289, 1.802462, 1.319405, 0.9884969, 0.9633994, 0.9417849, 0.6857789, 
    0.4423709, 0.2861043, 0.3679402, 0.4021524, 0.2277708, -0.01802987, 
    -0.01485604, 0.1121622, 0.08913156, -0.2376101, -0.4067992, -0.5872356, 
    -0.5981891, -0.4098431, -0.2638795, 0.1593463, 0.2269408, -0.04849863, 
    -0.4207153, 0.2405963, 0.8913937, 0.8175011, 0.4132853, 0.1068885, 
    0.04157298, -0.02758384, -0.1901975, -0.2603314, -0.3877401, -0.7005825, 
    -0.9951952, -0.980921, -0.7200809, -0.3746054,
  -0.4991982, -0.365751, -0.2326946, -0.2183228, -0.05469978, 0.1265175, 
    0.2115273, 0.002689421, -0.2817996, -0.4063928, -0.4051231, -0.3456017, 
    -0.3638794, -0.3830364, -0.3211385, -0.181425, -0.1018513, -0.0861938, 
    -0.08381772, -0.1419718, -0.1992309, -0.2328733, -0.2627074, -0.2396604, 
    -0.2139605, -0.3004189, -0.2796346, -0.3072228, -0.3420535, -0.379146, 
    -0.3961548, -0.3417279, -0.2544394, -0.2450319, -0.2371706, -0.2112591, 
    -0.186161, -0.3747027, -0.645618, -0.9804153, -1.256767, -1.363653, 
    -1.413911, -1.470634, -1.588782, -1.627503, -1.686894, -2.065735, 
    -1.694007, -1.279064, -0.724328, 0.008239985, 0.8552942, 0.9550658, 
    0.7539916, 0.6478882, 0.6612182, 0.699532, 0.5576211, 0.5679727, 
    0.6310261, 0.4982626, 0.3257041, 0.2064166, 0.2555215, 0.3047403, 
    0.1903197, 0.02402741, -0.1545371, -0.3196575, -0.5871052, -0.670097, 
    -0.7637492, -0.7089641, -0.5225219, -0.1913534, 0.01756573, 0.09207749, 
    -0.05925679, -0.4501424, -0.9289184, -0.5684204, 0.06859136, 0.4236857, 
    0.07560658, -0.3529739, -0.6837356, -0.7861126, -0.671334, -0.4407188, 
    -0.3713504, -0.5612748, -0.8623002, -1.026753, -0.9373002, -0.7090614,
  -0.2016397, -0.4725871, -0.6836548, -0.5668254, -0.4357052, -0.332792, 
    -0.06433511, -0.4224408, -0.4448854, -0.3926719, -0.2843224, -0.2277789, 
    -0.2282838, -0.2970496, -0.4127562, -0.4971637, -0.5078576, -0.467916, 
    -0.3809856, -0.2425255, -0.2362589, -0.2128212, -0.2563274, -0.2726033, 
    -0.3245074, -0.461454, -0.4844687, -0.4766888, -0.4823691, -0.4399374, 
    -0.4733033, -0.5170697, -0.5310181, -0.5725546, -0.5881959, -0.574345, 
    -0.619625, -0.462431, -0.3829388, -0.395292, -0.5112267, -0.8435996, 
    -1.012024, -1.227161, -1.50387, -1.841403, -2.046888, -2.297555, 
    -2.377892, -2.214351, -1.660803, -1.264172, -0.0567174, 0.3345093, 
    0.378959, 0.3322142, 0.2171101, 0.2154662, 0.2608437, 0.2428914, 
    0.1943561, 0.1522339, 0.1277058, 0.131254, 0.1381387, 0.1405964, 
    0.05633536, -0.09371347, -0.2821087, -0.4312299, -0.4579548, -0.4726359, 
    -0.4900998, -0.3535602, -0.2638628, -0.1710085, 0.04700905, 0.002738357, 
    -0.05491126, -0.06833863, 0.03130269, 0.3272178, 0.2855671, 0.1505736, 
    -0.1778769, -0.6342084, -0.9240351, -0.9114556, -0.4271946, 0.1431518, 
    0.4819052, 0.384444, 0.4904337, 0.3907266, 0.2183796, 0.03533936,
  1.104675, 0.6686563, 0.2207723, -0.1323202, -0.3966758, -0.4335728, 
    -0.5065386, -0.608052, -0.6426554, -0.5351518, -0.2711549, 0.3048543, 
    0.7179403, 0.9003292, 0.5055218, 0.3741412, 0.05648232, -0.2612264, 
    -0.4878705, -0.6097944, -0.5550903, -0.4505813, -0.332011, -0.2695758, 
    -0.3025188, -0.3643675, -0.3923459, -0.3588665, -0.3557577, -0.4104778, 
    -0.5879843, -0.773873, -0.9204062, -1.007109, -0.9345826, -0.9114546, 
    -0.7107382, -0.6754518, -0.5553508, -0.5697064, -0.6227012, -0.6340944, 
    -0.7331992, -0.8505332, -0.9998007, -1.088001, -1.213033, -1.302584, 
    -1.497929, -1.339953, -1.333117, -1.199247, -0.7491004, -0.3593223, 
    -0.106181, 0.02856839, 0.0001341105, -0.05229092, 0.06077871, 0.09660228, 
    0.1124389, 0.1218953, 0.1260619, 0.1391153, 0.1684936, 0.1997598, 
    0.1654988, 0.09059644, -0.05015886, -0.1472942, -0.2435019, -0.262317, 
    -0.2563438, -0.2969033, -0.1999469, -0.1160767, -0.08751225, 
    -0.009289622, 0.09958088, 0.1522505, 0.2570028, 0.4357625, 0.3728397, 
    0.3033407, -0.009810209, -0.3533489, -0.4593222, -0.4457822, -0.06251192, 
    0.1359406, 0.052526, 0.1276569, 0.1499884, 0.8780479, 1.377608, 1.373099,
  1.884818, 1.696912, 1.356286, 0.9442096, 0.5814982, 0.3433962, 0.1960491, 
    0.1139364, 0.05218494, 0.07020241, 0.2351439, 0.5696005, 0.8778034, 
    0.8960001, 0.7897015, 0.727999, 0.5908894, 0.3981647, 0.158793, 
    -0.03511989, -0.1523726, -0.2004676, -0.2163694, -0.2897909, -0.3461385, 
    -0.3614867, -0.3049273, -0.261129, -0.2336549, -0.2697877, -0.4019003, 
    -0.5873658, -0.7684692, -0.8916789, -0.9093225, -0.9051555, -0.7691367, 
    -0.6653931, -0.663554, -0.6033815, -0.5178347, -0.531946, -0.5716432, 
    -0.6855267, -0.7857057, -0.8498822, -0.9011517, -0.9409791, -0.9672159, 
    -1.002079, -1.020878, -0.970292, -0.8538697, -0.6891562, -0.5512168, 
    -0.4803835, -0.4686159, -0.4643841, -0.4006471, -0.2870078, -0.1649863, 
    -0.06217051, 0.07051179, 0.1564656, 0.1857462, 0.2184122, 0.1974161, 
    0.1279662, 0.02524817, 0.0170126, -0.1027467, -0.1386679, -0.1102664, 
    -0.1600873, -0.1581665, -0.1171834, -0.09232998, -0.003055573, 
    0.01489687, 0.01219475, 0.1385619, 0.2590536, 0.2141969, 0.1435413, 
    0.01435852, -0.1986125, -0.2410278, -0.06269097, -0.01540899, 
    -0.05658913, -0.08043337, 0.1760283, 0.494226, 0.8199582, 0.8178914, 
    1.413269,
  1.356254, 1.577999, 1.558842, 1.36615, 0.9918007, 0.6545776, 0.4925494, 
    0.3385617, 0.3916543, 0.3824911, 0.4715372, 0.4494506, 0.4728067, 
    0.4637084, 0.4535684, 0.4141966, 0.4540403, 0.4264199, 0.4024128, 
    0.3415241, 0.2799518, 0.2269083, 0.1495806, 0.03735757, -0.07603741, 
    -0.1203245, -0.1769003, -0.2718225, -0.3161744, -0.3186647, -0.3633424, 
    -0.3631471, -0.4390911, -0.551526, -0.6695924, -0.7966595, -0.8924115, 
    -0.9824668, -1.032939, -1.045748, -1.019951, -0.9894329, -0.946399, 
    -0.8841107, -0.8361126, -0.8011029, -0.7620404, -0.7315066, -0.6924114, 
    -0.6466269, -0.6113405, -0.5741009, -0.5328736, -0.4958945, -0.4759401, 
    -0.4653118, -0.4718548, -0.4665977, -0.4455202, -0.404, -0.3393028, 
    -0.2574342, -0.1728476, -0.1040813, -0.03396413, 0.05998117, 0.1440958, 
    0.2057657, 0.2161173, 0.1854858, 0.1365438, 0.049532, -0.02810472, 
    -0.09392506, -0.1175905, -0.1208783, -0.195504, -0.1873822, -0.03310148, 
    0.05467519, -0.003088474, -0.06651592, -0.1369262, -0.1483195, 
    -0.09405494, -0.01107967, 0.1712604, 0.4210324, 0.6045451, 0.7234247, 
    0.6861525, 0.932539, 1.012731, 1.172431, 1.300802, 1.465466,
  1.471277, 1.437374, 1.410128, 1.1724, 0.9346883, 0.69364, 0.4944701, 
    0.3106322, 0.1990762, 0.1442585, 0.1494506, 0.1883015, 0.2439818, 
    0.3042683, 0.36239, 0.3888386, 0.4045287, 0.4051147, 0.4050007, 
    0.4078327, 0.4208861, 0.4017618, 0.3483925, 0.2891478, 0.2187213, 
    -0.06669521, -0.1802369, -0.2374635, -0.2646609, -0.3164024, -0.3499475, 
    -0.3776816, -0.4102825, -0.4556601, -0.5197715, -0.6069459, -0.7133099, 
    -0.8152956, -0.9052532, -0.9710572, -1.013977, -1.042997, -1.06165, 
    -1.062415, -1.055693, -1.032027, -1.009436, -0.9664023, -0.915442, 
    -0.8696901, -0.8269166, -0.7763958, -0.720927, -0.655302, -0.5934693, 
    -0.5372031, -0.4864381, -0.4401816, -0.4073853, -0.371041, -0.3348267, 
    -0.2844525, -0.2236615, -0.1562299, -0.08391541, -0.010364, 0.05640036, 
    0.101957, 0.1326536, 0.1208047, 0.06709373, 0.09917372, 0.02982169, 
    -0.04701751, -0.09385997, -0.1141075, -0.08140898, -0.02834857, 
    -0.0003867149, 0.05394316, 0.1440308, 0.1559448, 0.1870482, 0.237618, 
    0.2956746, 0.3876507, 0.5191934, 0.6198117, 0.7909056, 0.8609419, 
    0.868608, 0.9295127, 1.084021, 1.276648, 1.397221, 1.475297,
  1.390157, 1.451322, 1.470235, 1.455554, 1.400378, 1.325509, 1.225753, 
    1.121374, 1.008354, 0.9049357, 0.8161172, 0.7414916, 0.6858438, 
    0.6432494, 0.6156453, 0.6031127, 0.5982299, 0.5994668, 0.6013222, 
    0.605131, 0.5965698, 0.5712931, 0.5332723, 0.4611204, 0.3621621, 
    0.2702676, 0.183435, 0.06769598, -0.04602468, -0.1443645, -0.2314414, 
    -0.3226361, -0.4059693, -0.4744264, -0.5412071, -0.5911583, -0.6396446, 
    -0.6899376, -0.720992, -0.7516561, -0.7784467, -0.799931, -0.8244752, 
    -0.8452272, -0.8499147, -0.8596152, -0.8651979, -0.8593222, -0.8410605, 
    -0.8224244, -0.7954388, -0.7527141, -0.699817, -0.6500123, -0.6124472, 
    -0.5801556, -0.5359336, -0.4847454, -0.4297324, -0.3617799, -0.2972128, 
    -0.2414837, -0.20164, -0.1703247, -0.158004, -0.1665326, -0.1910118, 
    -0.2177207, -0.2517865, -0.2935182, -0.3407024, -0.362968, -0.3794394, 
    -0.375289, -0.3085411, -0.3414187, -0.3198529, -0.2235152, -0.1127077, 
    -0.0674274, -0.01583278, 0.01405001, 0.03795958, 0.0802936, 0.1449096, 
    0.1889525, 0.2485717, 0.3099649, 0.3868855, 0.5436235, 0.6628785, 
    0.7983277, 0.9177775, 1.053064, 1.175199, 1.291377,
  1.078943, 1.138838, 1.175525, 1.201957, 1.22852, 1.238969, 1.235713, 
    1.223767, 1.202624, 1.168949, 1.126941, 1.078764, 1.033077, 0.9903522, 
    0.9455932, 0.8841023, 0.8256224, 0.7713418, 0.7154173, 0.6603556, 
    0.6052775, 0.5457723, 0.4875529, 0.4243042, 0.3632038, 0.2953815, 
    0.2151569, 0.141215, 0.08183992, 0.01497781, -0.07343352, -0.1428834, 
    -0.2014282, -0.257548, -0.3178997, -0.3744102, -0.4215456, -0.4624636, 
    -0.5044395, -0.5427696, -0.5788048, -0.6099245, -0.6401492, -0.6664674, 
    -0.6815553, -0.6993777, -0.7092408, -0.7201295, -0.7268841, -0.7286745, 
    -0.721692, -0.715914, -0.7039511, -0.6933391, -0.6848431, -0.6641399, 
    -0.6431438, -0.6205852, -0.5905234, -0.5602825, -0.535787, -0.510136, 
    -0.4886191, -0.4702434, -0.4547812, -0.445927, -0.4499635, -0.4590781, 
    -0.4668417, -0.4737102, -0.4802369, -0.4884889, -0.4889609, -0.4811809, 
    -0.4682903, -0.4539674, -0.4343222, -0.4046184, -0.3687135, -0.3244589, 
    -0.2736614, -0.2147259, -0.1487265, -0.07616788, 0.001664132, 0.08646229, 
    0.1781452, 0.273295, 0.371407, 0.4705443, 0.5675333, 0.6672891, 
    0.7637084, 0.8540728, 0.9362018, 1.011625,
  0.3112371, 0.2749746, 0.2390695, 0.204206, 0.1709542, 0.1408758, 0.1134667, 
    0.08716536, 0.06345081, 0.04144573, 0.02178407, 0.005150557, 
    -0.008423805, -0.02165651, -0.03394508, -0.0459404, -0.05818009, 
    -0.07204735, -0.08822596, -0.1094174, -0.1360123, -0.1687108, -0.207285, 
    -0.252744, -0.3019954, -0.3560971, -0.4118584, -0.468206, -0.5233326, 
    -0.5767021, -0.6276298, -0.674716, -0.7172949, -0.7548761, -0.7872496, 
    -0.8131933, -0.8336525, -0.8460546, -0.8521094, -0.8523703, -0.848887, 
    -0.8388119, -0.8240829, -0.8056583, -0.781846, -0.7545671, -0.7263284, 
    -0.6818781, -0.6401634, -0.5962825, -0.5549088, -0.4844656, -0.4493253, 
    -0.3901947, -0.3458748, -0.2811289, -0.2360773, -0.1851327, -0.1259696, 
    -0.1036228, -0.05598283, -0.0006443262, 0.02709007, 0.06639671, 
    0.09946978, 0.1358792, 0.1730537, 0.2119534, 0.2535388, 0.2984118, 
    0.350251, 0.4019437, 0.4446683, 0.5088611, 0.5182524, 0.5729887, 
    0.6047919, 0.6557522, 0.6897368, 0.7080798, 0.7162014, 0.7176828, 
    0.7119534, 0.7014061, 0.685114, 0.664297, 0.6396714, 0.6116439, 
    0.5821031, 0.5515203, 0.5196521, 0.4859769, 0.4514558, 0.4162998, 
    0.3810616, 0.3456938,
  -0.01905251, -0.06114197, -0.1000905, -0.1313899, -0.1557224, -0.1747978, 
    -0.1845796, -0.1857517, -0.182301, -0.1746025, -0.1643484, -0.1574966, 
    -0.153102, -0.1518002, -0.1508887, -0.1491959, -0.1469662, -0.1439224, 
    -0.1387955, -0.1321872, -0.1261978, -0.1225682, -0.1301203, -0.1456151, 
    -0.1701431, -0.2042091, -0.2382745, -0.2672946, -0.2953219, -0.323137, 
    -0.3484144, -0.3668394, -0.3773212, -0.3858333, -0.3927684, -0.3976183, 
    -0.4006133, -0.3994741, -0.3888459, -0.3717561, -0.3378367, -0.2865019, 
    -0.2107034, -0.1628189, -0.1212668, -0.06234694, -0.05674791, 
    -0.04340124, -0.05261302, -0.05163693, -0.08702111, -0.1135023, 
    -0.1479264, -0.1864845, -0.1435156, -0.194899, -0.1545344, -0.09952125, 
    -0.03964198, 0.04110348, 0.119831, 0.182331, 0.235342, 0.2601466, 
    0.2772526, 0.2852767, 0.2620183, 0.2252996, 0.1915919, 0.1862859, 
    0.2162338, 0.2464585, 0.2933497, 0.3396227, 0.3690505, 0.3742423, 
    0.3842845, 0.3751698, 0.363744, 0.3481677, 0.3448474, 0.3227769, 
    0.3017806, 0.270303, 0.2746811, 0.2491928, 0.2233137, 0.198835, 
    0.1825752, 0.1675203, 0.1549873, 0.1405015, 0.1193266, 0.09094048, 
    0.05856705, 0.02002573,
  0.178441, 0.07437205, -0.03939676, -0.1420667, -0.2257581, -0.2916437, 
    -0.3464453, -0.3653742, -0.3442479, -0.2894302, -0.2063899, -0.109808, 
    -0.002255917, 0.09339869, 0.1703681, 0.2190009, 0.22779, 0.1943748, 
    0.1308173, 0.05510104, -0.0119237, -0.04952121, -0.05196279, -0.0342055, 
    -0.03418933, -0.05124661, -0.05984026, -0.03762376, 0.006386995, 
    0.0479722, 0.06685257, 0.06478572, 0.05176473, 0.03719759, 0.02728558, 
    0.02474642, 0.02210903, 0.01672125, 0.001666546, -0.006862164, 
    -0.002614021, 0.0405345, 0.1336823, 0.1803617, 0.2094958, 0.2442939, 
    0.2165594, 0.2009181, 0.1689358, 0.1031641, 0.00337553, -0.09916341, 
    -0.1942479, -0.2526789, -0.2664812, -0.233099, -0.1907648, -0.10888, 
    -0.02647376, 0.08457756, 0.1685777, 0.2142808, 0.2396071, 0.23946, 
    0.1687731, 0.07015622, -0.03537744, -0.1090428, -0.1357517, -0.092978, 
    -0.01578021, 0.08016682, 0.1568418, 0.2195048, 0.2632065, 0.2980857, 
    0.2537999, 0.2997143, 0.3028388, 0.2538967, 0.2009997, 0.1546454, 
    0.1164127, 0.0950262, 0.09828138, 0.1361883, 0.1738997, 0.190534, 
    0.1933825, 0.2475004, 0.243969, 0.2773836, 0.2980535, 0.299746, 
    0.2909245, 0.2533593,
  0.181761, 0.07544577, -0.04527324, -0.1453221, -0.2236424, -0.276035, 
    -0.2940202, -0.2892188, -0.240016, -0.1440523, -0.02592087, 0.07442093, 
    0.1673896, 0.2483468, 0.3103094, 0.3299711, 0.3138254, 0.2479722, 
    0.1428286, 0.001520321, -0.1547463, -0.2458265, -0.2038662, -0.05077386, 
    0.1191475, 0.1716211, 0.1851141, 0.2075587, 0.1661849, 0.07547879, 
    -0.03596365, -0.1212338, -0.1401138, -0.08023441, 0.03579748, 0.1911849, 
    0.3462306, 0.4575262, 0.4794664, 0.4247303, 0.331794, 0.2125883, 
    0.2037344, 0.1814036, 0.1294827, 0.05887723, -0.03345656, -0.01182532, 
    0.0361886, -0.03054368, -0.01884115, -0.05818018, -0.104632, -0.1245376, 
    -0.1323175, -0.1161719, -0.09213221, -0.01327443, 0.06662452, 0.06574547, 
    0.09116864, 0.0573144, -0.03112943, -0.167604, -0.284987, -0.3760837, 
    -0.4559174, -0.5112395, -0.5365982, -0.52789, -0.5171809, -0.4881115, 
    -0.4344985, -0.3587985, -0.2878509, -0.2290127, -0.1709242, -0.1137464, 
    -0.07859015, -0.03466117, 0.008063436, 0.06076491, 0.07004231, 
    0.05366886, 0.05041353, 0.0438543, 0.06579429, 0.06992841, 0.0965234, 
    0.09820008, 0.1071357, 0.1807523, 0.2236397, 0.2677965, 0.2841539, 
    0.2554102,
  -0.1277279, -0.1486912, -0.1697848, -0.1396086, -0.08153605, -0.003866673, 
    0.05415726, 0.1145086, 0.3716373, 0.3635969, 0.3319569, 0.2557034, 
    0.1987368, 0.1791241, 0.1697171, 0.1134677, 0.05537701, -0.02190113, 
    -0.09237576, -0.06877577, -0.07798816, -0.06011701, 0.07756209, 
    0.3063383, 0.5623927, 0.7446353, 0.7637603, 0.6123929, 0.3507719, 
    0.07520223, -0.1224375, -0.1960546, -0.1430758, 0.01170945, 0.243464, 
    0.4952054, 0.6648831, 0.6733146, 0.5574944, 0.3494864, 0.106761, 
    -0.07022429, -0.1920834, -0.234303, -0.2490497, -0.2362075, -0.05476165, 
    -0.01703358, 0.1306548, 0.2814521, 0.5151756, 0.6312405, 0.6853094, 
    0.6173244, 0.4778387, 0.3360093, 0.1789943, 0.05202487, -0.05972643, 
    -0.1296809, -0.15805, -0.1518326, -0.1897883, -0.2404068, -0.2375911, 
    -0.2934991, -0.3413669, -0.4014093, -0.5502044, -0.6322521, -0.5761652, 
    -0.4334406, -0.4939874, -0.4441342, -0.2503841, -0.0355078, -0.07489586, 
    0.009088755, 0.08937824, 0.1338932, 0.1158431, 0.1676986, 0.2037827, 
    0.1784898, 0.1373602, 0.1352606, 0.0953517, 0.04675144, 0.002675891, 
    -0.02697891, -0.04820299, -0.04611969, -0.01696926, -0.02032213, 
    -0.04299468, -0.08785146,
  -0.05520171, -0.03593093, -0.06488609, -0.1473405, -0.1528418, -0.2094331, 
    -0.1502693, -0.0203383, -0.03000569, -0.0725193, -0.1554459, -0.2643325, 
    -0.3461848, -0.3462662, -0.2289975, -0.08065677, 0.06185484, 0.1084199, 
    0.0656805, -0.0140388, -0.006113052, 0.05521494, 0.1961818, 0.3419986, 
    0.4581935, 0.41835, 0.1862364, -0.1537209, -0.4386005, -0.5823169, 
    -0.6022718, -0.531178, -0.4075449, -0.2628996, -0.2023044, -0.1619072, 
    -0.1028576, -0.05853796, -0.1411552, -0.2035413, -0.2944758, -0.3238869, 
    -0.3479595, -0.4199634, -0.4482675, -0.5307868, -0.3495207, 0.114037, 
    0.6525784, 1.072109, 1.339362, 1.438679, 1.441869, 1.323021, 1.0961, 
    0.7872788, 0.4422593, 0.05861667, -0.3234146, -0.6106216, -0.71041, 
    -0.6832129, -0.6570244, -0.6460546, -0.5961359, -0.6017998, -0.6841404, 
    -0.8344171, -0.9028904, -0.8966242, -0.7415136, -0.5261815, -0.3676204, 
    -0.2558041, -0.07548165, 0.1009995, 0.2173406, 0.2688217, 0.2921941, 
    0.2731675, 0.2052476, 0.1822496, 0.08758804, 0.03817396, 0.06125339, 
    -0.005071484, -0.1251887, -0.2676691, -0.3252538, -0.331341, -0.3317153, 
    -0.2954199, -0.2561133, -0.2253515, -0.1342219, -0.1001074,
  -0.3818293, -0.4220473, -0.4396092, -0.423333, -0.3906833, -0.3515229, 
    -0.2929456, -0.1095145, 0.07347679, 0.09891629, 0.006354153, -0.2135025, 
    -0.3838964, -0.4191503, -0.3675878, -0.2685475, -0.1066983, 0.01828527, 
    0.06249118, 0.1079984, 0.1201079, 0.2154852, 0.2078841, 0.2190819, 
    0.2023666, 0.1128157, -0.08672822, -0.3606377, -0.5837822, -0.6273534, 
    -0.5531349, -0.4458919, -0.4054621, -0.2989353, -0.4551852, -0.493108, 
    0.02917361, -0.1336355, -0.1041436, -0.06970334, -0.1399016, -0.2393973, 
    -0.3272882, -0.4048104, -0.4085054, -0.3312919, -0.0871191, 0.3510157, 
    0.8440822, 1.256452, 1.494375, 1.510375, 1.393334, 1.171621, 0.9006252, 
    0.5384832, 0.07399751, -0.4096451, -0.8416927, -1.172194, -1.386777, 
    -1.472275, -1.425286, -1.29376, -1.130397, -1.090374, -1.168076, 
    -1.26832, -1.318076, -1.30416, -1.199717, -1.043385, -0.774147, 
    -0.4654231, -0.1793392, 0.0788478, 0.1831121, 0.2080633, 0.1867417, 
    0.1411687, 0.06328789, -0.07865545, -0.1691991, -0.2519953, -0.3995702, 
    -0.4310155, -0.4187922, -0.4233495, -0.4822036, -0.4540949, -0.395729, 
    -0.3004981, -0.2713474, -0.3220474, -0.3973404, -0.3832617,
  -1.159141, -1.221152, -1.068385, -0.7667575, -0.5346938, -0.4977636, 
    -0.4977962, -0.3650161, -0.1045181, 0.08615573, -0.001702338, -0.2191828, 
    -0.4556574, -0.6908462, -0.9116796, -1.03432, -0.9218684, -0.6999771, 
    -0.532692, -0.4687596, -0.494183, -0.5788183, -0.6879004, -0.818662, 
    -0.9078222, -0.9023208, -0.7889906, -0.6713312, -0.6192479, -0.6409603, 
    -0.686403, -0.7309016, -0.8349381, -0.9596125, -1.022357, -0.9375422, 
    -0.7017512, -0.4965752, -0.3832454, -0.4377863, -0.5670181, -0.6248957, 
    -0.622487, -0.6191665, -0.5780858, -0.4496027, -0.147552, 0.2801011, 
    0.6532781, 0.9240301, 1.014704, 0.9553777, 0.7444891, 0.4471095, 
    0.1230698, -0.2335057, -0.6271744, -0.9871516, -1.289365, -1.555902, 
    -1.832301, -1.97514, -1.908131, -1.771266, -1.591237, -1.41806, 
    -1.351865, -1.389203, -1.496234, -1.49931, -1.384775, -1.205348, 
    -1.000384, -0.6381118, -0.2535253, 0.007965654, 0.0557358, -0.05751294, 
    -0.1415787, -0.1510025, -0.2232193, -0.3759861, -0.5397882, -0.6095637, 
    -0.6024673, -0.5280206, -0.4636326, -0.470257, -0.5462499, -0.7038508, 
    -0.7233984, -0.5966895, -0.5377702, -0.6098731, -0.7743098, -0.9869888,
  -1.223431, -1.013535, -0.7331314, -0.5309342, -0.5416763, -0.6599219, 
    -0.6529231, -0.4857356, -0.2970151, -0.3319435, -0.6156838, -0.9126724, 
    -1.107806, -1.277044, -1.491774, -1.597031, -1.441872, -1.131504, 
    -0.9794854, -1.010166, -1.085963, -1.230706, -1.423317, -1.584873, 
    -1.624473, -1.401344, -1.069525, -0.7789483, -0.6812108, -0.7412367, 
    -0.8715753, -1.039853, -1.184791, -1.275954, -1.247373, -1.046006, 
    -0.7468031, -0.5887791, -0.6559666, -0.8490004, -0.9743913, -0.9141537, 
    -0.782155, -0.7759376, -0.7986264, -0.6524023, -0.331325, -0.04133475, 
    0.08613932, 0.07331383, 0.01885414, -0.05577141, -0.1269466, -0.2253514, 
    -0.4175389, -0.7834081, -1.208766, -1.505413, -1.692848, -1.937249, 
    -2.210768, -2.351296, -2.293744, -2.115716, -1.934352, -1.708376, 
    -1.583864, -1.600791, -1.679306, -1.709922, -1.6032, -1.393695, 
    -1.158685, -0.9009374, -0.6886978, -0.5631118, -0.5479262, -0.6119074, 
    -0.6143161, -0.4908788, -0.3127701, -0.3452571, -0.4844498, -0.6546646, 
    -0.7513933, -0.7362564, -0.7397395, -0.8937107, -1.171624, -1.383685, 
    -1.318092, -1.090618, -0.9782649, -1.089479, -1.214642, -1.268239,
  -1.138177, -1.020469, -0.9466895, -0.9229425, -0.9497328, -0.9016536, 
    -0.7402929, -0.5974542, -0.6110609, -0.7862403, -0.9682713, -1.201702, 
    -1.419053, -1.572487, -1.634645, -1.517653, -1.295631, -1.142816, 
    -1.135329, -1.218483, -1.240993, -1.28095, -1.431504, -1.540146, 
    -1.477858, -1.248431, -0.9785251, -0.7189713, -0.5986098, -0.7401136, 
    -0.9827569, -1.139837, -1.207138, -1.178948, -1.072242, -0.9265066, 
    -0.7753677, -0.7052993, -0.7577569, -0.8671484, -0.9117448, -0.9372166, 
    -1.011045, -1.060915, -1.030055, -0.9312434, -0.8002049, -0.7135024, 
    -0.6086683, -0.4926691, -0.4135025, -0.3974379, -0.345729, -0.3388771, 
    -0.5369402, -0.9557225, -1.397536, -1.620517, -1.697031, -1.875611, 
    -2.123366, -2.21928, -2.152191, -2.045517, -1.934173, -1.779844, 
    -1.677077, -1.743841, -1.835882, -1.774, -1.615162, -1.395859, -1.184938, 
    -1.081048, -1.04, -0.9584897, -0.8226168, -0.7059343, -0.5763121, 
    -0.3883559, -0.2834243, -0.3698827, -0.6484146, -0.8641046, -0.9662531, 
    -1.066612, -1.196071, -1.427777, -1.639268, -1.629941, -1.339235, 
    -1.073398, -1.090863, -1.200498, -1.242034, -1.222633,
  -1.044622, -0.9161229, -0.781992, -0.6004, -0.4413507, -0.3182387, 
    -0.2332451, -0.2614844, -0.4094338, -0.5774021, -0.7281837, -0.9103777, 
    -1.085784, -1.095892, -0.9413834, -0.8024514, -0.7436624, -0.7550223, 
    -0.8276298, -0.9249444, -0.9135838, -0.8862075, -0.8790947, -0.8438572, 
    -0.7183527, -0.6146579, -0.54319, -0.4469657, -0.3760023, -0.4344494, 
    -0.5960381, -0.7538347, -0.7980895, -0.7692156, -0.80779, -0.9218524, 
    -0.9832127, -0.9420342, -0.8673761, -0.8444428, -0.8266532, -0.8430433, 
    -0.9305272, -0.9237725, -0.832464, -0.826865, -0.8585382, -0.7840103, 
    -0.5536716, -0.356585, -0.2812107, -0.2112234, -0.1579032, -0.2923269, 
    -0.6661553, -1.124179, -1.363454, -1.46417, -1.602581, -1.819932, 
    -1.966563, -1.923268, -1.817084, -1.710963, -1.594997, -1.483326, 
    -1.487542, -1.496185, -1.446364, -1.332236, -1.210719, -1.066091, 
    -0.9262791, -0.8210385, -0.7210376, -0.630722, -0.4985766, -0.2318778, 
    0.1089097, 0.1484768, -0.006080508, -0.2213309, -0.4882417, -0.6842219, 
    -0.7915133, -0.8881445, -1.040098, -1.182041, -1.286598, -1.211826, 
    -1.041009, -0.940179, -0.9477794, -0.9782318, -1.040374, -1.0997,
  -0.346559, -0.1814711, -0.03337526, 0.1153064, 0.2217684, 0.2659252, 
    0.3515043, 0.3761137, 0.2492588, 0.1231513, -0.008375168, -0.1819267, 
    -0.2945244, -0.3090589, -0.3198657, -0.4019945, -0.5278416, -0.621217, 
    -0.7072518, -0.7559338, -0.6374283, -0.4930433, -0.3949964, -0.3319917, 
    -0.2702081, -0.2148857, -0.09421515, 0.01913166, 0.04722404, 0.04637742, 
    0.02901077, -0.03540993, -0.1651304, -0.3038023, -0.424196, -0.4531019, 
    -0.4030368, -0.3280041, -0.2865164, -0.2836683, -0.270973, -0.2385998, 
    -0.2875257, -0.3689873, -0.3500745, -0.297812, -0.2653577, -0.1681571, 
    -0.01976848, 0.03172874, -0.01412082, -0.03275681, -0.1195407, 
    -0.3786063, -0.7535577, -1.093824, -1.305072, -1.383929, -1.488226, 
    -1.540277, -1.372308, -1.109417, -1.03777, -1.018613, -1.000482, 
    -1.056781, -1.017995, -0.8405693, -0.7546482, -0.7367606, -0.6197686, 
    -0.4502046, -0.3000908, -0.1573007, 0.06628323, 0.2909904, 0.4769599, 
    0.6945386, 0.7535875, 0.4857652, 0.08244491, 0.06937551, 0.07243538, 
    -0.1371677, -0.3819268, -0.4939387, -0.6125908, -0.7774835, -0.8892673, 
    -0.9063246, -0.8356215, -0.7393651, -0.6143975, -0.5752535, -0.5890884, 
    -0.5040295,
  0.4296293, 0.5620999, 0.8152254, 0.9706776, 0.9677804, 1.044961, 1.16656, 
    1.130867, 0.9238025, 0.6820706, 0.4068103, 0.1024485, -0.06389284, 
    -0.2127047, -0.3605399, -0.4622488, -0.5197036, -0.5415132, -0.5776951, 
    -0.5347915, -0.3080986, -0.1448987, -0.1635022, -0.08671188, 0.1004462, 
    0.2878976, 0.4765532, 0.5949292, 0.6506093, 0.7279532, 0.7962472, 
    0.7472887, 0.5440986, 0.3588285, 0.2916083, 0.2823474, 0.2897692, 
    0.3588448, 0.5042546, 0.4807682, 0.2390528, 0.1423242, 0.1519761, 
    0.07673204, 0.1441801, 0.3099194, 0.286335, 0.2442615, 0.1214423, 
    0.01695037, -0.07606745, -0.1672132, -0.2710707, -0.4377372, -0.6082773, 
    -0.7885182, -0.9345632, -0.8983326, -0.762151, -0.6538827, -0.4320896, 
    -0.2860446, -0.4064221, -0.5168231, -0.5480731, -0.5873797, -0.4423921, 
    -0.221282, -0.1512132, -0.03225183, 0.1121655, 0.2780836, 0.5086172, 
    0.7191963, 0.9815984, 1.519814, 1.909561, 1.507494, 0.7413639, 
    0.05689138, -0.1186457, 0.3448472, 0.4936428, 0.1875718, -0.07273078, 
    -0.1933038, -0.3151951, -0.5099542, -0.5840263, -0.5011814, -0.4372327, 
    -0.3576756, -0.1897719, -0.10971, 0.02049851, 0.2863185,
  0.7400459, 1.0496, 1.314427, 1.318936, 1.310749, 1.300788, 1.210912, 
    1.024958, 0.7337143, 0.3110582, -0.1057224, -0.3223891, -0.323561, 
    -0.3137468, -0.2768161, -0.2397882, -0.2938738, -0.3509372, -0.2813574, 
    -0.1288507, 0.0782131, 0.269196, 0.4210677, 0.6021875, 0.7847723, 
    0.9426985, 1.083975, 1.220694, 1.396442, 1.429222, 1.311416, 1.075951, 
    0.7520574, 0.6004137, 0.5364813, 0.5377671, 0.7052636, 0.9333237, 
    1.053408, 0.7642645, 0.2299708, 0.0315007, 0.3311101, 0.5944564, 
    0.7960027, 0.8865952, 0.6734278, 0.3950911, 0.2035872, 0.002203941, 
    -0.209645, -0.3197687, -0.3312757, -0.437542, -0.6068618, -0.5831149, 
    -0.3654878, -0.02194953, 0.1875725, 0.1431875, 0.1736722, 0.1514392, 
    0.04999065, 0.07025433, 0.05139017, 0.1095121, 0.3351631, 0.3655832, 
    0.3163643, 0.5391343, 0.7368556, 0.8400943, 1.099502, 1.314932, 1.490843, 
    2.150625, 2.334333, 1.070417, -0.05479485, -0.4168065, 0.02476233, 
    0.2848374, 0.2590885, 0.2055894, 0.03413749, -0.179697, -0.3858006, 
    -0.441855, -0.3419855, -0.2110934, -0.1534927, -0.08861613, 0.06566429, 
    0.2066636, 0.3311753, 0.5442613,
  1.253132, 1.446735, 1.480508, 1.536172, 1.681713, 1.424584, 1.109854, 
    0.7481838, 0.1118557, -0.2559342, 0.0003484488, 0.3174708, 0.2581608, 
    0.1177963, 0.1528548, 0.08379555, -0.1922459, -0.3596776, -0.1912695, 
    0.1506088, 0.3968002, 0.6437241, 0.8721908, 0.901569, 0.9688869, 
    1.213369, 1.471442, 1.669424, 1.773151, 1.687686, 1.471459, 1.001732, 
    0.5320376, 0.5115461, 0.6085024, 0.7773178, 0.9798572, 1.074323, 
    0.8284084, 0.2724839, -0.0170832, 0.2355859, 0.5923895, 0.9106673, 
    1.121377, 0.8864813, 0.2690171, -0.1008723, -0.1767514, -0.2683692, 
    -0.3845152, -0.5608009, -0.656504, -0.5982357, -0.483099, -0.173431, 
    0.3211979, 0.6380761, 0.5612532, 0.3032616, 0.2980859, 0.3214422, 
    0.3474026, 0.4344306, 0.3981838, 0.4503485, 0.5661851, 0.6193261, 
    0.6866114, 0.8204495, 0.9982651, 1.115973, 1.135602, 1.253653, 1.55336, 
    1.798818, 1.14299, 0.24265, -0.2715265, -0.09893554, 0.2269598, 
    0.1133856, 0.175739, 0.3973863, 0.1472073, -0.1756606, -0.2265558, 
    -0.1344333, -0.1223403, -0.2113378, -0.133831, -0.004778385, 0.1899154, 
    0.4689518, 0.7117417, 0.9769273,
  1.049046, 1.107054, 1.248704, 1.617926, 1.448133, 0.8745837, 0.4698637, 
    0.1918522, -0.1145441, 0.3077542, 0.9264389, 0.806354, 0.2231998, 
    -0.08999991, -0.05053037, -0.2705011, -0.5127538, -0.3080663, 0.1029038, 
    0.5071681, 0.6840235, 0.8381415, 0.9502181, 0.9769924, 1.096719, 
    1.314118, 1.496491, 1.611156, 1.622436, 1.527137, 1.175185, 0.5463121, 
    0.1720117, 0.4501859, 0.5793198, 0.7203355, 0.7228909, 0.5114489, 
    0.1583238, -0.2904883, 0.1374251, 0.8054754, 0.8578191, 0.9406966, 
    1.013841, 0.6087468, -0.131211, -0.423903, -0.3813085, -0.4542251, 
    -0.4613052, -0.5873632, -0.704046, -0.3849705, -0.02051744, 0.2703843, 
    0.4972721, 0.5090561, 0.3486395, 0.2234278, 0.4476302, 0.6292382, 
    0.5952378, 0.5106348, 0.5020901, 0.5972073, 0.590957, 0.6520247, 
    0.8528225, 0.8801987, 0.882282, 0.9860092, 0.9357163, 0.952611, 1.018919, 
    0.5316458, -0.4498978, -0.4212985, -0.001279235, 0.1285875, 0.1364487, 
    0.03088229, 0.2290918, 0.4218003, 0.06338573, -0.04242516, 0.02110052, 
    -0.06701803, -0.2001723, -0.306455, -0.05360675, 0.2543036, 0.4113021, 
    0.6248276, 0.8591539, 0.9985254,
  0.7098539, 0.8160553, 0.8995657, 0.8340383, 0.5145884, 0.1434803, 
    -0.1709406, -0.126686, 0.2955633, 1.110749, 1.284658, 0.6585362, 
    -0.2036231, -0.829681, -0.6547135, -0.3274347, -0.333164, -0.2372167, 
    0.006403208, 0.283161, 0.580459, 0.7543524, 0.7301011, 0.7289617, 
    0.8467348, 0.9434969, 1.089054, 1.166493, 0.9990945, 0.6937385, 0.222075, 
    -0.1597753, -0.119069, 0.3348209, 0.3556541, 0.4391832, 0.4058824, 
    0.2595932, -0.05489242, -0.3568618, 0.3288152, 0.8948632, 0.90056, 
    0.832217, 0.6425686, 0.1793525, -0.5995214, -0.8081964, -0.5514744, 
    -0.4100032, -0.3789647, -0.6641698, -0.8061619, -0.3574966, -0.06443021, 
    0.04688165, 0.190713, 0.235407, 0.4091212, 0.6022038, 0.7721421, 
    0.7891668, 0.6254461, 0.5548081, 0.5429916, 0.6028224, 0.6459864, 
    0.7631252, 0.8502182, 0.7716864, 0.6332912, 0.5904202, 0.5674386, 
    0.392633, 0.1793022, -0.2389097, -0.6764431, -0.07172179, 0.178913, 
    -0.1710383, -0.2423111, -0.1421157, 0.1037013, 0.1732488, 0.05681002, 
    0.06109118, -0.196722, -0.3811455, -0.2847426, -0.09756839, 0.1315659, 
    0.3379949, 0.4934963, 0.6117578, 0.7544175, 0.7640204,
  0.3280182, 0.2695203, 0.07459736, 0.003780365, -0.01633406, -0.2715591, 
    -0.3403254, 0.07555997, 0.3616278, 0.6534574, 0.9562573, 0.5421295, 
    -0.2632744, -0.963177, -0.7205826, 0.1455634, 0.08763683, -0.3692479, 
    -0.2854102, 0.0993228, 0.5494534, 0.7661854, 0.6550851, 0.6083395, 
    0.6252353, 0.6601639, 0.7148185, 0.5353894, 0.123003, -0.2697377, 
    -0.456471, -0.3337009, -0.09016266, 0.2430406, 0.2063707, 0.1940498, 
    0.1355376, -0.1216893, -0.4040785, -0.2331639, 0.5905504, 0.7841537, 
    0.6983464, 0.3812237, 0.1639881, -0.2024021, -0.9542413, -0.886191, 
    -0.5419529, -0.2774024, -0.3188249, -0.6665299, -0.6891048, -0.2506282, 
    -0.03597957, 0.009397954, 0.2798733, 0.5118557, 0.7613837, 0.8279037, 
    0.8545153, 0.7988837, 0.6399807, 0.6722072, 0.6701565, 0.6369531, 
    0.6212792, 0.6986231, 0.6277899, 0.4961169, 0.4297426, 0.3573799, 
    0.3165436, 0.09092331, -0.07086086, -0.1446896, -0.3254976, -0.01462567, 
    -0.002809137, -0.3809345, -0.2992284, -0.02343088, 0.2453352, 0.1658269, 
    0.215827, 0.1228583, -0.3116136, -0.2170506, 0.1129948, 0.2418523, 
    0.2947495, 0.3507879, 0.4094143, 0.4330959, 0.4446032, 0.3714426,
  0.1060777, -0.1356397, -0.3239861, -0.1011324, -0.06539053, -0.4143163, 
    -0.2027767, 0.3058986, 0.2161359, 0.3006904, 0.8914621, 0.3838446, 
    -0.3636327, -0.5158462, -0.4346452, 0.5180893, 0.4346094, -0.4719498, 
    -0.4868749, 0.05490553, 0.5749743, 0.7091539, 0.542129, 0.3553617, 
    0.242846, 0.176228, -0.01921558, -0.1715102, -0.3785415, -0.5475855, 
    -0.4163015, -0.2369562, -0.1086359, 0.1199938, -0.005006313, -0.1460218, 
    -0.01529264, 0.01292968, 0.06319025, 0.392715, 0.5351955, 0.3547432, 
    0.1407948, -0.4865327, -0.6332774, -0.7564547, -1.235394, -1.01928, 
    -0.7742122, -0.4160742, -0.269134, -0.5104426, -0.582513, -0.3460546, 
    -0.01695293, 0.07567394, 0.4005276, 0.7474512, 0.8708073, 0.7964423, 
    0.7833237, 0.8079003, 0.7037013, 0.6635482, 0.6255109, 0.6637762, 
    0.6143786, 0.60043, 0.5232327, 0.3629138, 0.2995348, 0.2578201, 
    0.1574931, -0.09224653, -0.146152, 0.04142857, 0.1409736, 0.1068914, 
    -0.266253, -0.2211362, 0.07269543, 0.2124251, 0.3093002, 0.2748438, 
    0.4106023, 0.1207746, -0.2443452, 0.09753251, 0.3053125, 0.3130112, 
    0.3023828, 0.3246486, 0.3204007, 0.3054268, 0.2463772, 0.1298742,
  -0.08908796, -0.2431741, -0.2965589, -0.02217758, 0.0132553, -0.08235025, 
    0.3249417, 0.3227443, 0.06058604, 0.1333561, 0.3800684, 0.127269, 
    -0.2968682, -0.2807551, -0.3338146, 0.5262436, 0.4929591, -0.5931411, 
    -0.5888119, 0.1420311, 0.70152, 0.5926173, 0.2052803, 0.005817413, 
    -0.01914954, -0.04255509, -0.3408296, -0.3038013, -0.3326099, -0.4265881, 
    -0.3677994, -0.1920344, -0.09577787, -0.1266208, -0.4417254, -0.381927, 
    -0.1609472, -0.3356867, -0.1701269, -0.1968684, -0.3112237, -0.2169369, 
    -0.5932877, -1.164186, -1.181178, -1.035426, -1.118158, -0.9612238, 
    -0.7306086, -0.1902928, 0.07448579, -0.2896418, -0.5822525, -0.2888931, 
    0.1574936, 0.2382065, 0.5662175, 0.8655015, 0.8728744, 0.8708236, 
    0.8006412, 0.7520084, 0.7527245, 0.7780665, 0.7107813, 0.6366441, 
    0.5604072, 0.4887602, 0.4051499, 0.3448472, 0.3087633, 0.2547433, 
    0.1187081, 0.03620529, 0.1490774, 0.1843648, 0.3191799, 0.2231023, 
    -0.1740983, -0.08446634, 0.2133366, 0.2271063, 0.1587794, 0.07959628, 
    0.1111068, -0.1994565, -0.1003027, 0.2445378, 0.3224676, 0.3881902, 
    0.2900783, 0.1804919, 0.1232328, 0.08714867, 0.03739309, -0.03560519,
  -0.02709222, -0.098984, -0.163779, -0.02116853, 0.1303615, 0.1596421, 
    0.3185449, 0.07442057, 0.1686427, 0.2921453, 0.2674383, 0.1760974, 
    -0.07435846, 0.04551446, 0.1725327, 0.4850652, 0.194424, -0.4293877, 
    -0.1272232, 0.3112534, 0.6341375, 0.3654687, 0.09064764, 0.003294468, 
    -0.1602311, -0.1969985, -0.4162368, -0.3502212, -0.2756771, -0.2567642, 
    -0.2272883, 0.08902013, 0.3213444, -0.1381605, -0.8114517, -0.6580177, 
    -0.4952898, -0.7384372, -0.5493096, -0.9678482, -0.921901, -0.6626236, 
    -1.162982, -1.140863, -1.213421, -1.009238, -0.6404882, -0.48305, 
    -0.2917742, 0.009430408, 0.3442286, 0.009056091, -0.2973893, 0.02487645, 
    0.2256902, 0.2264064, 0.4578354, 0.6636135, 0.5815822, 0.5749088, 
    0.5911849, 0.6506411, 0.6641669, 0.6338936, 0.5752344, 0.4473052, 
    0.4028063, 0.3739488, 0.3060777, 0.32862, 0.2930901, 0.245466, 0.1335192, 
    0.05515003, 0.001211643, 0.1366605, 0.03635105, 0.1974024, 0.0530175, 
    0.23806, 0.1499578, 0.09250337, 0.1584702, 0.09819996, 0.04068047, 
    -0.005706251, 0.1867091, 0.2949285, 0.2702052, 0.1889387, 0.1071682, 
    0.03251004, 0.08605838, 0.08249402, 0.01727581, 0.01307702,
  -0.2566175, -0.3197682, -0.1662857, 0.02642266, 0.08384453, 0.1107325, 
    0.07199538, -0.006113291, 0.09251964, -0.02662095, 0.07412755, 0.2535224, 
    0.01789427, 0.2268457, 0.2688543, 0.1803287, -0.01692033, -0.1880143, 
    -0.01241201, 0.116901, 0.3649969, 0.1980372, 0.06397149, -0.01600899, 
    -0.2367935, -0.1770767, -0.1769628, -0.2126073, -0.1785741, -0.06068671, 
    0.07988945, 0.2429103, 0.2405015, -0.1448987, -0.8971125, -0.6610775, 
    -0.2576592, -0.5225356, -0.4327245, -0.8815038, -0.9682063, -0.7593683, 
    -0.957562, -0.520355, -0.5408299, -0.4458432, -0.2142187, -0.2280697, 
    -0.1662533, 0.02132821, 0.244489, -0.06760424, -0.2674088, 0.01170909, 
    0.2184799, 0.3587306, 0.3656642, 0.3726792, 0.3484931, 0.3557521, 
    0.3224022, 0.3438865, 0.4323148, 0.4689195, 0.369359, 0.3265531, 
    0.2779691, 0.2809966, 0.3325915, 0.3242581, 0.1605053, 0.06301141, 
    0.05606151, 0.02792025, -0.09231091, 0.02995456, 0.1498438, 0.09976238, 
    0.131631, 0.1343979, 0.0912827, 0.1233139, 0.1566961, 0.1073797, 
    0.04100585, 0.1029526, 0.1269923, 0.1177801, 0.2381901, 0.1297265, 
    0.1469957, 0.003620028, -0.02273083, -0.1039808, -0.1719332, -0.196249,
  -0.4325128, -0.4057389, -0.1655697, 0.03011715, 0.04208022, -0.002971858, 
    0.005589306, -0.03008777, -0.1067153, -0.3055108, -0.003248632, 
    0.3707592, 0.2328672, 0.254564, 0.2513578, 0.2191473, 0.1700588, 
    0.1484931, 0.2486883, 0.4095282, 0.4566474, 0.272614, 0.142422, 
    0.02264661, -0.07305664, 0.06634778, 0.1818262, 0.08076836, 0.03960626, 
    0.1926497, 0.4596582, 0.3036362, -0.1520116, -0.3373137, -0.7917085, 
    -0.3675715, 0.06517589, -0.08340807, -0.03059232, -0.0708431, -0.1857674, 
    -0.4698825, -0.815309, -0.7038182, -0.6194756, -0.6723077, -0.6199477, 
    -0.5859469, -0.5869074, -0.3721611, -0.3920177, -0.5759698, -0.4705502, 
    -0.2646582, -0.1245542, -0.04042339, -0.004729748, 0.02691096, 
    0.01511079, 0.01662448, -0.02596992, -0.00590156, 0.0977931, 0.2331284, 
    0.1914455, 0.238418, 0.1993717, 0.1838772, 0.1475002, 0.005817413, 
    -0.05442023, -0.01350236, -0.08926725, -0.2666762, -0.3240329, 
    -0.004762232, 0.01162773, -0.05033515, 0.030215, 0.00261081, 0.08926439, 
    0.1471583, 0.1155014, 0.2487534, 0.1395737, -0.122812, -0.1362076, 
    -0.0202733, 0.05124363, 0.004091948, 0.05887705, -0.02680004, 0.01063454, 
    -0.1701921, -0.3397557, -0.4213802,
  -0.1595799, -0.1835873, -0.104746, 0.06232762, 0.1372464, 0.01807304, 
    -0.004664581, -0.06490221, -0.04776354, 0.1028387, 0.3428777, 0.2773013, 
    0.1228421, 0.1148486, 0.397419, 0.4885654, 0.4758368, 0.6475008, 
    0.5744373, 0.527692, 0.4728745, 0.3714583, 0.2290107, 0.1186426, 
    0.06647789, 0.05778664, 0.1266667, 0.001585424, -0.1018975, -0.004224777, 
    0.07337904, -0.004192591, -0.02343094, 0.2583222, -0.1547627, -0.1420019, 
    -0.03988594, 0.08161467, 0.4228909, 0.4418857, 0.01052189, -0.276686, 
    -0.4058526, -0.4605889, -0.4344006, -0.4601007, -0.3884692, -0.3304288, 
    -0.3831143, -0.295387, -0.2819107, -0.2151299, -0.1688082, -0.2204523, 
    -0.2089446, -0.2457128, -0.2543226, -0.2627863, -0.3211521, -0.3629978, 
    -0.3594662, -0.2182064, -0.1910906, -0.1053321, -0.004339099, 0.05747736, 
    -0.004973888, 0.118838, 0.1975164, 0.1108302, 0.06535494, 0.1090236, 
    -0.01285148, -0.2379328, -0.3249771, -0.1011327, 0.004189581, 0.01208347, 
    0.02762709, 0.0678452, 0.0897039, 0.0735743, -0.09122086, -0.3561456, 
    -0.1447685, -0.3923924, -0.2744722, -0.07126629, -0.04486656, 
    -0.02839512, 0.009170055, -0.03736314, -0.02175432, -0.1646256, 
    -0.1967545, -0.1808365,
  0.1127999, 0.09183609, 0.2000227, 0.09499362, -0.00554347, -0.05914047, 
    0.01673841, -0.03959297, -0.03902331, 0.06078138, 0.01231131, 
    -0.03145492, 0.09294295, 0.0344615, 0.2376842, 0.5115457, 0.6086657, 
    0.7925203, 0.7423415, 0.7355537, 0.7144922, 0.5514065, 0.3435781, 
    0.0831449, 0.1116439, 0.1485093, 0.1076889, -0.1136002, -0.3004498, 
    -0.3033624, -0.1194761, 0.00617528, 0.03963864, 0.4045639, 0.1243067, 
    0.06131887, -0.09055305, 0.05493832, 0.03742528, 0.06540442, 0.006143093, 
    -0.05354071, -0.04867458, -0.008619308, 0.1063871, 0.2774813, 0.365144, 
    0.4450264, 0.5127027, 0.5301342, 0.5322177, 0.4468336, 0.3837798, 
    0.3292387, 0.1651108, 0.02202821, -0.1347101, -0.251491, -0.3112566, 
    -0.3570412, -0.4442155, -0.4630629, -0.4377865, -0.4485935, -0.4721287, 
    -0.375563, -0.2389419, -0.08788398, -0.06228179, 7.176399e-005, 
    0.1034573, 0.1637272, 0.07736668, -0.008684993, -0.04535484, -0.06125638, 
    0.09614923, 0.4103256, 0.3087955, 0.2842677, 0.2334383, -0.04530585, 
    -0.1760186, -0.2648711, -0.1085868, -0.0254488, 0.07972693, 0.0946362, 
    0.1040602, 0.08304715, 0.04564452, 0.004531384, -0.04605456, 0.04901379, 
    0.1847724, 0.2098539,
  -0.06125653, -0.2547622, -0.04017895, -0.2480891, -0.5955337, -0.5767186, 
    -0.2992121, -0.2436948, -0.2803483, -0.1430109, -0.04226226, -0.06482086, 
    0.02287447, 0.02044773, -0.1431103, 0.2870994, 0.5047102, 0.6026106, 
    0.6709385, 0.5893135, 0.5659572, 0.4863346, 0.6926346, 0.3468499, 
    0.1061759, 0.03807664, 0.01716158, -0.05542958, -0.4499116, -0.6191683, 
    -0.3740335, -0.0591079, 0.01278329, 0.3152084, 0.229043, 0.3754458, 
    0.2302804, 0.2548897, 0.2584701, 0.3418036, 0.3080797, 0.1576896, 
    0.05511761, 0.08460951, 0.08109379, 0.1090565, 0.1094799, 0.1727772, 
    0.3003817, 0.3478746, 0.4513412, 0.5189197, 0.6150949, 0.6677809, 
    0.5271232, 0.3877513, 0.2504957, 0.1519606, -0.04231095, -0.2395763, 
    -0.3630791, -0.4489515, -0.417327, -0.4217706, -0.5172133, -0.499375, 
    -0.3525002, -0.1474057, -0.03059244, 0.05173159, 0.1281314, 0.3209212, 
    0.5168688, 0.3266829, 0.3808661, 0.1517319, 0.3876858, 0.5660062, 
    0.4290926, -0.1162856, -0.1034107, 0.03583097, 0.5929763, 0.4433489, 
    0.3467185, 0.2874084, 0.2477283, 0.1726136, 0.2348375, 0.2486892, 
    0.1900947, 0.07443702, -0.1168879, -0.07893229, 0.05775404, 0.04352885,
  0.03280282, -0.2218195, -0.4319919, -0.4722912, -0.8072197, -0.8870538, 
    -0.5356541, -0.430999, -0.3527923, -0.09260428, 0.1131902, 0.06846367, 
    -0.05272773, -0.07478142, -0.325841, -0.1183219, 0.1907768, 0.4232974, 
    0.6600323, 0.69628, 0.9164779, 0.5699286, 0.8545809, 0.6540928, 0.294034, 
    -0.1510832, -0.1056409, -0.004160024, -0.2618259, -0.6340933, -0.8004994, 
    -0.4765553, -0.4639411, -0.0127697, 0.04782629, 0.2366271, 0.2437243, 
    0.149323, 0.181859, 0.1855698, 0.177855, 0.2378483, 0.221817, 0.1451883, 
    0.1070542, 0.09050179, 0.04502535, 0.02700806, 0.06537056, 0.1307516, 
    0.09072876, 0.08236265, 0.06636381, 0.1839738, 0.363678, 0.3933816, 
    0.3583879, 0.2539291, 0.1768293, 0.02098656, -0.195859, -0.2956963, 
    -0.390358, -0.3887463, -0.4784594, -0.6560965, -0.6059663, -0.3682383, 
    -0.156227, 0.07206082, 0.1283922, 0.2351143, 0.8759508, 0.7555885, 
    0.05669594, -0.04017878, -0.1892998, -0.2969813, -0.293906, -0.1339285, 
    0.2269769, 0.3297112, 0.3224514, 0.2381904, 0.2074113, 0.1433334, 
    0.1617255, 0.1825256, 0.2352924, 0.3586326, 0.5457745, 0.5555413, 
    0.3794173, 0.1982651, 0.123086, 0.1368717,
  0.2067132, 0.08683944, -0.08845282, -0.1206963, -0.3146582, -0.6419525, 
    -0.6528254, -0.4973564, -0.3873806, -0.3854756, -0.1453224, 0.02730155, 
    -0.1874444, -0.3566013, -0.4151461, -0.3167415, -0.1437435, 0.1130762, 
    0.3019595, 0.314476, 0.5159896, 0.735993, 1.09353, 0.7612379, 0.592325, 
    0.1838942, -0.1887465, -0.4238214, -0.5004491, -0.810475, -0.9835699, 
    -0.494524, -0.7623954, -0.5767021, -0.3936942, -0.258863, -0.1283131, 
    -0.1750736, -0.1459732, -0.1449962, -0.104583, -0.1142349, -0.01872683, 
    0.02967787, 0.01960325, 0.02805066, 0.04553103, 0.04992533, 0.01013041, 
    0.09411478, 0.07141018, 0.05288744, -0.009758472, -0.03697205, 
    -0.02551365, 0.07279301, 0.261986, 0.2149971, 0.149909, 0.1115794, 
    -0.01298189, -0.1168394, -0.2219987, -0.2080827, -0.2254982, -0.3344502, 
    -0.4646082, -0.6224704, -0.5233496, 0.0413478, 0.5468492, 0.5348866, 
    0.3974354, -0.07730436, -0.5193467, -0.520582, -0.3646252, -0.1465102, 
    0.1629791, 0.4098535, 0.3607814, 0.1647694, 0.07386804, 0.05056071, 
    0.02261472, 0.06439543, 0.05202484, 0.08340502, 0.150218, 0.2571664, 
    0.4123096, 0.540565, 0.4540436, 0.1983466, 0.2545483, 0.3058829,
  0.3248284, 0.1455636, 0.03125668, 0.1169994, -0.02178669, -0.4757578, 
    -0.7988045, -0.7028415, -0.5477486, -0.4303169, -0.4452889, -0.06127274, 
    -0.1995376, -0.6438246, -0.6226009, -0.410605, -0.2827239, -0.05044937, 
    0.3285222, 0.1835504, 0.1409085, 0.8456122, 1.37932, 0.9100491, 
    0.8162013, 0.5698957, -0.03965807, -0.5349869, -0.9408625, -1.455625, 
    -1.482562, -0.4599867, -0.5491304, -0.8467541, -0.8706965, -0.7388766, 
    -0.5471444, -0.4325285, -0.369801, -0.4267023, -0.4461682, -0.4514737, 
    -0.2718186, -0.1561291, -0.182008, -0.1636651, -0.06914997, -0.04693317, 
    -0.1439059, -0.1311781, -0.09623289, -0.06861305, 0.02806711, 0.05261087, 
    0.03490329, 0.1133537, 0.1897209, 0.2476311, 0.2565341, 0.2419505, 
    0.1241443, -0.05647135, -0.190733, -0.3080831, -0.2442331, -0.1876569, 
    -0.4210877, -0.6927178, -0.4677013, -0.1090916, -0.1388121, -0.07131493, 
    -0.1988865, -0.8108819, -0.6399181, -0.3128679, -0.09533841, 0.1622788, 
    0.2803125, 0.3200426, 0.3334538, 0.3740304, 0.2342842, 0.02676463, 
    -0.1667249, -0.1496351, -0.08804607, -0.06107712, -0.04091215, 
    -0.00603199, 0.1218152, 0.2159719, 0.1634347, 0.1774807, 0.1680574, 
    0.2759676,
  0.6165434, 0.3666406, -0.1324801, -0.2932706, -0.2549572, -0.5285578, 
    -0.9597752, -1.016953, -1.032968, -0.734271, -0.4728947, 0.06857741, 
    0.102855, -0.5553157, -0.7599709, -0.5101985, -0.7126398, -0.6229258, 
    0.1400459, 0.3666732, 0.1131904, 0.3378322, 0.6572168, 0.8467516, 
    0.6568426, 0.1200425, 0.1238022, 0.1054914, -0.3751398, -1.25346, 
    -1.416709, -0.6234636, -0.4789319, -0.8641046, -1.09612, -1.024749, 
    -0.8472588, -0.700465, -0.5964124, -0.5191174, -0.4642508, -0.4682224, 
    -0.4778415, -0.4029882, -0.312884, -0.2896906, -0.188014, -0.1234465, 
    -0.08324528, -0.0605886, -0.09349895, -0.1815848, -0.09164357, 
    -0.01887321, -0.05949855, -0.02310514, 0.02699244, 0.2006904, 0.3236072, 
    0.3489325, 0.1971912, 0.04004645, -0.08576798, -0.2827573, -0.266253, 
    -0.2187448, -0.1164823, -0.1298759, -0.05993789, -0.08031562, -0.3102797, 
    -0.2184178, -0.2342058, -0.7198013, -0.5826755, -0.2910581, -0.088893, 
    0.1626368, 0.334284, 0.4141016, 0.3983626, 0.3861232, 0.2164944, 
    0.06260407, -0.07136393, -0.1418067, -0.117197, -0.082757, -0.03496981, 
    -0.04743814, 0.02149057, 0.1295314, 0.109838, 0.2080472, 0.0913806, 
    0.2320869,
  -0.07974577, 0.437051, 0.2550846, -0.1853123, -0.2822523, -0.5118259, 
    -0.9333106, -1.109417, -1.328167, -1.017505, -0.6431241, -0.4310158, 
    -0.2345311, -0.4648045, -0.5187762, -0.4874771, -0.9633723, -0.6795671, 
    -0.07899714, 0.02020526, 0.1749091, 0.2900455, 0.1030016, 0.3488997, 
    0.03195643, -0.4423925, -0.1160904, 0.1394436, -0.2352471, -0.4796644, 
    -0.806113, -0.7778094, -0.342392, -0.2941337, -0.3341892, -0.4506279, 
    -0.6223077, -0.632122, -0.6741307, -0.6669041, -0.603281, -0.5334243, 
    -0.5074641, -0.4941342, -0.4474542, -0.4366636, -0.3151625, -0.2474868, 
    -0.2300715, -0.2055925, -0.108506, -0.06250978, -0.09068334, -0.1218033, 
    -0.1347754, -0.001767457, 0.1341375, 0.1670314, 0.104157, 0.1642808, 
    0.1190659, -0.06416965, -0.2468681, -0.3436129, -0.4035096, -0.5162868, 
    -0.1552668, -0.03311527, -0.0672785, 0.01909828, 0.1146551, 0.1146877, 
    -0.3191991, -0.7164158, -0.5754166, -0.3704035, -0.1987889, -0.05402979, 
    0.1919989, 0.3954495, 0.2292872, 0.2187078, 0.2433823, 0.007867962, 
    -0.2307876, -0.3619073, -0.3177341, -0.1976985, -0.1168066, -0.07035446, 
    -0.08905554, -0.08055925, -0.05039954, 0.04774404, -0.1270278, -0.3913832,
  -0.4561946, -0.1163344, 0.1366277, 0.02520195, 0.03436536, -0.3158625, 
    -0.7055272, -0.9634212, -1.372454, -0.9583757, -0.4815852, -0.5987726, 
    -0.5889259, -0.4439548, -0.4017187, -0.7132421, -0.9619076, -0.6890234, 
    -0.3217219, -0.1729751, 0.03210354, -0.03355443, -0.1123633, -0.06164703, 
    -0.2178636, -0.2080824, 0.1281803, 0.009023666, -0.08480781, 0.2672434, 
    0.1737211, -0.1210382, 0.1138577, 0.1223693, 0.1347561, 0.164623, 
    -0.08571887, -0.139658, -0.2886165, -0.5363703, -0.7026951, -0.7675227, 
    -0.7148861, -0.6874446, -0.5181576, -0.3147395, -0.2424088, -0.1893, 
    -0.07247061, -0.03886056, -0.07481435, -0.1097101, -0.2050389, 
    -0.2128026, -0.009335804, 0.2579169, 0.3238181, 0.2284894, 0.0597232, 
    0.1122463, 0.1187404, -0.1592707, -0.4343357, -0.4786553, -0.5122321, 
    -0.4506273, -0.2722425, -0.1403091, -0.07216135, -0.02082668, 0.03496754, 
    -0.01477218, -0.4006282, -0.5784926, -0.359173, -0.2591242, -0.07680005, 
    -0.01905298, -0.04468775, -0.01626968, -0.07442391, -0.01843441, 
    -0.0252378, -0.1969987, -0.3097916, -0.4884374, -0.4600521, -0.2011165, 
    -0.1468846, -0.05879873, -0.06584632, -0.1850681, -0.1338634, 0.05718422, 
    0.1677638, -0.1642511,
  0.3948473, 0.3455307, 0.2116114, 0.09784192, 0.05990247, -0.2836685, 
    -0.5812433, -0.9954524, -1.668971, -1.111501, -0.4149836, -0.4221776, 
    -0.6190687, -0.4489191, -0.3332616, -0.562054, -0.7384373, -0.6587498, 
    -0.48624, -0.3313081, -0.01036096, -0.1607517, -0.2869077, -0.09493113, 
    -0.2021253, -0.4490006, -0.2424085, -0.07569313, -0.10569, 0.02098656, 
    0.06532228, -0.09527314, 0.05199313, 0.2439356, 0.3030324, 0.5098209, 
    0.3197498, 0.268497, 0.2745025, 0.1886785, -0.003818244, -0.3023533, 
    -0.470843, -0.5830172, -0.5816662, -0.4650323, -0.3341403, -0.1984141, 
    -0.03983688, 0.1113348, 0.1693915, 0.1176988, -0.08664691, -0.3287696, 
    -0.1970638, 0.2068752, 0.4748765, 0.4140368, 0.1331937, 0.07796872, 
    0.1154037, -0.201328, -0.5749444, -0.5704684, -0.4402275, -0.4247165, 
    -0.5325295, -0.4358658, -0.3073503, 0.002920054, 0.2255926, 0.282575, 
    0.1432033, -0.06167956, -0.283343, -0.3439224, -0.08988594, 0.2337303, 
    0.3073145, 0.1626855, -0.05069327, -0.240586, -0.3932385, -0.476295, 
    -0.4781995, -0.6648526, -0.6673434, -0.3578705, -0.2236258, -0.09577775, 
    0.01257175, -0.01519518, -0.08459604, -0.1506605, 0.07974297, 0.3391017,
  0.2337956, 0.3696681, 0.5355046, 0.549486, 0.2993882, -0.0248957, 
    -0.3978449, -0.8456804, -1.23458, -1.192864, -0.6320573, -0.3375422, 
    -0.2910905, -0.2892188, -0.1205013, -0.1899673, -0.3425716, -0.5029393, 
    -0.5732519, -0.3056086, 0.003571272, 0.009007454, -0.1408622, -0.1239841, 
    -0.1444921, -0.4285254, -0.3268978, -0.07465155, -0.05290693, 0.04972994, 
    0.1139061, 0.05462897, 0.2854564, 0.3969798, 0.3128645, 0.2874744, 
    0.02500659, -0.0959406, 0.01410198, 0.2022698, 0.3627995, 0.318073, 
    0.2111883, 0.1099679, -0.01097941, -0.1253023, -0.09463787, 0.01903367, 
    0.04627967, 0.05251336, 0.1964912, 0.3564196, 0.2421787, -0.06771708, 
    -0.04411697, 0.3864977, 0.757575, 0.7324772, 0.3811104, 0.1599841, 
    0.1452868, -0.1882422, -0.7292415, -0.7017674, -0.248268, -0.3659275, 
    -0.4084406, -0.2957453, -0.4266372, -0.4768325, -0.1404881, 0.1507228, 
    0.2936915, 0.2469304, 0.05807936, 0.1693751, 0.4111882, 0.534691, 
    0.5663314, 0.5667869, 0.3916732, 0.1127839, -0.2371352, -0.6997647, 
    -0.970598, -0.935637, -0.6524177, -0.2609465, -0.1813564, -0.2540128, 
    -0.1962492, -0.07230794, 0.03475595, -0.04533839, -0.1008723, 0.06623393,
  0.1436589, 0.4032293, 0.6637273, 0.5954981, 0.303213, 0.2335027, 0.2061752, 
    0.1325425, -0.2114354, -0.743955, -0.8611587, -0.4466405, -0.09909809, 
    0.1212795, 0.1014389, 0.00298515, -0.1425389, -0.277744, -0.1646417, 
    0.1735585, 0.0693264, -0.0923599, -0.0388117, 0.01870782, -0.01374661, 
    -0.06031238, -0.02492839, 0.08003598, 0.02004245, -0.001344264, 
    0.1343652, 0.2429592, 0.3111559, 0.2134507, 0.03872752, 0.1451402, 
    -0.004241228, -0.1631118, -0.2481705, -0.0308032, 0.1648669, 0.2026759, 
    0.1817937, 0.09489599, 0.01509452, -0.03983712, -0.07513952, 0.006777763, 
    0.1436594, 0.125788, 0.1134834, 0.2605863, 0.3637276, 0.282917, 0.288825, 
    0.6471102, 1.146671, 1.315795, 0.9686925, 0.3890862, 0.0473702, 
    -0.2623625, -0.7064219, -0.6367122, -0.2966568, -0.5952734, -0.6412369, 
    -0.3849706, -0.513893, -0.7676366, -0.4008071, 0.05977228, 0.3705145, 
    0.4066795, 0.245726, 0.2549708, 0.5284082, 0.8608139, 1.182705, 1.273021, 
    0.924079, 0.4236557, 0.03140295, -0.4276139, -1.010231, -1.478199, 
    -1.448316, -0.8248138, -0.3090425, -0.1830008, -0.1394787, -0.0180428, 
    0.1688061, 0.1710029, 0.01543617, 0.03184259,
  0.6276759, 0.9392484, 0.9212795, 0.7033269, 0.4588771, 0.3233139, 
    0.2753485, 0.460635, 0.5986068, 0.3431705, 0.05527997, -0.09096026, 
    -0.08905584, 0.04365897, 0.2866115, 0.2532457, 0.2170477, 0.07027031, 
    -0.1041274, 0.1122954, -0.1559179, -0.212119, 0.005280077, 0.007835422, 
    -0.1230727, -0.149147, -0.04239243, 0.1111883, 0.09828139, 0.03791356, 
    0.1058172, 0.1843164, 0.2069894, 0.1803615, 0.1318427, 0.189379, 
    0.06963396, -0.1823661, -0.3023207, -0.3733822, -0.4413505, -0.5018651, 
    -0.3216733, -0.2214452, -0.3155695, -0.3223404, -0.188128, -0.08163381, 
    -0.03723264, -0.008684635, -0.04476857, -0.1056893, 0.01372814, 
    0.3094628, 0.5933499, 0.8431547, 1.182852, 1.461499, 1.417472, 0.975121, 
    0.335098, -0.3003187, -0.7829692, -0.5908942, 0.0654366, -0.1735446, 
    -0.5936619, -0.5825943, -0.6258886, -0.7493747, -0.5652115, -0.2808039, 
    0.08792982, 0.4331609, 0.5179918, 0.1877996, 0.133047, 0.2883366, 
    0.9561425, 1.322207, 1.341348, 0.9962958, 0.4943427, 0.07671535, 
    -0.3892026, -1.017669, -1.443157, -1.384774, -1.029111, -0.6285257, 
    -0.2401953, 0.0252347, 0.2233791, 0.4261794, 0.460603, 0.5380762,
  0.7445543, 0.8117251, 0.6704657, 0.5442775, 0.5167872, 0.4798731, 
    0.2818751, 0.3156479, 0.6626205, 0.779987, 0.6783433, 0.416006, 
    0.2009666, 0.2185613, 0.3050684, 0.2336001, 0.3730048, 0.3128647, 
    -0.01410455, -0.1187761, -0.06999648, -0.08065736, -0.06088221, 
    0.02749687, 0.03765312, 0.04821628, 0.04315443, 0.07013988, 0.04914379, 
    0.06039071, 0.1664941, 0.1517483, 0.1525133, 0.1862534, 0.0975652, 
    0.04017591, 0.1103585, 0.1801, 0.04668474, 0.2234764, 0.5109932, 
    0.4319243, 0.2548895, 0.2903386, 0.1381414, -0.2077082, -0.2595962, 
    -0.0009862185, 0.1666734, 0.1180569, 0.09759796, -0.0543716, -0.1769135, 
    0.06668973, 0.5590401, 0.9246483, 1.162084, 1.454484, 1.671345, 1.488028, 
    0.8172925, -0.008879662, -0.5190203, -0.4439216, 0.08473992, -0.1108165, 
    -0.1992607, -0.3242934, -0.5727147, -0.7087173, -0.53541, -0.3492284, 
    -0.2330011, -0.2219012, 0.09740245, 0.2662989, 0.3445379, 0.2763087, 
    0.2524318, 0.5633204, 1.339167, 1.519977, 1.214704, 0.7935289, 0.3400942, 
    -0.2879653, -0.9241469, -1.450725, -1.621477, -1.248773, -0.5906024, 
    -0.2579846, -0.03505182, 0.3505273, 0.6292057, 0.6167879,
  0.7171774, 0.7694235, 0.7549059, 0.405931, 0.2247462, 0.1502508, 0.1034409, 
    0.1387599, 0.3144436, 0.4237698, 0.5742903, 0.6422428, 0.6150455, 
    0.6075423, 0.4833238, 0.4056382, 0.5333074, 0.5535223, 0.2798407, 
    0.09785831, 0.1977766, 0.1932034, -0.008619308, -0.04797482, 0.03902054, 
    0.02194691, -0.001767635, -0.02743477, -0.04087865, -0.01571596, 
    0.008502841, 0.06104183, 0.1114163, 0.09553099, -0.1042414, -0.1497983, 
    0.03685561, -0.1146253, -0.5515227, -1.053575, 0.7686257, 1.300414, 
    0.739542, 0.3349841, 0.2002183, -0.2174252, -0.62999, -0.3576268, 
    -0.02723947, 0.01590833, 0.1200263, 0.3375556, 0.4151596, 0.4426012, 
    0.8282944, 1.384056, 1.614004, 1.605068, 1.646865, 1.592145, 1.198966, 
    0.5693591, 0.03666067, -0.218011, -0.2593356, -0.2664323, -0.2437271, 
    -0.3257909, -0.510182, -0.5472263, -0.4430923, -0.2856542, -0.2417739, 
    -0.2426366, -0.09774727, 0.2184637, 0.35681, 0.3616276, 0.3178776, 
    0.5224839, 0.9569572, 1.069685, 1.408698, 1.449339, 1.062051, 0.3960679, 
    -0.1596452, -0.6751074, -1.142458, -1.187102, -0.8111091, -0.4187589, 
    -0.1487722, 0.09494495, 0.28352, 0.4426508,
  0.3910551, 0.1802316, 0.1647856, 0.3473215, 0.4399478, 0.1613998, 
    -0.1340427, -0.1296647, -0.004160047, 0.1992089, 0.2712467, 0.2667872, 
    0.2162989, 0.2090074, 0.2495184, 0.2906318, 0.4324775, 0.5618882, 
    0.542552, 0.4139552, 0.3480536, 0.3565173, 0.2500401, 0.1419663, 
    0.02844119, -0.07819974, -0.06644833, -0.04986322, -0.04390615, 
    -0.06078437, -0.02126616, 0.05697298, 0.1132879, 0.0498116, -0.2792087, 
    -0.3389418, -0.01897073, -0.3793063, -0.8372159, -1.793044, -0.3492765, 
    0.6467032, 0.3911688, 0.08519626, 8.821487e-005, -0.3412859, -0.8115654, 
    -0.821478, -0.5079198, -0.3406184, -0.1822362, 0.1909408, 0.4399642, 
    0.5821193, 1.02141, 1.659251, 1.919375, 1.623167, 1.401813, 1.446621, 
    1.369522, 0.9124579, 0.2561754, 0.02170241, -0.01687157, -0.02592134, 
    -0.03842109, -0.1140721, -0.127093, -0.08996731, -0.1057225, -0.1153579, 
    -0.1045183, -0.1081153, -0.2157977, -0.1141047, -0.07854153, 0.1845444, 
    0.3939844, 0.5527086, 0.7189034, 0.647094, 1.085603, 1.29226, 0.7933499, 
    0.1040757, -0.236403, -0.4098241, -0.7422458, -1.028395, -1.015992, 
    -0.6640062, -0.1975517, 0.2543037, 0.5484931, 0.5751536,
  0.3558502, 0.2225819, 0.2703357, 0.5104883, 0.5159085, 0.2167547, 
    -0.1284275, -0.2592869, -0.2499282, -0.1551691, -0.05321604, 
    0.0005599856, 0.008795679, -0.01273763, -0.0749284, -0.1233822, 
    -0.1636163, -0.09385741, -0.09462214, -0.05020475, 0.0388577, 0.1078193, 
    0.1251214, 0.06480217, -0.005168915, -0.08423805, -0.1507257, -0.1756771, 
    -0.194183, -0.2073829, -0.2232355, -0.1850032, -0.08116198, -0.05381835, 
    -0.192474, -0.2826428, -0.245029, -0.3871677, -0.4226174, -0.9903107, 
    -0.7179952, -0.4084888, -0.1142347, -0.1957772, -0.7327423, -0.340961, 
    -0.4881783, -0.4032643, -0.04818606, 0.2280672, 0.3599684, 0.3371007, 
    0.2999744, 0.3439521, 0.540892, 1.157054, 1.474632, 1.4586, 1.350609, 
    1.342894, 1.100902, 0.8663803, 0.4812242, 0.2514713, 0.2508204, 
    0.2960516, 0.2341212, 0.09149423, 0.0523504, 0.1008855, 0.06423187, 
    -0.04271781, -0.1718524, -0.4011328, -0.6428974, -0.626572, -0.4269302, 
    0.01800795, 0.2804427, 0.2451565, 0.2491608, 0.08976984, 0.7558172, 
    1.117765, 0.6775627, 0.08091497, -0.338161, -0.4881281, -0.5830337, 
    -0.7087498, -0.825205, -0.8924083, -0.7613697, -0.3970468, 0.07453489, 
    0.391283,
  -0.3702729, -0.01747417, 0.355118, 0.3097725, 0.3072657, 0.4624578, 
    0.192894, 0.03690445, -0.1818293, -0.2796322, -0.2816828, -0.2246191, 
    -0.1908464, -0.1570248, -0.08796537, -0.0560807, -0.04916328, 
    -0.07107091, -0.1053319, -0.1135515, -0.1586523, -0.1467869, -0.1441503, 
    -0.132285, -0.1318781, -0.1699314, -0.1661881, -0.1779558, -0.1968035, 
    -0.207041, -0.2334733, -0.2034439, -0.1278579, -0.1105891, -0.1162369, 
    -0.1656184, -0.1888282, -0.2654717, -0.3428643, -0.3700447, -0.2649674, 
    -0.2145448, -0.2951097, -0.4142022, -0.5529711, -0.6672959, -0.8907495, 
    -1.816759, -1.650271, -1.451427, -1.168337, -0.7883394, -0.1568773, 
    0.06089509, 0.2770737, 0.4131087, 0.5261297, 0.6010484, 0.5802963, 
    0.6545963, 0.7078841, 0.6056542, 0.4522036, 0.3111884, 0.247907, 
    0.2477117, 0.195368, 0.07562512, 0.01945651, 0.05532891, 0.06641275, 
    0.09294271, -0.05129528, -0.1520603, -0.1769302, -0.1775814, -0.1081965, 
    0.04390311, 0.2196354, 0.2157788, 0.1609774, 0.1489167, 0.430053, 
    0.4515042, 0.3386137, 0.01008177, -0.3404059, -0.8152928, -1.1289, 
    -1.184238, -1.034157, -0.8767511, -0.9036554, -0.9967377, -0.9668874, 
    -0.7346931,
  -0.6113862, -0.5634041, -0.4509535, -0.0267179, 0.06123734, 0.1080146, 
    0.197565, -0.05941731, -0.1927505, -0.2612728, -0.2500586, -0.179925, 
    -0.1639744, -0.1606541, -0.1335059, -0.1138933, -0.08189428, -0.07909495, 
    -0.04149729, 0.03864592, 0.08381176, 0.05399442, -0.04113901, -0.1285253, 
    -0.1168227, -0.1309177, -0.1025, -0.1098729, -0.163535, -0.210996, 
    -0.2722427, -0.3518, -0.3843033, -0.413177, -0.3692316, -0.3179458, 
    -0.3238704, -0.2261978, -0.1867772, -0.1566339, -0.08428669, -0.2129819, 
    -0.2561779, -0.4255466, -0.6219984, -0.8857517, -0.9601169, -0.9698019, 
    -0.8803, -0.7295027, -0.6562934, -0.6379652, -0.305738, 0.00425446, 
    0.1801009, 0.2410385, 0.2331935, 0.2134181, 0.2052963, 0.2363508, 
    0.2632389, 0.2689683, 0.3065659, 0.3544662, 0.3066635, 0.2112534, 
    0.09561212, 0.03062188, 0.08698581, 0.1858464, 0.2387762, 0.2506738, 
    0.1535386, 0.01821959, 0.003278255, 0.009007156, 0.05785155, 0.1255436, 
    0.2887763, 0.4507561, 0.5853264, 0.5619378, 0.2494043, 0.01791029, 
    -0.1275163, -0.1743584, -0.1344657, -0.4238396, -0.5180449, -0.650825, 
    -0.783587, -0.4187436, -0.2783952, -0.2193616, -0.3840754, -0.5501724,
  0.01836602, -0.2483985, -0.4328545, -0.4199963, -0.2594171, 0.06402063, 
    0.128669, 0.0548408, -0.09245741, -0.2015723, -0.2071873, 0.1086818, 
    0.2377345, 0.1960678, 0.0854882, 0.08413744, 0.02170241, -0.006210685, 
    0.08542329, 0.2198959, 0.3093652, 0.2749416, 0.1169503, -0.0410409, 
    -0.07338119, 0.02347708, 0.06476915, 0.05850267, -0.06934556, -0.2221613, 
    -0.369606, -0.5613216, -0.7294366, -0.7491797, -0.5389743, -0.4183204, 
    -0.3121841, -0.2557388, -0.2671483, -0.313421, -0.3638607, -0.3368263, 
    -0.3350683, -0.3353448, -0.4905207, -0.6186944, -0.7031508, -0.5624605, 
    -0.4609468, -0.1618419, -0.1051044, -0.2082288, -0.2750745, -0.1687598, 
    -0.109759, -0.009645045, 0.01743829, 0.04569346, 0.1185288, 0.1322983, 
    0.1640366, 0.2335353, 0.3178777, 0.3755274, 0.3699124, 0.3218816, 
    0.2229233, 0.1815171, 0.1950099, 0.3151271, 0.3370346, 0.4039454, 
    0.3224187, 0.2567122, 0.2310615, 0.3486723, 0.2640364, 0.2933171, 
    0.3184636, 0.3532617, 0.3818752, 0.4160874, 0.1669501, -0.2295015, 
    -0.5913019, -0.6970474, -0.6256766, -0.4185004, -0.1756787, -0.1607699, 
    -0.2869902, -0.3232841, -0.6278906, -0.4928637, 0.2239487, 0.2647691,
  0.6572988, 0.6771063, 0.642487, 0.7099024, 0.8258694, 0.909691, 0.8765693, 
    0.638304, 0.4009994, 0.1312403, 0.04408216, 0.05148774, 0.09240574, 
    0.1662339, 0.06382501, 0.02232099, 0.1170151, 0.1367579, 0.2214747, 
    0.3397363, 0.3918197, 0.362637, 0.2506092, 0.1105378, 0.03034592, 
    0.04312205, 0.1310939, 0.2022362, 0.1685125, 0.003945448, -0.1518163, 
    -0.3123145, -0.4663669, -0.5253353, -0.4832292, -0.4956802, -0.2665949, 
    -0.2268977, -0.3354262, -0.3534927, -0.2962173, -0.3047134, -0.3587986, 
    -0.4131118, -0.501035, -0.5915459, -0.6329035, -0.6220477, -0.5782647, 
    -0.5298761, -0.4885674, -0.4321547, -0.3505795, -0.2921486, -0.2465753, 
    -0.1521417, -0.09058589, -0.07123363, -0.04693353, -0.02175444, 
    0.003294408, 0.05656589, 0.10834, 0.1970606, 0.2279201, 0.2556382, 
    0.2289941, 0.2002182, 0.1948471, 0.3431543, 0.2763086, 0.3271388, 
    0.4452214, 0.3733628, 0.355866, 0.3574772, 0.4215398, 0.6262441, 
    0.4623929, 0.3383042, 0.3723374, 0.2422103, -0.09564686, -0.6491957, 
    -0.9950452, -0.994638, -0.9787533, -0.879225, -0.7614996, -0.6027932, 
    -0.3647242, -0.1548438, 0.06317425, 0.199306, 0.254467, 0.08194089,
  0.6107821, 0.8236728, 1.032722, 1.043203, 0.910163, 0.792357, 0.6767155, 
    0.5067611, 0.4162502, 0.3257878, 0.178164, 0.114834, 0.07140946, 
    0.04557949, 0.03628594, 0.03125665, 0.06861016, 0.1116928, 0.1396876, 
    0.2285874, 0.2952703, 0.3206446, 0.3205957, 0.2843001, 0.1827542, 
    0.2890855, 0.2475165, 0.2186425, 0.1906154, 0.1271877, 0.003994286, 
    -0.1411229, -0.309222, -0.3962825, -0.4816992, -0.5073177, -0.534287, 
    -0.5758886, -0.6214126, -0.6563247, -0.6914321, -0.6911228, -0.6768162, 
    -0.6621678, -0.6446384, -0.6270441, -0.5993259, -0.5632095, -0.5193456, 
    -0.4656024, -0.4060807, -0.3414811, -0.2758234, -0.1976984, -0.1501399, 
    -0.1138606, -0.08554018, -0.07769519, -0.08142245, -0.07894844, 
    -0.07940418, -0.08936512, -0.08843726, -0.09104154, -0.03301746, 
    -0.0225845, 0.002138853, 0.0338282, 0.1203191, 0.2428776, 0.332461, 
    0.3676823, 0.4042383, 0.3362044, 0.3768621, 0.4358139, 0.2954329, 
    0.3273503, 0.2798569, 0.1897527, 0.176748, -0.04257131, -0.3187425, 
    -0.5363209, -0.5862556, -0.5692151, -0.5006281, -0.4036881, -0.2578218, 
    -0.06122303, 0.04225969, 0.298851, 0.4416237, 0.5466857, 0.5701234, 
    0.6890042,
  0.7299874, 0.7860583, 0.8326889, 0.7944241, 0.6988184, 0.6016178, 
    0.5218652, 0.3804265, 0.3141341, 0.2688216, 0.2221582, 0.2086979, 
    0.2017969, 0.187295, 0.1824285, 0.1809311, 0.1776108, 0.1892807, 
    0.199616, 0.2217514, 0.258226, 0.309642, 0.3370509, 0.3356349, 0.3137924, 
    0.2926012, 0.2413151, 0.1371321, 0.02232099, -0.04914701, -0.140244, 
    -0.1705663, -0.1949152, -0.2200944, -0.2504655, -0.2956151, -0.3691666, 
    -0.4572525, -0.5349055, -0.598675, -0.6643651, -0.7159765, -0.751328, 
    -0.7574641, -0.7628677, -0.7644628, -0.7530369, -0.7340102, -0.7057876, 
    -0.6677343, -0.6096125, -0.5433039, -0.4633397, -0.3820897, -0.307578, 
    -0.2553319, -0.2112564, -0.1750747, -0.1371028, -0.1250096, -0.1284275, 
    -0.1186783, -0.1108332, -0.1145116, -0.1134374, -0.1078224, -0.09013033, 
    -0.03573585, 0.05344057, 0.1411197, 0.2076725, 0.3518783, 0.4117254, 
    0.4198959, 0.3873602, 0.4075263, 0.3898013, 0.3801988, 0.4051175, 
    0.355443, 0.2780015, 0.209235, 0.1534894, 0.08726287, 0.0622139, 
    0.04751611, 0.04727227, 0.04286122, 0.05098331, 0.06869173, 0.09297562, 
    0.1962636, 0.337328, 0.504353, 0.5826571, 0.6607168,
  0.5571355, 0.6095607, 0.6319078, 0.6459378, 0.6461003, 0.6138738, 
    0.5720443, 0.522207, 0.4634668, 0.409056, 0.3598535, 0.3209864, 
    0.2841863, 0.249144, 0.2290268, 0.2249741, 0.2299057, 0.24584, 0.2709376, 
    0.3047267, 0.3362696, 0.3571355, 0.3480861, 0.3123438, 0.2549708, 
    0.188711, 0.1093653, 0.04548192, -0.01696944, -0.08283842, -0.1542578, 
    -0.2113705, -0.2762631, -0.3275163, -0.3701433, -0.4099707, -0.4420019, 
    -0.4655045, -0.4842057, -0.4912533, -0.4987077, -0.5021908, -0.4955176, 
    -0.4948176, -0.4869562, -0.473854, -0.4539322, -0.4414159, -0.416302, 
    -0.3895767, -0.3652115, -0.3342219, -0.2973566, -0.247438, -0.2128189, 
    -0.1739191, -0.1405207, -0.111468, -0.09099266, -0.07640928, -0.05749655, 
    -0.03947896, -0.01989901, 0.003180385, 0.005084515, 0.008144379, 
    0.01852846, 0.01675451, 0.02144194, 0.02503914, 0.01756859, 0.002562046, 
    -0.002239451, 0.0003484488, 0.02254879, 0.02910817, 0.030931, 0.04782557, 
    0.09208012, 0.1105211, 0.1032292, 0.1249576, 0.1075912, 0.1027086, 
    0.08517918, 0.06061862, 0.04103854, 0.02399755, -0.0007745028, 
    0.05697262, 0.114069, 0.1816145, 0.2448144, 0.3281478, 0.4101952, 
    0.4898666,
  0.2102604, 0.2297917, 0.2400293, 0.2562728, 0.2756087, 0.2861556, 
    0.2948308, 0.3066146, 0.3105861, 0.30917, 0.3095281, 0.3099025, 
    0.3069728, 0.2951075, 0.2905828, 0.291006, 0.2917221, 0.2822332, 
    0.2747788, 0.2638087, 0.2533921, 0.2363186, 0.2150295, 0.1933661, 
    0.1656969, 0.1412177, 0.1094794, 0.07253277, 0.04287767, 0.004840732, 
    -0.03807932, -0.07914376, -0.1188736, -0.1536067, -0.1907974, -0.2259048, 
    -0.2632746, -0.295013, -0.3216569, -0.3422949, -0.3555924, -0.3652604, 
    -0.3711849, -0.3752213, -0.3708919, -0.3694595, -0.365895, -0.3605891, 
    -0.3507583, -0.3434178, -0.3339126, -0.3227798, -0.3146255, -0.3054458, 
    -0.2908788, -0.2724542, -0.2537205, -0.233587, -0.2149509, -0.1941176, 
    -0.1729913, -0.1518813, -0.1278904, -0.1180271, -0.106227, -0.08903956, 
    -0.08583319, -0.08907205, -0.08918595, -0.08975559, -0.09537089, 
    -0.0984633, -0.1009698, -0.0964939, -0.09514299, -0.09195295, 
    -0.09367818, -0.0933364, -0.08903953, -0.08430323, -0.07561186, 
    -0.06677395, -0.0571548, -0.04501286, -0.03042954, -0.01630196, 
    -0.0003840327, 0.01805669, 0.03753912, 0.0588932, 0.08589512, 0.1057845, 
    0.1289127, 0.153457, 0.1725326, 0.1920964,
  0.1296897, 0.1430202, 0.1579943, 0.1736846, 0.1891961, 0.2065949, 0.223815, 
    0.2397165, 0.254365, 0.2669296, 0.2763209, 0.2827983, 0.2878928, 
    0.2920272, 0.2938504, 0.292418, 0.2881544, 0.2808304, 0.2695835, 
    0.2550327, 0.2381543, 0.2184927, 0.1953808, 0.1689159, 0.1389029, 
    0.1055046, 0.0711621, 0.03558266, -1.311302e-005, -0.03362346, 
    -0.06606174, -0.09628677, -0.1238258, -0.148777, -0.1695933, -0.186748, 
    -0.199769, -0.2095838, -0.213913, -0.2124305, -0.2060995, -0.1934538, 
    -0.1758265, -0.1525517, -0.1252732, -0.09628439, -0.06947899, 
    -0.03993797, -0.01052713, 0.02264309, 0.04840803, 0.06945324, 0.0682168, 
    0.09666586, 0.0240097, 0.1037621, 0.08663988, 0.09090424, 0.06766224, 
    -0.003936052, 0.05753851, 0.02768826, 0.03281522, 0.01497674, 
    0.009817362, 0.006529331, 0.002151012, -0.002699137, -0.01156974, 
    0.00530839, 0.01041889, 0.01004505, 0.001776695, -0.02061939, 0.03125238, 
    0.03271866, 0.02868128, 0.02825785, 0.05687189, 0.07552338, 0.09368753, 
    0.1112492, 0.127444, 0.1389837, 0.1461132, 0.1489453, 0.1476433, 
    0.1436718, 0.1380403, 0.1315135, 0.1249053, 0.1179886, 0.1119494, 
    0.1107287, 0.1134629, 0.1198266,
  0.3112659, 0.380146, 0.4452014, 0.5041203, 0.5451202, 0.5649438, 0.5661967, 
    0.5571148, 0.5431175, 0.5276389, 0.5079291, 0.4824085, 0.4536817, 
    0.4215529, 0.3846554, 0.348799, 0.3165072, 0.2899772, 0.2662956, 
    0.2433463, 0.2176464, 0.1895702, 0.1565136, 0.1219758, 0.08922845, 
    0.06063163, 0.03875649, 0.0224154, 0.01051712, 0.0007998943, -0.01417398, 
    -0.03884792, -0.07603884, -0.1273069, -0.1894169, -0.2551723, -0.3190722, 
    -0.3698206, -0.4015265, -0.4115524, -0.4252729, -0.3306603, -0.2133918, 
    -0.1596479, -0.08464813, -0.02388954, 0.06048536, 0.1260285, 0.1831894, 
    0.1829774, 0.2257512, 0.2281115, 0.2381051, 0.2603869, 0.2052931, 
    0.3015495, 0.3194693, 0.3221548, 0.3355664, 0.3344434, 0.337357, 
    0.3103223, 0.2635937, 0.1983757, 0.1431675, 0.07666373, 0.02568686, 
    -0.03396493, -0.0869597, -0.151836, -0.2360806, -0.2961559, -0.3370254, 
    -0.384975, -0.3905082, -0.4036098, -0.4084435, -0.3856735, -0.389873, 
    -0.3667121, -0.259275, -0.2212379, -0.02099371, -0.01306605, 0.1013542, 
    0.179121, 0.2525911, 0.2869011, 0.2963407, 0.283108, 0.2601104, 0.236918, 
    0.2190623, 0.2125521, 0.2220087, 0.2530465,
  0.372366, 0.4372091, 0.4772809, 0.4760931, 0.4395378, 0.3886591, 0.3462598, 
    0.32069, 0.2957714, 0.2521354, 0.1740918, 0.07736325, -0.007158756, 
    -0.06173205, -0.07763457, -0.05844498, -0.01884508, 0.01650667, 
    0.03403652, 0.03631508, 0.0393912, 0.05547193, 0.08068347, 0.08714509, 
    0.05081698, -0.003903091, -0.04169583, -0.05058265, -0.03964496, 
    -0.03588581, -0.04763722, -0.07063508, -0.09161568, -0.1037412, 
    -0.1119442, -0.1302061, -0.1550589, -0.1926236, -0.2283645, -0.2421994, 
    -0.2286735, -0.1704888, 0.02005482, 0.05789614, 0.07057548, 0.1360703, 
    0.1761096, 0.219306, 0.2554228, 0.2623894, 0.2362498, 0.1839062, 
    0.1586459, 0.1593456, 0.1543814, 0.1432487, 0.1264682, 0.1297879, 
    0.106708, 0.05247641, -0.04893875, -0.1832976, -0.3383112, -0.4650688, 
    -0.5702934, -0.6339811, -0.6870573, -0.7288217, -0.7598925, -0.7628391, 
    -0.7228329, -0.6283669, -0.5005016, -0.3964634, -0.3886194, -0.4255986, 
    -0.4452767, -0.6074839, -0.5535936, -0.4670553, -0.316843, -0.155026, 
    -0.001428962, 0.1037142, 0.2038281, 0.2801952, 0.3592644, 0.4466504, 
    0.5018101, 0.5380888, 0.5375834, 0.4789734, 0.4194365, 0.3680534, 
    0.3323765, 0.3379583,
  0.4409375, 0.5050161, 0.5692089, 0.5875194, 0.5396516, 0.4271027, 0.300459, 
    0.1956086, 0.1224475, 0.06639242, 0.02334261, 0.01417875, 0.06312084, 
    0.1558299, 0.2468138, 0.2872257, 0.2949407, 0.2497098, 0.1726267, 
    0.04236972, -0.08878255, -0.1228979, -0.05614948, 0.04459906, 0.1052115, 
    0.08929372, 0.06504224, 0.07095063, 0.08572924, 0.08688486, 0.07345712, 
    0.04378593, 0.007571578, -0.02629888, -0.06082022, -0.08183265, 
    -0.09434891, -0.1091444, -0.1138806, -0.08997178, -0.05479908, 
    -0.04690456, 0.03846359, 0.1097202, 0.08633089, 0.04253197, 0.2370305, 
    0.2454941, 0.2226753, 0.1606805, 0.1358432, 0.1351919, 0.1008983, 
    0.09188144, 0.1400096, 0.1952507, 0.2215527, 0.2118034, 0.1594923, 
    0.01011062, -0.1260383, -0.1915658, -0.2580861, -0.3566374, -0.4804003, 
    -0.6150521, -0.671628, -0.714874, -0.7079887, -0.6433563, -0.542624, 
    -0.4393687, -0.3571258, -0.3314428, -0.3225241, -0.3622692, -0.3812473, 
    -0.3464165, -0.2506802, -0.1306772, -0.08541322, 0.08159518, 0.193444, 
    0.2758008, 0.3457714, 0.3911491, 0.4188346, 0.4166698, 0.4156609, 
    0.3684279, 0.4125358, 0.4700718, 0.474189, 0.4977076, 0.4766145, 0.4466506,
  0.08468699, 0.1542509, 0.2804387, 0.3373885, 0.3059597, 0.2529168, 
    0.1502805, 0.0588913, -0.1124153, -0.09130478, -0.06195927, -0.06375074, 
    -0.06370163, -0.05421257, -0.03274465, 0.009883404, -0.02535439, 
    -0.1760702, -0.2769175, -0.2549771, -0.2940561, -0.350518, -0.1879044, 
    0.05908489, 0.3375357, 0.5649284, 0.647903, 0.5716176, 0.4187045, 
    0.241864, 0.1303248, 0.07078743, 0.0381701, 0.004901886, -0.0629859, 
    -0.1417456, -0.2414041, -0.337904, -0.3807263, -0.3213329, -0.2416306, 
    -0.1867805, -0.2280073, -0.3032346, -0.4042773, -0.4689097, -0.2095513, 
    -0.08547974, 0.008482695, 0.02021813, 0.02042973, 0.00288409, 0.03950512, 
    0.1655631, 0.2761913, 0.2818879, 0.2373567, 0.1730826, 0.02894197, 
    -0.1025033, -0.1778452, -0.1646127, -0.1613411, -0.1849414, -0.1961719, 
    -0.3150848, -0.4474741, -0.5082811, -0.529261, -0.5401982, -0.6287237, 
    -0.5300748, -0.6233039, -0.8029101, -0.7983853, -0.7040819, -0.6526335, 
    -0.4752897, -0.3613411, -0.203382, -0.01215482, 0.1484407, 0.3019402, 
    0.3998404, 0.4637402, 0.5282422, 0.5590038, 0.5365916, 0.5156933, 
    0.47694, 0.4452668, 0.2295929, 0.1896842, 0.1311718, 0.08319008, 
    0.06810224,
  -0.05040368, -0.007662773, -0.008053541, 0.04162109, 0.08322215, 0.0998559, 
    0.1286483, 0.2358255, 0.284915, 0.3068871, 0.2282743, 0.07264328, 
    -0.1656056, -0.4149706, -0.5345516, -0.4137502, -0.2070274, -0.07672119, 
    0.003730774, -0.05175447, -0.08171916, -0.1394175, -0.09364915, 
    0.02568686, 0.2451034, 0.3991241, 0.4072299, 0.2648144, 0.01691437, 
    -0.2112112, -0.3592749, -0.3924947, -0.4007626, -0.436553, -0.5039511, 
    -0.5561328, -0.5294719, -0.4483042, -0.4139457, -0.2950001, -0.2712045, 
    -0.2734494, -0.3423309, -0.4654918, -0.4458466, -0.4955211, -0.3446755, 
    -0.2995093, 0.04598284, 0.2930046, 0.3250684, 0.2333853, 0.1336946, 
    0.1248893, 0.1530793, 0.1473828, 0.1001496, 0.007132053, -0.1316701, 
    -0.2296191, -0.2290007, -0.1270476, -0.02253914, -0.0956023, -0.3629525, 
    -0.661325, -0.8775846, -1.033688, -1.080059, -1.080775, -1.083688, 
    -0.9418424, -1.025664, -1.171042, -1.242314, -1.09946, -0.8555632, 
    -0.6057584, -0.350957, -0.1154426, 0.1796745, 0.3400098, 0.4017774, 
    0.4275097, 0.4222201, 0.4092481, 0.3512403, 0.2450065, 0.1756055, 
    0.1341503, 0.07249659, 0.0427441, 0.0735873, 0.07291996, 0.05859697, 
    -0.02515954,
  -0.7177215, -0.7395964, -0.6720183, -0.5827603, -0.4676887, -0.3582158, 
    -0.2295053, -0.1120899, -0.01537776, 0.01891613, 0.05296552, 0.02205721, 
    -0.1068979, -0.241517, -0.4353808, -0.5743456, -0.4945288, -0.3563616, 
    -0.1728816, -0.03691196, -0.09994888, -0.06791711, -0.1256638, 
    -0.1603808, -0.1341602, -0.1225228, 0.001435757, -0.08277702, -0.177048, 
    -0.1854948, -0.179603, -0.2374967, -0.2922819, -0.337301, -0.5879369, 
    -0.6746233, -0.4312799, -0.7838027, -0.6620893, -0.5544887, -0.4767547, 
    -0.5846164, -0.7423472, -0.9015272, -0.9682913, -0.9085575, -0.6769336, 
    -0.4592742, -0.2798634, -0.2367319, -0.2818815, -0.2784474, -0.1977345, 
    -0.1668749, -0.2245898, -0.2955533, -0.3521126, -0.3816373, -0.4063933, 
    -0.4310027, -0.4133269, -0.3466765, -0.3264617, -0.4328582, -0.6983367, 
    -0.9990691, -1.170342, -1.226071, -1.287644, -1.321937, -1.385739, 
    -1.461244, -1.488718, -1.439076, -1.366957, -1.226494, -1.020374, 
    -0.7267221, -0.3894174, -0.05424488, 0.2229688, 0.2599642, 0.2340363, 
    0.1055696, -0.04688808, -0.1523894, -0.3130991, -0.473532, -0.6181935, 
    -0.7113413, -0.7401336, -0.6899057, -0.5731414, -0.4759083, -0.5308074, 
    -0.6564096,
  -1.42542, -1.526429, -1.577503, -1.516094, -1.308232, -1.066842, 
    -0.8624154, -0.8554004, -0.9477017, -0.951901, -0.837985, -0.6893197, 
    -0.6087533, -0.6785449, -0.8918751, -1.174329, -1.381816, -1.48696, 
    -1.52822, -1.544854, -1.477097, -1.301462, -1.025176, -0.8550912, 
    -0.8067189, -0.7913055, -0.7812794, -0.7932748, -0.8380177, -0.902959, 
    -0.9197884, -0.9145637, -1.001982, -1.206784, -1.480124, -1.7186, 
    -1.767982, -1.619853, -1.416175, -1.261211, -1.253512, -1.359095, 
    -1.509323, -1.610625, -1.596449, -1.44679, -1.25877, -1.124167, 
    -1.070879, -1.032061, -0.9444467, -0.7859831, -0.6585745, -0.6592907, 
    -0.7620901, -0.8786263, -0.905791, -0.8852181, -0.9128223, -1.080954, 
    -1.165052, -1.037806, -0.9298958, -0.9324511, -1.025599, -1.188083, 
    -1.299492, -1.373971, -1.391777, -1.408102, -1.393226, -1.395635, 
    -1.430107, -1.520993, -1.583037, -1.438685, -1.15929, -0.8285612, 
    -0.5850392, -0.4844368, -0.5540821, -0.6529753, -0.6334766, -0.4936002, 
    -0.3995573, -0.4673633, -0.7062631, -0.9918913, -1.139417, -1.212269, 
    -1.248402, -1.252617, -1.222311, -1.159909, -1.152747, -1.26043,
  -1.164417, -1.164515, -1.152878, -1.150957, -1.036374, -0.8085419, 
    -0.5997363, -0.5629036, -0.6056123, -0.6426241, -0.691957, -0.7718723, 
    -0.8880668, -1.036716, -1.206524, -1.334942, -1.400795, -1.466176, 
    -1.600828, -1.700193, -1.628903, -1.394691, -1.15418, -1.03665, 
    -1.058493, -1.1575, -1.260739, -1.372425, -1.495326, -1.541778, 
    -1.485154, -1.402292, -1.422149, -1.54334, -1.629311, -1.700665, 
    -1.760951, -1.75532, -1.636423, -1.47713, -1.391908, -1.433412, 
    -1.494464, -1.577634, -1.63128, -1.534779, -1.386488, -1.324103, 
    -1.336163, -1.308998, -1.217201, -1.161277, -1.18543, -1.262334, 
    -1.307809, -1.269056, -1.220163, -1.247197, -1.425029, -1.556296, 
    -1.481881, -1.258102, -1.05986, -1.081931, -1.189824, -1.220033, 
    -1.232679, -1.23416, -1.209128, -1.179408, -1.305449, -1.555336, 
    -1.803968, -1.905678, -1.845277, -1.5985, -1.249574, -0.9569474, 
    -0.8286432, -0.8061985, -0.7620572, -0.7103157, -0.6477998, -0.5955697, 
    -0.5951464, -0.6819303, -0.8238249, -0.9706836, -1.118372, -1.186911, 
    -1.201462, -1.212952, -1.17127, -1.083314, -1.054212, -1.11292,
  -1.00138, -0.968715, -0.8843725, -0.788002, -0.6587377, -0.5151179, 
    -0.4385715, -0.4210749, -0.4430964, -0.5366511, -0.6671362, -0.7828262, 
    -0.9074194, -1.001055, -1.063067, -1.087204, -1.047898, -1.052373, 
    -1.154734, -1.217624, -1.163702, -1.11336, -1.143927, -1.168438, 
    -1.120961, -1.090378, -1.151137, -1.245733, -1.300453, -1.223337, 
    -1.079245, -1.069724, -1.249102, -1.37249, -1.358965, -1.370521, 
    -1.49098, -1.560235, -1.445863, -1.256426, -1.167706, -1.233021, 
    -1.379539, -1.503757, -1.505141, -1.432305, -1.352813, -1.332549, 
    -1.351348, -1.330564, -1.270668, -1.211521, -1.161895, -1.120245, 
    -1.089581, -1.062872, -1.103253, -1.131589, -1.150599, -1.128513, 
    -1.093438, -1.028936, -1.07573, -1.204994, -1.284584, -1.263686, 
    -1.261455, -1.306817, -1.287758, -1.336391, -1.513197, -1.67796, 
    -1.615362, -1.357794, -1.097589, -0.8703425, -0.7023571, -0.5953095, 
    -0.5184867, -0.4165013, -0.3254209, -0.4159319, -0.6568499, -0.78351, 
    -0.7499161, -0.6720841, -0.6063771, -0.65973, -0.8337209, -1.02669, 
    -1.078496, -1.069821, -1.044366, -0.9715137, -0.9107388, -0.9463185,
  -0.5860977, -0.4571915, -0.2570126, -0.06318116, 0.06198144, 0.08019423, 
    0.04881406, 0.05377817, 0.02039623, -0.08974361, -0.1824682, -0.2748835, 
    -0.3791642, -0.4484837, -0.5102186, -0.6080542, -0.7004044, -0.7728, 
    -0.8512993, -0.893487, -0.8427379, -0.7925916, -0.8198214, -0.8061986, 
    -0.6673474, -0.5864394, -0.6215141, -0.6391251, -0.5983374, -0.5551732, 
    -0.5576148, -0.6701143, -0.8308403, -0.8353326, -0.7551403, -0.7459772, 
    -0.7633924, -0.6895971, -0.6005344, -0.5635881, -0.5910294, -0.7379043, 
    -0.9273739, -0.990427, -0.8742325, -0.7783504, -0.7880671, -0.8192682, 
    -0.7934055, -0.7516251, -0.7689915, -0.784405, -0.7137017, -0.6157687, 
    -0.5631318, -0.5606253, -0.5788059, -0.5479467, -0.4419568, -0.4134414, 
    -0.5098119, -0.6821589, -0.8468072, -0.9105768, -0.857924, -0.8423638, 
    -0.8913221, -0.9029758, -0.8717744, -0.8793428, -0.7717094, -0.5424452, 
    -0.3392389, -0.1884091, -0.172133, -0.2497692, -0.3019986, -0.1811173, 
    -0.0001924038, 0.02674484, -0.1285775, -0.4310193, -0.7187312, 
    -0.7242324, -0.5282688, -0.4368296, -0.5040497, -0.63001, -0.7697561, 
    -0.8575816, -0.8276011, -0.7433723, -0.7218721, -0.6639459, -0.6097305, 
    -0.5883763,
  -0.2856584, -0.04112697, 0.2497096, 0.3883488, 0.4565289, 0.5235047, 
    0.5732934, 0.5848167, 0.510875, 0.4506373, 0.4006047, 0.2364445, 
    0.001792908, -0.1956029, -0.3393202, -0.5120902, -0.6029108, -0.5386367, 
    -0.4596326, -0.5066864, -0.5328262, -0.5277319, -0.5379858, -0.5456514, 
    -0.4602349, -0.3424778, -0.2248836, -0.119952, -0.08165431, -0.06656647, 
    -0.0528295, -0.06386471, -0.02852941, 0.05705023, 0.09562421, 0.09887934, 
    0.1663113, 0.2141464, 0.1164577, -0.0009577274, -0.03676486, -0.09776735, 
    -0.2216444, -0.2595024, -0.1793268, -0.09379625, -0.09036207, -0.1482882, 
    -0.1669407, -0.0977838, -0.1370084, -0.254668, -0.2287245, -0.06754208, 
    0.04660177, 0.08208346, 0.05737638, 0.05441403, 0.1337919, 0.08844638, 
    -0.07507896, -0.3014135, -0.3993461, -0.2341444, -0.03264689, 
    -0.07958698, -0.1929822, -0.1509576, -0.09402418, -0.04999709, 0.1357772, 
    0.303632, 0.2860377, 0.1973495, 0.2754095, 0.421031, 0.4925642, 
    0.5407414, 0.4830439, 0.2426628, 0.01772785, -0.007598162, -0.00295949, 
    0.05036139, 0.1523962, 0.1259151, -0.07537103, -0.2203908, -0.1960092, 
    -0.1590624, -0.1699836, -0.1687143, -0.1742325, -0.2685359, -0.3911922, 
    -0.4010391,
  0.3014185, 0.6419296, 0.9841175, 1.123685, 1.257556, 1.39932, 1.423946, 
    1.329381, 1.11667, 0.7794145, 0.4389846, 0.08273435, -0.173353, 
    -0.3183887, -0.4055634, -0.4075166, -0.3389291, -0.2147915, -0.1854783, 
    -0.2951463, -0.3854299, -0.3831837, -0.3517873, -0.226023, 0.04987288, 
    0.3630078, 0.5666862, 0.6886916, 0.7544632, 0.8214228, 0.8940139, 
    0.8665237, 0.8090369, 0.7913611, 0.7764846, 0.78459, 0.7670445, 
    0.7272333, 0.7745805, 0.7455925, 0.5217969, 0.269209, 0.1732943, 
    0.1353875, 0.1501501, 0.308125, 0.4910026, 0.5137405, 0.3035192, 
    0.2740757, 0.3752315, 0.3784379, 0.4517615, 0.5113155, 0.3866407, 
    0.2901564, 0.3411492, 0.4926465, 0.6585971, 0.533939, 0.250247, 
    0.1033559, 0.2326205, 0.5105176, 0.6779003, 0.5958855, 0.403193, 
    0.3128772, 0.3553576, 0.4199083, 0.4823432, 0.5431831, 0.6470249, 
    0.8218949, 1.074157, 1.618851, 1.896487, 1.277347, 0.6347688, 0.1508496, 
    0.1089063, 0.4151238, 0.6852409, 0.7524446, 0.644079, 0.357572, 
    0.04569006, -0.0458951, 0.02695656, 0.1260939, 0.1148961, 0.01709318, 
    -0.05323553, -0.1711884, -0.1777644, 0.06351161,
  0.6512406, 0.9924349, 1.331579, 1.498522, 1.622773, 1.523571, 1.220267, 
    0.8413931, 0.3303742, -0.07999337, -0.2318654, -0.2604787, -0.1511523, 
    -0.02758455, 0.02739584, 0.04223967, -0.01860023, -0.142347, -0.33486, 
    -0.3590951, -0.2421354, -0.03638995, 0.2677767, 0.4711621, 0.6822134, 
    0.9290882, 1.098652, 1.268525, 1.399596, 1.408418, 1.310241, 1.116914, 
    0.9871289, 0.9458202, 0.8591666, 0.7859405, 0.777884, 0.8651562, 0.96916, 
    0.6316763, 0.2029655, 0.01992494, 0.1261262, 0.2887562, 0.5489613, 
    0.7028838, 0.6901885, 0.5856314, 0.4989615, 0.5803579, 0.7961946, 
    0.811608, 0.7108756, 0.5535839, 0.3941764, 0.4952832, 0.7106803, 
    0.7975942, 0.7640494, 0.535257, 0.3887403, 0.4852084, 0.6869012, 
    0.7986201, 0.7557166, 0.6929885, 0.5704463, 0.4935094, 0.5781447, 
    0.6955602, 0.7468134, 0.8523308, 1.17873, 1.459313, 1.625736, 2.325507, 
    2.501825, 1.153958, 0.1558463, -0.01231772, 0.2972853, 0.6729199, 
    0.8189485, 0.5742872, 0.1889356, -0.1588997, -0.2346323, -0.02763343, 
    0.09279299, 0.07526362, 0.10653, 0.06237316, 0.04072595, 0.07069016, 
    0.1467972, 0.3733922,
  0.8128938, 1.179479, 1.466312, 1.739212, 1.857392, 1.384882, 1.037275, 
    0.6454134, 0.01756503, 0.02552414, 0.4800813, 0.8009146, 0.8681185, 
    0.7175324, 0.5444205, 0.227233, -0.1878223, -0.4375131, -0.4923308, 
    -0.2528614, 0.02969065, 0.2423209, 0.5118684, 0.6124869, 0.7737012, 
    1.174857, 1.408353, 1.515644, 1.542336, 1.529234, 1.349091, 0.8426141, 
    0.5567741, 0.6367872, 0.6651237, 0.748278, 0.7558465, 0.8504428, 
    0.6217806, 0.08864251, 0.0328645, 0.2731314, 0.1818228, 0.210664, 
    0.5271354, 0.4730663, 0.2263702, 0.2913281, 0.5250684, 0.8068879, 
    0.9047069, 0.6202505, 0.3182324, 0.2093782, 0.1492057, 0.2740917, 
    0.3453971, 0.3758169, 0.3769725, 0.2997753, 0.4213572, 0.589326, 
    0.7164584, 0.7487659, 0.6459991, 0.602868, 0.4675326, 0.5708692, 
    0.8448439, 0.8350292, 0.9516634, 1.184834, 1.337454, 1.53804, 1.818281, 
    2.319926, 1.751713, 0.4848661, 0.006562423, 0.2035026, 0.4137727, 
    0.5404166, 0.4083852, -0.04348624, -0.3537402, -0.2351366, -0.05774415, 
    0.04223967, -0.01537752, -0.00930655, 0.1316603, 0.06557953, 0.06990862, 
    0.2366732, 0.3180044, 0.4807487,
  0.7101269, 1.093899, 1.380455, 1.584102, 1.220463, 0.7194364, 0.5958041, 
    0.39722, 0.187552, 0.8290557, 1.292663, 1.207653, 0.9922718, 0.4580436, 
    0.09453452, -0.2773407, -0.6370738, -0.5726858, -0.4636523, -0.2068166, 
    0.007864594, 0.1301463, 0.4960971, 0.7140168, 0.9609562, 1.266897, 
    1.281383, 1.32554, 1.409866, 1.395772, 0.9360871, 0.3748889, 0.3782422, 
    0.6621126, 0.6924675, 0.6348015, 0.4678574, 0.1758008, -0.1949675, 
    -0.4609018, 0.01279615, 0.2163607, -0.04262364, 0.1970085, 0.5435252, 
    0.428421, 0.3023794, 0.4793164, 0.6247103, 0.5924839, 0.2770704, 
    -0.1030567, -0.2609018, -0.2769988, -0.36834, -0.2519011, -0.006311923, 
    0.2505728, 0.3227246, 0.1432649, 0.2904003, 0.4252148, 0.372757, 
    0.2720897, 0.1941275, 0.3355988, 0.4326527, 0.6177764, 0.7829621, 
    0.678177, 0.8389355, 1.007572, 1.076452, 1.265953, 1.419127, 1.267712, 
    0.2532749, -0.2234347, 0.06857415, 0.2207063, 0.234899, 0.240498, 
    0.1153677, 0.008515477, -0.1121874, -0.004651666, 0.06043625, 
    -0.06093419, -0.07301122, 0.1142772, 0.1643749, 0.03813794, 0.02820956, 
    0.02337557, 0.09684569, 0.3663607,
  0.7136259, 0.9439969, 1.020788, 1.004902, 0.7044144, 0.4556674, 0.1505404, 
    -0.09501648, 0.2056022, 1.250638, 1.405537, 0.8937361, 0.5327179, 
    0.04844064, -0.4206675, -0.6966924, -0.9134411, -0.8233858, -0.6953257, 
    -0.4974253, -0.2085904, 0.09025407, 0.5375516, 0.7619493, 0.8686876, 
    0.8925481, 0.9252634, 1.067582, 1.090629, 0.8133497, 0.2043324, 
    0.0343132, 0.4375194, 0.5831901, 0.2758007, 0.1968132, -0.0499804, 
    -0.2887011, -0.5414516, -0.5420541, -0.07078123, 0.1870141, 0.3378935, 
    0.7344429, 0.7346056, 0.3508978, 0.2356145, 0.333694, 0.1663761, 
    -0.2812955, -0.6430143, -0.7041309, -0.7599089, -0.7254201, -0.6477019, 
    -0.2308725, 0.1384145, 0.1256379, 0.04209302, -0.06737963, 0.119388, 
    0.1865754, 0.03546868, 0.005618408, 0.07160148, 0.369925, 0.5879263, 
    0.659606, 0.6077507, 0.6564323, 0.7946483, 0.7738957, 0.7745144, 
    0.7401071, 0.6546264, 0.3237019, -0.4313607, -0.2310351, 0.01194979, 
    -0.1869596, 0.001142502, 0.1136751, 0.05890614, 0.08016269, -0.1088021, 
    -0.3575814, -0.2127734, -0.1607391, -0.09692067, 0.07051099, -0.04622078, 
    -0.1226531, -0.0301888, -0.04978514, 0.1701529, 0.4791367,
  0.5486031, 0.545609, 0.4961295, 0.6630406, 0.5254745, 0.2515005, 
    -0.002584636, -0.100127, 0.2569205, 0.8281929, 0.9410195, 0.4390984, 
    0.07469416, -0.09880869, -0.7523568, -1.175403, -1.121774, -0.9351531, 
    -0.6333137, -0.3246548, 0.004137278, 0.2888374, 0.5655298, 0.6555526, 
    0.6582224, 0.7305527, 0.7523794, 0.5467644, 0.3852901, 0.2582712, 
    -0.03064537, 0.05731118, 0.2643912, 0.1957064, -0.07319033, -0.1473606, 
    -0.3925107, -0.633038, -0.6794076, -0.3982553, 0.01424384, 0.3308134, 
    0.5936232, 0.5939968, 0.392597, -0.02138424, -0.2391415, -0.2575333, 
    -0.6624482, -1.091989, -1.227324, -0.9032683, -0.8243946, -0.6463673, 
    -0.2231576, 0.1644075, 0.3019888, -0.09475593, -0.1399545, 0.01196607, 
    0.1545116, 0.1943066, 0.1421581, 0.2274609, 0.4256705, 0.6397168, 
    0.7275749, 0.7342481, 0.6234245, 0.5938346, 0.5557806, 0.450784, 
    0.4827824, 0.3593459, 0.2588248, 0.009785652, -0.3624806, 0.02630544, 
    0.003616512, -0.1984993, 0.05638339, 0.1947297, 0.1304557, 0.2035188, 
    -0.0004688501, -0.3434049, -0.2503222, -0.02581063, 0.04010734, 
    0.2057486, 0.1808301, 0.1617546, 0.2047559, 0.2237988, 0.3564482, 
    0.4293973,
  0.2618194, 0.08774757, 0.1521521, 0.4069042, 0.3557324, 0.01917639, 
    0.06347972, 0.3649772, 0.4639356, 0.3876166, 0.5508657, 0.2878931, 
    -0.04501635, -0.006588608, -0.734437, -1.076494, -0.8176403, -0.5275849, 
    -0.1749804, 0.103112, 0.3547072, 0.4473171, 0.4820011, 0.5397813, 
    0.5818222, 0.601028, 0.3339062, 0.03867435, 0.2012396, 0.1419301, 
    -0.1579394, -0.3034147, -0.3081348, -0.3431444, -0.4777801, -0.5881807, 
    -0.6241014, -0.5637658, -0.2458951, -0.02001643, -0.07885504, 0.01260042, 
    0.0373559, -0.06495523, 0.1234074, -0.3983042, -0.976136, -1.055531, 
    -1.425013, -1.425257, -1.122409, -0.5841277, -0.4694955, -0.3402963, 
    -0.04011727, 0.05892245, 0.1829947, -0.05457039, 0.03289706, 0.2726757, 
    0.2783723, 0.309134, 0.3635285, 0.4239779, 0.6141146, 0.7626009, 
    0.7009473, 0.6114289, 0.4984074, 0.4005561, 0.337291, 0.2619982, 
    0.2281275, 0.07713461, -0.07105827, -0.1398239, 0.1360061, 0.2231152, 
    -0.1980925, -0.1298633, 0.2376822, 0.2188345, -0.02039069, 0.06842765, 
    0.0177929, -0.3381967, -0.1538706, 0.225052, 0.3494172, 0.3816438, 
    0.2976106, 0.3475782, 0.3456569, 0.3294299, 0.3135607, 0.2578802,
  -0.05640984, -0.1948538, -0.1523733, -0.06464505, 0.1272655, 0.02689111, 
    0.1725292, 0.1836132, 0.03625, -0.000159502, 0.1879755, 0.2194531, 
    -0.2732715, -0.7880827, -1.299232, -0.9820932, -0.6233204, -0.3507781, 
    0.0793165, 0.2741896, 0.4605829, 0.2849801, 0.2003772, 0.4102731, 
    0.423245, 0.2742214, -0.02117229, -0.06386399, -0.01703787, -0.3540494, 
    -0.6364062, -0.7322885, -0.6759245, -0.5918425, -0.6180144, -0.566403, 
    -0.6393683, -0.7491667, -0.2017058, -0.2570605, -0.6600072, -0.6238737, 
    -0.5396448, -0.2836392, 0.05130506, -0.6649382, -1.353105, -1.229115, 
    -1.414906, -1.146384, -0.5485157, 0.05081701, 0.072106, -0.07255542, 
    0.1142447, 0.2879101, 0.4003124, 0.3416536, 0.4324902, 0.495446, 
    0.4095085, 0.402819, 0.4952995, 0.5457552, 0.593444, 0.5934602, 
    0.5899608, 0.4644234, 0.3693225, 0.3129749, 0.2629256, 0.2025251, 
    0.0556016, -0.0610652, -0.04739237, 0.02155256, 0.3288281, 0.1661164, 
    -0.1857715, -0.03295588, 0.1929882, 0.1174347, -0.07323903, 0.08672184, 
    -0.05614917, -0.1741016, 0.2841015, 0.4361848, 0.4315461, 0.459069, 
    0.362975, 0.3260608, 0.2546253, 0.2175972, 0.1974797, 0.1250515,
  -0.1765273, -0.1148255, -0.01337624, 0.1170117, 0.1446809, -0.1065724, 
    -0.08243501, -0.3011361, -0.2663379, -0.01404309, 0.03703117, 
    -0.006669998, -0.5275522, -0.9602669, -0.7972463, -0.1759897, -0.1869109, 
    -0.1858367, 0.1700065, 0.2358268, 0.2019401, -0.151071, -0.2020963, 
    0.02674484, -0.09353518, -0.2633431, -0.2908007, -0.164743, -0.1963184, 
    -0.4743945, -0.5122039, -0.3391896, 0.05928063, -0.04662752, -0.2866992, 
    -0.2640431, -0.4529916, -0.5252897, 0.01245427, -0.3099578, -0.7498341, 
    -0.5232227, -0.3648406, 0.1550325, 0.2601919, -0.3216602, -0.7208138, 
    -0.6068327, -0.7429655, -0.3500947, 0.3134147, 0.5237176, 0.3588248, 
    0.1859407, 0.1835806, 0.2963085, 0.2595247, 0.2366568, 0.286966, 
    0.2597689, 0.2826205, 0.3487663, 0.4120963, 0.391133, 0.431253, 
    0.3908558, 0.391881, 0.3056345, 0.2779651, 0.2472517, 0.1195989, 
    0.06526923, -0.02896881, -0.181654, -0.2100229, 0.1195021, 0.04956374, 
    0.1739942, 0.0003287792, 0.1317251, 0.09134433, 0.02905592, 0.002428308, 
    0.0883007, -0.1380177, -0.004602909, 0.3850455, 0.3823762, 0.3227897, 
    0.2012078, 0.1097689, 0.01515627, 0.03820276, 0.03530526, 0.01147723, 
    -0.06921983,
  -0.1479628, -0.1325819, -0.09687191, 0.1527864, 0.083955, -0.04024747, 
    -0.2082976, -0.4593881, -0.2481414, -0.1687305, -0.1039193, -0.1793588, 
    -0.3310027, -0.04682299, 0.231416, 0.3323436, -0.1084766, -0.3365852, 
    -0.1379688, -0.01601245, -0.03090502, -0.1879851, -0.2113249, -0.1363249, 
    -0.1662078, -0.1493621, 0.005211473, 0.02809554, -0.1585092, -0.3392872, 
    -0.2716602, -0.154961, 0.02340817, -0.1728485, -0.2875456, -0.1708138, 
    -0.1208463, -0.2372851, -0.2305794, -0.681312, -0.9063932, -0.1510384, 
    0.09761083, 0.473864, 0.4342318, 0.1323597, -0.04830396, -0.1846646, 
    -0.3057584, 0.08802414, 0.2850131, 0.1279653, 0.113854, 0.08432937, 
    -0.01355477, 0.1365917, 0.199759, 0.2579134, 0.2620637, 0.2358106, 
    0.2340853, 0.2505242, 0.3188508, 0.3107131, 0.2966173, 0.248245, 
    0.1912625, 0.2092314, 0.2288437, 0.2067571, 0.1436713, 0.0496769, 
    -0.005710602, -0.1038716, -0.07480145, 0.004153568, 0.07840484, 
    0.0528352, 0.07679355, 0.06347966, 0.08611971, 0.0665722, 0.105358, 
    0.1828482, 0.02889317, 0.1357942, 0.2447462, 0.2627799, 0.2450554, 
    0.0688346, 0.117793, 0.009508491, -0.01376629, -0.1181283, -0.1534641, 
    -0.1942196,
  -0.3311164, -0.2658496, -0.2054005, 0.1069694, 0.2391309, 0.1119661, 
    -0.08959621, -0.3002247, -0.2706186, -0.574362, -0.3923634, -0.1531218, 
    -0.2165006, 0.07791674, 0.1946485, 0.1952833, -0.008330226, -0.06788421, 
    0.07567045, 0.1796581, 0.1170605, 0.04710606, -0.0582325, -0.05445647, 
    0.09853834, 0.2094107, 0.4621776, 0.4165396, -0.0251433, -0.2192839, 
    0.07280591, -0.02367836, -0.204196, -0.2724907, -0.0744108, 0.1640006, 
    0.1351593, -0.0931282, -0.01607755, -0.06415701, -0.1425264, 0.2390007, 
    0.03076506, -0.1111621, -0.1440558, -0.3633268, -0.5309702, -0.543926, 
    -0.5316374, -0.3685514, -0.4777961, -0.5812466, -0.4813607, -0.5076628, 
    -0.4674772, -0.2911913, -0.1364063, -0.02019542, -0.03915691, 0.02212229, 
    0.09795234, 0.1280305, 0.1526236, 0.2526887, 0.2314323, 0.247806, 
    0.1869172, 0.158548, 0.06209636, -0.1007292, -0.1054659, -0.1287894, 
    -0.2158005, -0.4271941, -0.3454553, 0.00475578, 0.004462808, -0.05660489, 
    -0.02664071, -0.006653711, -0.007744133, 0.05796218, 0.1139843, 
    0.2717317, 0.1360058, -0.0155077, 0.1112337, 0.3058951, 0.2189485, 
    0.09331363, 0.1477734, -0.003414631, -0.07859397, -0.2075979, -0.266989, 
    -0.3535448,
  -0.06422204, -0.063034, -0.03176766, 0.1453808, 0.1223176, -0.03596687, 
    -0.01741219, -0.02553393, -0.05725592, -0.2706512, -0.1253549, 
    0.02018559, -0.2128549, -0.2664688, 0.02930021, 0.2933955, 0.3072625, 
    0.352103, 0.4125358, 0.35194, 0.265856, 0.1304069, -0.03005856, 
    -0.1069954, 0.02975577, 0.1337596, 0.2365266, 0.01894849, -0.2509896, 
    -0.3427378, 0.001956299, -0.07284838, -0.05556324, 0.09669828, 
    -0.02548552, -0.04097998, -0.02856135, 0.08341783, 0.4278029, 0.7301784, 
    0.3747261, 0.2990432, 0.2132189, 0.07593107, 0.03393888, -0.05092454, 
    -0.1034639, -0.1122367, -0.1881809, -0.2061331, -0.175746, -0.2421196, 
    -0.3486462, -0.4133272, -0.3946912, -0.4530737, -0.4539521, -0.3319631, 
    -0.2564261, -0.1518685, -0.08551097, 0.05986667, 0.04866862, 0.1091666, 
    0.1204948, 0.1877311, 0.1290559, 0.1193066, 0.1401399, 0.07073885, 
    0.06055009, -0.02498055, -0.2320118, -0.4148406, -0.3857553, -0.1122201, 
    -0.03134447, -0.06796557, -0.03827807, 0.002395809, 0.1577343, 0.1729361, 
    0.06748372, -0.2024057, -0.06415677, -0.1500626, 0.06076121, 0.1730177, 
    0.101517, 0.03034171, -0.009209059, -0.04132169, -0.002128899, 
    -0.02908206, -0.04055655, 0.005651116,
  0.1198926, 0.2357616, 0.1276074, 0.03773105, 0.06196606, 0.04121411, 
    0.06175447, 0.03813797, 0.05610663, -0.06728196, -0.2317189, 0.05976892, 
    0.06486315, -0.1739559, -0.1798966, 0.0840528, 0.2613478, 0.341247, 
    0.4031771, 0.3394564, 0.2315462, -0.04454434, -0.03437173, -0.001998663, 
    0.00654608, 0.03895175, 0.1566113, -0.1323373, -0.5021946, -0.5391574, 
    -0.07787764, 0.002916589, -0.01184577, 0.08421493, -0.1051083, 
    -0.07592487, -0.04719806, 0.2114782, 0.1286653, 0.2086937, 0.1938663, 
    0.2514837, 0.3283391, 0.4416041, 0.5110214, 0.5773787, 0.6065619, 
    0.638365, 0.7232122, 0.7531114, 0.7247427, 0.5598502, 0.3989291, 
    0.2012079, -0.02496409, -0.142233, -0.2387824, -0.2708141, -0.3113574, 
    -0.3080696, -0.3569467, -0.2986785, -0.2906543, -0.2839323, -0.2524871, 
    -0.09006843, -0.01664722, 0.08572911, 0.1565787, 0.1501171, 0.1900259, 
    0.1780143, 0.03582674, 0.07529628, 0.0528841, -0.0472787, -0.01495451, 
    0.1789908, 0.1814322, 0.2780468, 0.3814812, 0.06064785, -0.1488085, 
    -0.2260861, -0.01591539, 0.05382681, 0.09747934, 0.02010369, -0.01899123, 
    -0.01313162, 0.006350994, -0.02680346, -0.08145845, -0.06453127, 
    -0.1426075, -0.0322721,
  0.3259311, 0.2996447, 0.178991, 0.04329753, -0.03036797, -0.03277671, 
    0.02497077, 0.1069368, 0.2061555, 0.1348176, -0.22236, -0.1015267, 
    -0.02209969, -0.211748, -0.4100721, -0.1317358, 0.1719913, 0.3259141, 
    0.4444371, 0.4680208, 0.3790722, -0.1127083, -0.09124032, -0.02349925, 
    -0.1650521, -0.3354622, 0.008596927, -0.06392911, -0.4228652, -0.71419, 
    -0.4687145, -0.07737303, -0.06827474, -0.1012175, -0.1113582, 0.1347029, 
    0.1043649, 0.1928899, 0.1852565, 0.2247581, 0.2617865, 0.2727237, 
    0.1805525, 0.2093122, 0.283824, 0.3432474, 0.4186058, 0.5527043, 
    0.7173686, 0.7989283, 0.8035831, 0.7788923, 0.7273459, 0.5514998, 
    0.3439314, 0.2352726, 0.06476498, -0.03464913, -0.1631806, -0.2950006, 
    -0.3300428, -0.3512669, -0.3464164, -0.3561001, -0.2860482, -0.1392221, 
    -0.06361973, -0.01448256, -0.029603, 0.03001618, -0.0321908, -0.01736343, 
    0.2247268, 0.4166209, 0.2440131, 0.0772981, 0.184671, 0.5106804, 
    0.5432329, -0.04366541, -0.1581028, 0.008352041, 0.5277696, 0.3772483, 
    0.3146832, 0.2437525, 0.1726911, 0.1543806, 0.1390324, 0.1001329, 
    0.1115267, 0.05600917, 0.01429355, 0.1795443, 0.1729199, 0.198099,
  0.5782096, 0.5494986, 0.3863313, 0.1778352, -0.0007454157, 0.01061516, 
    0.07350577, 0.1536328, 0.2177768, 0.2120637, 0.0001170039, -0.2387987, 
    -0.2681119, -0.2319793, -0.397963, -0.270359, 0.02257705, 0.3827169, 
    0.5358748, 0.6168003, 0.6280143, 0.2903353, 0.2290559, 0.1525585, 
    0.08603823, -0.2706186, 0.06408167, 0.0198437, -0.1638639, -0.5228651, 
    -0.9129202, -0.5298963, -0.2747693, -0.04620445, -0.1146297, 0.07744408, 
    0.2119005, 0.2371769, 0.2936385, 0.2640324, 0.2285993, 0.2238953, 
    0.1684594, 0.1174178, 0.07384682, 0.07794809, 0.1203966, 0.1718616, 
    0.1761909, 0.2680368, 0.297936, 0.3093619, 0.2687364, 0.3076525, 
    0.2108755, 0.1309271, 0.1341667, 0.03349924, 0.01665354, -0.0462532, 
    -0.126348, -0.1509733, -0.08948278, -0.06438541, -0.06907272, -0.1304665, 
    -0.08145881, 0.04572296, 0.05364919, 0.1938021, 0.1841016, -0.01788402, 
    0.09962821, 0.2851267, -0.002633333, -0.1173143, -0.1901665, -0.1872046, 
    -0.3144999, -0.2211885, 0.1088083, 0.3649116, 0.3835311, 0.2893088, 
    0.2479515, 0.1647325, 0.1296411, 0.07246351, 0.05312729, 0.07680941, 
    0.2043481, 0.3454947, 0.3243685, 0.2423209, 0.3185904, 0.4966342,
  0.2857943, 0.5398799, 0.5215366, 0.37274, 0.1381373, -0.03860426, 
    -0.09604216, -0.00338316, 0.007150173, -0.0746069, -0.1634733, 
    -0.2084603, -0.2419889, -0.356312, -0.5211068, -0.3583305, -0.1411111, 
    0.2109723, 0.5280461, 0.7483587, 0.4967805, 0.5098176, 0.7004427, 
    0.3147981, 0.1507844, 0.09557617, 0.149629, -0.03796893, -0.2516243, 
    -0.6211882, -0.965817, -0.8216281, -0.6887989, -0.4809055, -0.4273736, 
    -0.2537732, -0.04802799, 0.07498646, 0.2391465, 0.289032, 0.3051622, 
    0.2254908, 0.09617758, -0.01746178, -0.06088614, -0.03726959, 
    -0.07307696, -0.0332334, 0.05534077, 0.1783228, 0.1841331, 0.2000837, 
    0.1232772, 0.1240101, 0.02301788, -0.1234841, -0.07481813, -0.1182098, 
    -0.09996462, -0.01882839, 0.01989269, -0.01860046, -0.04023123, 
    -0.02561522, 0.01126623, -0.009176731, -0.09426832, -0.1961727, 
    -0.1243131, 0.2035514, 0.6736685, 0.8727086, 0.4260614, -0.08749723, 
    -0.3181272, -0.3844533, -0.3640432, -0.4749322, -0.2763476, 0.03496432, 
    0.09407878, 0.2107785, 0.2804878, 0.3411155, 0.2260764, 0.1481466, 
    0.09935188, -0.02960253, -0.09499979, -0.1322055, -0.1019988, 0.1462603, 
    0.2564325, -0.05554652, -0.2164037, -0.05929041,
  -0.07507896, 0.1317737, 0.1794946, 0.2920434, 0.3210475, 0.08465409, 
    -0.1531062, -0.2086725, -0.1023731, -0.07590818, -0.1645484, 0.004169941, 
    -0.1408008, -0.4439585, -0.5569791, -0.3812143, -0.2560188, -0.05600357, 
    0.4675159, 0.7286005, 0.3361518, 0.7934115, 1.256887, 0.5141141, 
    -0.03733408, 0.1246777, 0.07962567, -0.305433, -0.9645314, -1.615768, 
    -1.531768, -0.881963, -0.6059375, -0.7354947, -0.7804335, -0.5241184, 
    -0.3246067, -0.1762016, 0.02402616, 0.1579456, 0.2096381, 0.2577503, 
    0.1435413, -0.08064508, -0.2313447, -0.2233858, -0.1778622, -0.1521297, 
    -0.1341283, 0.00945878, 0.1287298, 0.1594911, 0.0618515, -0.05339932, 
    -0.07992935, -0.2414365, -0.3925757, -0.3308246, -0.3518038, -0.3269184, 
    -0.2311821, -0.1812797, -0.1725392, -0.2311168, -0.2561817, -0.1574345, 
    -0.1726532, -0.3175426, 0.01081085, 0.1555533, 0.1044791, 0.002444744, 
    -0.04096353, -0.3307428, -0.5596814, -0.5715625, -0.4270639, -0.3762826, 
    -0.3309863, -0.1324676, -0.03949869, 0.1199903, 0.2052934, 0.1736689, 
    0.06826448, -0.03795314, -0.1893208, -0.2563291, -0.395586, -0.4752893, 
    -0.5730267, -0.4742966, -0.08108473, -0.05048561, -0.2066708, -0.2574518,
  -0.2361627, 0.0359571, 0.131644, 0.1495957, 0.1711295, -0.07242513, 
    -0.255433, -0.4701471, -0.5664363, -0.3881645, -0.2103152, 0.03929353, 
    0.196927, 0.0696972, -0.1862598, -0.3418097, -0.5257455, -0.3272922, 
    0.1924503, 0.118232, -0.01555705, 0.508483, 1.160794, 1.083824, 
    0.1808453, -0.1936165, -0.08936858, 0.09157228, -0.291387, -1.230205, 
    -1.638831, -1.105921, -0.7233528, -0.9204232, -0.8824023, -0.6972623, 
    -0.5851207, -0.3876598, -0.2379692, -0.02571297, 0.03983092, 0.09709001, 
    0.06266606, -0.06376624, -0.2218879, -0.4269986, -0.5020641, -0.444707, 
    -0.3619434, -0.1868947, 0.03060174, 0.0898304, 0.08875608, -0.001673698, 
    -0.06796598, -0.2397106, -0.4633923, -0.4749811, -0.4694963, -0.3720188, 
    -0.3529761, -0.3218238, -0.2368793, -0.2661586, -0.2814584, -0.2358036, 
    -0.11235, 0.01531839, 0.08760089, 0.1827018, -0.1292936, -0.3700975, 
    -0.1853158, -0.1786914, -0.5719533, -0.7756153, -0.6834277, -0.4567026, 
    -0.2815235, -0.02325529, 0.1080924, 0.0586783, 0.1018587, 0.1601596, 
    0.1233432, -0.06137359, -0.2850232, -0.3359675, -0.6167779, -0.7463832, 
    -0.8333459, -0.9073687, -0.4646947, -0.29072, -0.3433077, -0.313669,
  -0.1993301, -0.04350281, 0.08748686, 0.05529296, 0.07698894, -0.08542985, 
    -0.1795703, -0.3489879, -0.7130179, -0.5488415, -0.2683244, -0.2563607, 
    -0.1411427, 0.007148445, 0.09708971, -0.05253583, -0.4369109, -0.2660122, 
    -0.134974, -0.2647429, -0.1176888, 0.1135124, 0.3312209, 0.4837599, 
    0.1756537, 0.01437485, 0.1436881, 0.2278345, -0.3086073, -0.7845996, 
    -1.237952, -1.344854, -1.014808, -1.11196, -0.7591928, -0.5637337, 
    -0.5308887, -0.3150684, -0.2939258, -0.1613249, -0.1351205, -0.1118132, 
    -0.0363574, -0.04205418, 0.0126009, -0.1088836, -0.4206999, -0.5316536, 
    -0.5049772, -0.4759083, -0.2329882, -0.04190743, -0.1082816, -0.2268524, 
    -0.2450814, -0.367754, -0.5502738, -0.5914193, -0.6029751, -0.4816208, 
    -0.4270477, -0.3294082, -0.2324684, -0.2871881, -0.3727508, -0.3916297, 
    -0.1357069, -0.0789355, -0.06038094, -0.008281231, 0.3195181, 0.3936066, 
    0.1927278, 0.02340812, -0.2504036, -0.5067676, -0.5914519, -0.4751107, 
    -0.2343555, 0.05501619, 0.127054, 0.04800122, 0.1170605, 0.07132478, 
    -0.06492198, -0.258965, -0.473483, -0.5289842, -0.726397, -0.8578749, 
    -1.013066, -1.16082, -0.7297502, -0.408314, -0.3146126, -0.1748831,
  -0.03531575, -0.06682634, 0.06360996, 0.1934439, 0.328942, 0.18319, 
    0.06302401, -0.1466602, -0.6909148, -0.7031053, -0.4076954, -0.4413868, 
    -0.4865527, -0.2853971, -0.06012052, -0.1464324, -0.3234343, -0.374525, 
    -0.2650358, -0.01873052, 0.1826029, -0.0413053, -0.3457488, -0.4015919, 
    -0.4938929, -0.01630497, 0.3809115, -0.1237612, -0.4519012, -0.0744431, 
    -0.004163504, -0.3743457, -0.5166798, -0.7229785, -0.7103646, -0.5741992, 
    -0.5563445, -0.3611296, -0.2714975, -0.2481414, -0.275599, -0.2558562, 
    -0.2353322, -0.3367646, -0.1616343, 0.06351227, -0.08466476, -0.2995086, 
    -0.3660288, -0.4067351, -0.2715951, -0.03723639, -0.06596357, -0.2555631, 
    -0.3526823, -0.5710254, -0.8471323, -0.8844532, -0.7832813, -0.6320931, 
    -0.5205209, -0.4497038, -0.3269012, -0.1591287, -0.2741175, -0.3094053, 
    -0.09143543, 0.05394198, 0.05804354, 0.01658846, 0.2640657, 0.423164, 
    0.1632519, 0.003160732, -0.09934577, -0.263685, -0.3578907, -0.4023569, 
    -0.42625, -0.3145153, -0.07219744, 0.143281, 0.1328319, -0.09028018, 
    -0.2436817, -0.3436329, -0.5073861, -0.6427051, -0.8581999, -0.9798472, 
    -0.9946098, -1.136098, -0.9519992, -0.6567843, -0.2892057, 0.01383775,
  0.2240102, 0.3584176, 0.413561, 0.3352245, 0.4175161, 0.424873, 0.2911816, 
    -0.03886402, -0.6546518, -0.7834604, -0.422946, -0.308737, -0.3644825, 
    -0.2519337, -0.2285286, -0.3341603, -0.4618293, -0.5279915, -0.48875, 
    -0.2536101, 0.02360344, -0.3465947, -0.3995085, -0.2413225, -0.4554989, 
    -0.5057588, -0.3946917, -0.1454401, 0.1057486, 0.1611688, 0.2308946, 
    0.1161817, 0.1296097, -0.03668356, -0.1282036, -0.03748035, -0.1974577, 
    -0.1384245, 0.02348951, 0.00224936, -0.0289681, -0.03468084, -0.08064437, 
    -0.1286588, -0.1319797, -0.07948971, -0.026088, -0.01059294, -0.0134244, 
    -0.03780568, -0.02633107, 0.02687502, 0.03789377, -0.1048959, -0.2967416, 
    -0.5671355, -0.9141896, -1.150583, -1.063604, -0.8838999, -0.6313446, 
    -0.3797169, -0.2644823, -0.05588937, 0.02217054, -0.0333463, 
    -0.005677104, 0.05332349, 0.1555046, 0.2692253, 0.3194856, 0.2756217, 
    0.1304719, 0.04499018, -0.06069016, -0.09239591, -0.04340503, 0.05264008, 
    0.126338, 0.009296894, -0.115768, -0.01192713, 0.236315, 0.2833033, 
    -0.05920959, -0.480238, -0.6891403, -0.8874642, -1.163897, -1.344658, 
    -1.315199, -1.047507, -0.7229302, -0.5790501, -0.3155566, 0.01291007,
  0.2115103, 0.4729198, 0.6237334, 0.6828485, 0.7822946, 0.7470083, 
    0.5585644, 0.4240266, -0.1150357, -0.6679006, -0.5099741, -0.4554004, 
    -0.3719693, -0.349232, -0.2245086, -0.1984181, -0.2520314, -0.3872851, 
    -0.5774707, -0.41445, -0.2248182, -0.2032363, -0.1414523, -0.05945313, 
    -0.1854625, -0.3036592, -0.3310027, -0.3017221, -0.2758105, -0.184974, 
    -0.1423144, 0.1032261, 0.2995479, 0.2917027, 0.3127964, 0.4047887, 
    0.2102408, 0.3096548, 0.4220895, 0.3529981, 0.4613476, 0.4591014, 
    0.3263865, 0.2430856, 0.1710474, 0.1332219, 0.1223981, 0.1250513, 
    0.1094587, 0.1399274, 0.3299179, 0.43747, 0.3263049, 0.1774774, 
    0.003714442, -0.2913215, -0.6555142, -1.027113, -1.082679, -1.001689, 
    -0.8248665, -0.4016244, -0.1093394, -0.01445007, 0.1133657, 0.2901236, 
    0.2623242, 0.09111646, 0.1377147, 0.3827995, 0.5363964, 0.5695996, 
    0.5857291, 0.5049024, 0.3282747, 0.3917675, 0.5217968, 0.5749381, 
    0.6906119, 0.6931672, 0.5564806, 0.4676299, 0.4977241, 0.4979839, 
    0.1466331, -0.3104146, -0.5838356, -0.8640761, -1.158948, -1.517803, 
    -1.693584, -1.307956, -0.7437793, -0.4087858, -0.2273732, -0.04745775,
  0.2144563, 0.2886589, 0.4693232, 0.755602, 0.9513215, 0.8247917, 0.5230664, 
    0.7668326, 0.6453646, 0.09248376, -0.2961718, -0.2301236, -0.09255862, 
    0.06295896, 0.1416536, 0.09359042, -0.01420581, 0.09284163, 0.4510612, 
    0.6541209, 0.3934277, 0.3515169, 0.5535839, 0.4804719, 0.6028841, 
    0.7707715, 0.6373245, -0.06003922, -0.2844369, -0.223532, -0.413636, 
    -0.2643523, 0.02036452, 0.06616545, 0.03556645, 0.1033232, 0.1409539, 
    0.2727897, 0.4800162, 0.5527214, 0.6718132, 0.8029491, 0.846569, 
    0.5941929, 0.3567252, 0.3879423, 0.3538277, 0.3701034, 0.4286809, 
    0.3475935, 0.4190125, 0.5749211, 0.5472195, 0.4785182, 0.2943878, 
    -0.02607155, -0.2497041, -0.6243458, -0.9109018, -0.8639951, -0.8251109, 
    -0.6140924, -0.1083137, 0.2526237, 0.2629751, 0.2021679, 0.3797557, 
    0.3978547, 0.1510611, 0.2818716, 0.4131867, 0.476289, 0.5529166, 
    0.5672233, 0.3954622, 0.3997916, 0.4897493, 0.664668, 0.9040722, 
    0.9865429, 0.935371, 0.8387402, 0.7895703, 0.8099475, 0.5986514, 
    0.1007671, -0.4086893, -0.8333149, -1.216144, -1.58154, -1.673158, 
    -1.365524, -0.9216601, -0.4414031, -0.01824227, 0.1474316,
  0.26055, 0.4655633, 0.6187698, 0.7024934, 0.9067904, 0.7024771, 0.2996451, 
    0.26055, 0.4140006, 0.36667, 0.2009798, 0.3225945, 0.3192741, 0.02471021, 
    0.0167675, 0.1781445, 0.2141145, 0.31361, 0.7611361, 1.076891, 0.8486198, 
    0.6476105, 0.5896354, 0.3906445, 0.2438183, 0.3806347, 0.3299836, 
    -0.1565886, -0.08562505, 0.1047558, -0.04620451, -0.1107878, 0.1145378, 
    0.2144401, 0.1796092, 0.0970248, 0.003485918, 0.06992507, 0.2836295, 
    0.7048534, 0.6192253, 0.5453808, 0.7646841, 0.7495149, 0.5423373, 
    0.4900746, 0.3976591, 0.3415229, 0.4091988, 0.3634629, 0.4022977, 
    0.4938014, 0.4067571, 0.341783, 0.104104, -0.1855114, -0.1565399, 
    -0.2320933, -0.6526017, -0.7294736, -0.6688449, -0.7031391, -0.3140602, 
    0.1387072, 0.3714552, 0.07495451, 0.07734716, 0.2237988, 0.1637077, 
    0.2052605, 0.3093782, 0.2243521, 0.2297558, 0.4008658, 0.5126334, 
    0.4264843, 0.2444368, 0.2480501, 0.6336458, 0.7907423, 0.8824576, 
    1.00487, 1.005814, 1.047204, 1.015465, 0.6610217, 0.2007999, -0.2872536, 
    -0.9306133, -1.503415, -1.646172, -1.462464, -1.15003, -0.5687956, 
    0.0406934, 0.2623404,
  0.06715816, 0.277054, 0.2605664, 0.2890331, 0.6329623, 0.6570832, 
    0.3010774, -0.02694994, -0.03660154, 0.04839185, 0.1066438, 0.1948925, 
    0.18, -0.08697598, -0.3708464, -0.1906218, 0.2103222, 0.4768912, 
    0.7076855, 1.087048, 1.323978, 1.090905, 0.7167675, 0.3550487, 0.1817903, 
    0.2989615, 0.1646191, -0.194707, -0.1821257, 0.02477539, 0.08646166, 
    0.009394526, 0.007050991, 0.04515302, 0.1051791, 0.03704745, 0.0300163, 
    0.106822, 0.2514997, 0.6820014, 1.031758, 1.012113, 0.917272, 0.9340853, 
    0.9515983, 0.9399284, 0.8528513, 0.8457383, 0.8191758, 0.6410346, 
    0.5374377, 0.5491076, 0.4810901, 0.4486194, 0.07864881, -0.4786916, 
    -0.5528941, -0.3868625, -0.5199029, -0.6798801, -0.5676408, -0.4421852, 
    -0.2864561, 0.03603792, 0.4013376, 0.1156772, 0.05838549, 0.1076692, 
    0.2253937, 0.4190135, 0.3763703, 0.1395051, -0.03888023, -0.1607226, 
    0.05306306, 0.2150585, 0.2691275, 0.2590852, 0.1828971, 0.1437858, 
    0.4670929, 0.8342642, 1.030944, 1.140368, 1.123555, 0.923017, 0.5875351, 
    0.07544208, -0.6694477, -1.298939, -1.509991, -1.531849, -1.330937, 
    -0.738636, -0.08533239, 0.08174169,
  0.05112576, 0.1634631, 0.1944206, 0.254593, 0.3868032, 0.431888, 0.2334015, 
    -0.09556973, -0.2293425, -0.227601, -0.177422, -0.08248377, -0.0572722, 
    -0.2062794, -0.4178677, -0.4311817, -0.1754363, 0.1488802, 0.3235058, 
    0.5055045, 0.9341667, 1.239798, 1.071032, 0.7637404, 0.6503614, 
    0.4905794, 0.3582226, 0.1444531, 0.07176429, 0.0773958, 0.01460302, 
    -0.06552386, -0.06633782, -0.07843137, -0.2025688, -0.1992154, 
    0.05342126, -0.05139649, -0.3443332, -0.9491668, 0.4108591, 1.290677, 
    1.442582, 1.514391, 1.773587, 1.735111, 1.408109, 1.331986, 1.306481, 
    1.017907, 0.7231314, 0.6606313, 0.7632843, 0.7977406, 0.5778354, 
    0.185957, 0.01741838, -0.047019, -0.3892229, -0.8072243, -0.7618632, 
    -0.3603492, 0.04269528, 0.04087245, 0.02609384, 0.03419924, 0.09829426, 
    0.1226432, 0.2309602, 0.2783724, 0.204593, 0.1637076, 0.1019075, 
    0.09393227, 0.06666988, 0.1127474, 0.2192414, 0.2767772, 0.2235708, 
    0.1384474, -0.2350553, 0.03504539, 0.1988149, 0.745332, 0.9960318, 
    1.040531, 0.9059927, 0.5807806, -0.009323359, -0.6146457, -0.9868305, 
    -1.21541, -1.290426, -1.004798, -0.4406378, -0.06379843,
  -0.1474901, -0.1498665, 0.0554558, 0.1832715, 0.3106477, 0.40194, 
    0.3964224, 0.1703483, -0.09524423, -0.1391082, -0.08819687, -0.1043916, 
    -0.2292776, -0.3307258, -0.375127, -0.3705862, -0.3642221, -0.2622364, 
    -0.1199514, 0.1148471, 0.4598828, 0.7622101, 0.8340847, 0.6446643, 
    0.398701, 0.211071, 0.1264194, 0.08302718, 0.07807937, 0.07184563, 
    0.08659178, 0.0926466, 0.09704137, -0.009339571, -0.3896129, -0.4946423, 
    -0.200843, -0.2702444, -0.5412407, -1.292006, -0.7607069, 0.1433303, 
    0.6030632, 1.25666, 2.155195, 2.603144, 2.401127, 2.085908, 1.858743, 
    1.530081, 1.205911, 1.034004, 0.8983755, 0.726468, 0.4967806, 0.2832716, 
    0.2042348, 0.1532905, -0.0949192, -0.3950169, -0.358103, 0.08358026, 
    0.1366081, 0.1204134, 0.04575527, 0.05841804, 0.1718295, 0.1873079, 
    0.09204419, 0.06938794, 0.1655305, 0.289147, 0.4017773, 0.5010288, 
    0.5348178, 0.2879264, 0.2070832, 0.1925324, 0.2784536, 0.2143422, 
    -0.162334, -0.7209611, -1.147003, -0.5167451, -0.1015918, 0.3446483, 
    0.8380566, 1.06055, 0.7701528, 0.1977901, -0.2255988, -0.3836555, 
    -0.4390435, -0.4932747, -0.4206831, -0.2725552,
  -0.05222678, -0.06581712, -0.04565096, 0.1254096, 0.2849315, 0.3415559, 
    0.2411978, 0.06789052, -0.1328419, -0.2089975, -0.1718556, -0.1469207, 
    -0.2495249, -0.3107393, -0.279375, -0.1945443, -0.2344207, -0.3397918, 
    -0.4249967, -0.2385061, 0.0512892, 0.3063346, 0.4689158, 0.3893585, 
    0.2527212, 0.1615592, 0.08480155, -0.01501954, -0.1337206, -0.1850553, 
    -0.2037566, -0.192461, -0.1235484, -0.1214813, -0.2279266, -0.3823371, 
    -0.4284315, -0.5612926, -0.6936982, -1.125371, -1.259892, -0.7666152, 
    -0.2370903, 0.207978, 0.5223331, 1.897008, 2.388121, 2.628908, 2.748082, 
    2.668477, 2.316149, 1.859492, 1.415401, 1.013675, 0.4430534, -0.03412771, 
    -0.2436492, -0.2566699, -0.2002243, -0.1060514, 0.1282748, 0.05877614, 
    0.04653645, -0.0088346, 0.02490562, 0.1246126, 0.1846549, 0.1143424, 
    0.03616855, 0.05421867, 0.1568716, 0.1947134, 0.1712924, 0.2441928, 
    0.3805531, 0.435778, 0.4238964, 0.3399934, 0.3297396, 0.1804229, 
    -0.1393359, -0.741436, -1.057712, -0.7177224, -0.8235815, -0.5145966, 
    0.03945625, 0.6286978, 0.8539095, 0.606595, 0.2055209, -0.07874012, 
    -0.1720021, -0.172523, -0.1072564, 0.005422831,
  -0.03038406, -0.2356415, -0.2281055, -0.1694466, 0.01653969, 0.2158072, 
    0.1731314, 0.07490551, -0.05056646, -0.1209604, -0.1188771, -0.1611621, 
    -0.219463, -0.2875131, -0.3393523, -0.3388966, -0.3122364, -0.3211069, 
    -0.3440724, -0.2847625, -0.1669726, -0.03521812, 0.04018879, 0.08029306, 
    0.09980798, 0.07905602, 0.04803383, 0.003274739, -0.07148117, -0.1421191, 
    -0.2190724, -0.2404428, -0.186504, -0.1156381, -0.1220834, -0.2714485, 
    -0.5206836, -0.7696258, -1.049835, -1.308363, -1.378464, -1.263165, 
    -0.9891412, -0.651511, -0.2587535, 0.1474471, 0.5184278, 0.4418001, 
    0.7927928, 1.203844, 1.515172, 1.532912, 1.580309, 1.052868, 0.5375521, 
    0.1331086, -0.05852547, -0.1609343, -0.08821303, -0.1080371, -0.1341275, 
    -0.1502734, -0.1385709, -0.07813805, -0.01231781, 0.03927726, 0.08175775, 
    0.08800775, 0.07516593, 0.05781568, 0.01982731, 0.03945649, 0.1052605, 
    0.2099317, 0.3357292, 0.3962598, 0.4501657, 0.4204458, 0.4089552, 
    0.2314975, 0.05446243, -0.1514614, -0.2209764, -0.2315722, -0.5662079, 
    -0.7237608, -0.5714004, -0.08917308, 0.4304392, 0.7591501, 0.7597525, 
    0.5772655, 0.3541372, 0.2787467, 0.2778352, 0.1851921,
  0.1811391, -0.3107717, -0.5924282, -0.4457, -0.3260872, -0.1577115, 
    -0.04060549, 0.05433255, 0.0896028, 0.1112988, 0.07122707, 0.005146444, 
    -0.1160938, -0.2401171, -0.3644172, -0.4346648, -0.3936654, -0.3213022, 
    -0.2109831, -0.08235359, 0.02179682, 0.09694338, 0.1559116, 0.1591667, 
    0.1598991, 0.1283073, 0.09785485, 0.03079748, -0.08472989, -0.222295, 
    -0.3824674, -0.4678516, -0.4863574, -0.5326791, -0.5673308, -0.6419077, 
    -0.7231901, -0.7434701, -0.8149058, -0.9664193, -1.292543, -1.628871, 
    -1.529538, -1.286374, -1.011748, -0.7874485, -0.5629365, -0.1493788, 
    0.4486194, 1.124955, 1.595805, 1.442548, 1.559948, 1.117468, 0.7048208, 
    0.4263216, 0.2047395, 0.0786653, 0.03764963, 0.03143215, 0.04489243, 
    0.04619458, 0.04601556, 0.07500318, 0.128942, 0.1208365, 0.08825187, 
    0.09090486, 0.1039582, 0.1072949, 0.1641958, 0.2422394, 0.2886751, 
    0.2770869, 0.2471876, 0.2639682, 0.3354686, 0.4266471, 0.3464551, 
    0.1981153, 0.1104195, 0.03872418, 0.06362629, 0.08839837, 0.001354069, 
    -0.1924608, -0.3730607, -0.5544238, -0.06956053, 0.3705926, 0.469583, 
    0.9160028, 1.218314, 1.241833, 1.040595, 0.717386,
  0.7114453, 0.2342969, -0.2144988, -0.5297008, -0.7798305, -0.6582322, 
    -0.6116827, -0.4448856, -0.2130663, -0.008232713, 0.1638867, 0.231481, 
    0.1309766, 0.01989251, -0.1185515, -0.2574512, -0.3247526, -0.2494761, 
    -0.1334115, -0.006474689, 0.1045767, 0.1425326, 0.1044466, 0.08362913, 
    0.1075869, 0.1875682, 0.1675814, 0.1043813, -0.0278614, -0.206019, 
    -0.4191701, -0.5609018, -0.6036915, -0.6170541, -0.6208465, -0.7072885, 
    -0.6839161, -0.6557586, -0.6718067, -0.784502, -0.9602343, -1.047051, 
    -1.090036, -1.044121, -0.9636198, -0.9048634, -0.8356901, -0.6500462, 
    -0.2516084, 0.3265812, 0.6658065, 0.8099632, 0.8054063, 0.7134311, 
    0.5871778, 0.4962109, 0.4399121, 0.355407, 0.3016469, 0.2650749, 
    0.2533072, 0.2531933, 0.1918652, 0.1463899, 0.08423173, -0.001152456, 
    -0.08529955, -0.1170378, -0.07081388, 0.01790682, 0.1853059, 0.3546418, 
    0.3973827, 0.3012891, 0.2442091, 0.2796421, 0.1881056, 0.1529168, 
    0.1225131, 0.009362102, -0.01659834, 0.02134107, 0.1260288, 0.4379585, 
    0.5137399, 0.2957877, 0.1809444, 0.08030844, -0.1022253, -0.2499967, 
    0.2311392, 0.5776887, 0.7586129, 0.7054553, 1.204707, 1.113138,
  0.9061391, 0.8655468, 0.6832552, 0.4340689, 0.1203807, -0.1908496, 
    -0.4576956, -0.5129364, -0.4553192, -0.2286589, -0.04101253, 0.1322135, 
    0.158483, 0.0198274, -0.01148769, -0.1672169, -0.2341602, -0.1937468, 
    -0.079017, 0.01898104, 0.1327669, 0.1763704, 0.1602734, 0.1173859, 
    0.09054589, 0.118932, 0.1932162, 0.2247428, 0.1658398, 0.02236646, 
    -0.1330697, -0.3044239, -0.4322397, -0.4843391, -0.5351366, -0.6699837, 
    -0.5902638, -0.6250619, -0.786276, -0.8405241, -0.7813444, -0.7103646, 
    -0.6710417, -0.6862924, -0.7124643, -0.7314747, -0.7025033, -0.6378874, 
    -0.5427704, -0.4133759, -0.2683566, -0.1556776, -0.0644176, 0.01675129, 
    0.0995965, 0.1804882, 0.2412956, 0.2549837, 0.2545606, 0.2320996, 
    0.2065136, 0.2398469, 0.2544954, 0.3022981, 0.2626334, 0.1858919, 
    0.07371737, -0.03725266, -0.09278655, 0.03904933, 0.02230138, 0.08419916, 
    0.1598664, 0.1452506, 0.09202796, 0.02160144, 0.03882158, 0.1599483, 
    0.07259452, -0.009339213, 0.005244065, -0.03375316, 0.05179286, 0.158612, 
    0.2346709, 0.2361362, 0.2321483, 0.2135451, 0.1831076, 0.1464386, 
    0.3422065, 0.408711, 0.5177116, 0.5496287, 0.7090192, 0.4674666,
  0.2133486, 0.2860701, 0.4375846, 0.5110875, 0.3841341, 0.3219596, 
    0.1375356, -0.02761728, -0.09895509, -0.1279426, -0.1188931, -0.1051563, 
    -0.1060678, -0.1161588, -0.1219532, -0.1659962, -0.1566049, -0.1118783, 
    -0.05042, 0.03638013, 0.09748039, 0.08734043, 0.06393546, 0.06206363, 
    0.0646354, 0.007360101, 0.04163742, 0.05005193, 0.05867827, 0.0270865, 
    -0.06086922, -0.1741179, -0.331019, -0.4420542, -0.5427215, -0.6213673, 
    -0.6938608, -0.7572722, -0.7960581, -0.8157846, -0.7762501, -0.7309211, 
    -0.6789355, -0.6300262, -0.578366, -0.5269337, -0.4582325, -0.3748504, 
    -0.2953092, -0.2265104, -0.1661751, -0.1382779, -0.1237109, -0.08328128, 
    -0.05990887, -0.03614581, -0.01322913, 0.01920915, 0.06754887, 
    0.07840478, 0.08149737, 0.09044921, 0.1212108, 0.1465364, 0.1916373, 
    0.2096386, 0.1654654, 0.120039, 0.06981105, 0.04113269, 0.04640615, 
    0.04036772, 0.03755212, -0.01506841, 0.02039701, -0.06337565, 
    -0.06807959, -0.08324873, -0.05123381, -0.05955085, -0.08643901, 
    -0.1621387, -0.2455378, -0.2762668, -0.2105925, -0.07836592, 0.04756176, 
    0.1662794, 0.3309271, 0.4590354, 0.4655132, 0.5744653, 0.4926949, 
    0.4191594, 0.3289409, 0.2696149,
  0.2106967, 0.1622753, 0.1845411, 0.2204134, 0.108483, 0.1286978, 0.1280793, 
    0.1088898, 0.06295887, 0.02614245, 0.01878566, 0.008352757, 0.01829743, 
    0.01806957, 0.01548168, 0.01330072, 0.01870435, 0.02959302, 0.03154615, 
    0.02020174, 0.01352857, -0.006067783, -0.03219084, -0.05377286, 
    -0.05694669, -0.1178191, -0.1363737, -0.1395314, -0.1476857, -0.1683562, 
    -0.195814, -0.1884084, -0.2037728, -0.2389941, -0.2817676, -0.3257944, 
    -0.3760873, -0.4348276, -0.4943165, -0.5506316, -0.6074838, -0.6374968, 
    -0.6327768, -0.6116017, -0.5854949, -0.5540658, -0.5137013, -0.453724, 
    -0.4043588, -0.3501759, -0.2909474, -0.2374806, -0.1767058, -0.1181446, 
    -0.04280284, 0.03996083, 0.1143911, 0.163431, 0.2064323, 0.2376496, 
    0.2618684, 0.273229, 0.2847526, 0.2932649, 0.2877474, 0.2812533, 
    0.2815788, 0.2525747, 0.2145376, 0.1741079, 0.09964508, 0.08006504, 
    0.05420239, 0.002688721, -0.0026986, -0.03249997, -0.05779314, 
    -0.04244459, -0.06790042, -0.08679724, -0.1013482, -0.1205213, 
    -0.1301892, -0.1046515, -0.04838526, 0.03393865, 0.124401, 0.1858269, 
    0.2484572, 0.2726753, 0.2777207, 0.2907255, 0.3153183, 0.3323922, 
    0.3082712, 0.2645216,
  0.5816766, 0.5842155, 0.5672071, 0.5379916, 0.5128125, 0.4655958, 
    0.4038282, 0.3626333, 0.3043489, 0.2466503, 0.1812044, 0.1210644, 
    0.0744009, 0.04702467, 0.03970043, 0.05268872, 0.07319654, 0.07313143, 
    0.06806958, 0.05604159, 0.0389843, 0.01730461, -0.01498705, -0.05719082, 
    -0.1074838, -0.1556283, -0.1905567, -0.2693653, -0.3165496, -0.3650033, 
    -0.3977833, -0.4202929, -0.4296679, -0.4285449, -0.4273568, -0.4354298, 
    -0.4466277, -0.4549936, -0.4586718, -0.4751432, -0.4787728, -0.4757943, 
    -0.4729949, -0.4748667, -0.4713184, -0.4549122, -0.4414519, -0.4255176, 
    -0.4012663, -0.3682911, -0.3303517, -0.2828093, -0.2216602, -0.1589812, 
    -0.08756194, -0.02291349, 0.04619458, 0.1140982, 0.169453, 0.219632, 
    0.2720409, 0.3157258, 0.3459178, 0.3666862, 0.3829622, 0.3782746, 
    0.3603709, 0.3341503, 0.3088899, 0.2801952, 0.2432486, 0.1985383, 
    0.1646679, 0.1353385, 0.0589388, 0.03792644, 0.03437805, -0.02076519, 
    -0.045228, -0.06280613, -0.04988301, -0.04086578, -0.02966797, 
    -0.01897466, -0.002796292, 0.0222688, 0.0492382, 0.08818674, 0.1313509, 
    0.1906284, 0.2661328, 0.3290561, 0.3865918, 0.4578646, 0.5146518, 
    0.5567089,
  0.5252961, 0.5275911, 0.5311393, 0.5276563, 0.5125682, 0.5031608, 
    0.4801139, 0.4554558, 0.4307976, 0.3954785, 0.3620149, 0.3329784, 
    0.2963573, 0.2695506, 0.2400097, 0.2049837, 0.1753287, 0.1397004, 
    0.1107128, 0.08537102, 0.06839511, 0.05184236, 0.03958648, 0.01823232, 
    0.0003123879, -0.01817709, -0.03674805, -0.06119472, -0.08718765, 
    -0.1213022, -0.1517059, -0.1756642, -0.1950327, -0.2187955, -0.2450488, 
    -0.2753385, -0.2984668, -0.3188118, -0.342575, -0.3539844, -0.3639616, 
    -0.370944, -0.3825001, -0.3869109, -0.3841603, -0.389336, -0.3881642, 
    -0.3775683, -0.360853, -0.3454721, -0.3277475, -0.3052214, -0.2757943, 
    -0.2430795, -0.2041635, -0.1649382, -0.1179819, -0.07636401, -0.04218432, 
    0.001744717, 0.05034497, 0.1007845, 0.1408723, 0.1669954, 0.1939159, 
    0.2120963, 0.2329622, 0.2512076, 0.2659049, 0.2744335, 0.2665722, 
    0.2523795, 0.2450878, 0.2363801, 0.2273795, 0.2059602, 0.1889192, 
    0.1779003, 0.1682324, 0.1616406, 0.1589876, 0.1581087, 0.1609895, 
    0.1720735, 0.18861, 0.2083527, 0.232539, 0.2602245, 0.2898144, 0.3212759, 
    0.3509471, 0.3859243, 0.4185741, 0.4525261, 0.483011, 0.5100455,
  -0.4349256, -0.4031706, -0.3701134, -0.3375111, -0.3066363, -0.2784629, 
    -0.2539182, -0.2333455, -0.217021, -0.2062135, -0.1990185, -0.194447, 
    -0.1914849, -0.1891246, -0.1879852, -0.1868622, -0.1854298, -0.1834271, 
    -0.1805954, -0.1776005, -0.1745569, -0.171204, -0.1675906, -0.1636843, 
    -0.1582969, -0.1507286, -0.1400355, -0.124736, -0.1047487, -0.07888627, 
    -0.0471642, -0.010674, 0.0301137, 0.07449961, 0.122108, 0.1721883, 
    0.2238655, 0.2750864, 0.3244681, 0.3704157, 0.4139051, 0.4540901, 
    0.4901905, 0.5217986, 0.5484753, 0.5692921, 0.5870495, 0.5833869, 
    0.5785856, 0.5680552, 0.5578504, 0.5129762, 0.5039105, 0.5306191, 
    0.4682488, 0.4806833, 0.495739, 0.4679067, 0.3909535, 0.3152215, 
    0.3105824, 0.3203647, 0.2796743, 0.2560582, 0.2282422, 0.2008982, 
    0.1760285, 0.1566925, 0.1389842, 0.09375286, 0.05674124, 0.01532078, 
    -0.03000784, -0.0401969, -0.1125946, -0.176362, -0.2161746, -0.2378368, 
    -0.3375926, -0.3747191, -0.4153781, -0.4529252, -0.4882944, -0.5166149, 
    -0.537431, -0.5549443, -0.5672164, -0.5741986, -0.5765098, -0.574101, 
    -0.5668746, -0.5547326, -0.5374961, -0.5172331, -0.4930634, -0.4650359,
  -0.259614, -0.1886506, -0.1152139, -0.04657793, 0.009623528, 0.04318428, 
    0.05234909, 0.03691721, -0.001087666, -0.05069685, -0.1024873, -0.148581, 
    -0.177845, -0.1890104, -0.1846321, -0.1699507, -0.1488082, -0.1228155, 
    -0.09467423, -0.06210554, -0.03427351, -0.01542583, -0.009045638, 
    -0.01208931, -0.01754177, -0.01907194, -0.01313114, 0.003731012, 
    0.03519249, 0.0802927, 0.1363964, 0.1986213, 0.2629437, 0.3235564, 
    0.3777719, 0.4233937, 0.4589901, 0.4831104, 0.4948444, 0.4981165, 
    0.5068245, 0.4978247, 0.4118547, 0.3785858, 0.366786, 0.2936573, 0.36869, 
    0.3576059, 0.3454466, 0.3218617, 0.3837759, 0.2895374, 0.2983756, 
    0.2978065, 0.2685423, 0.3562696, 0.3505735, 0.3279824, 0.3334184, 
    0.3310584, 0.3266799, 0.3151894, 0.2918005, 0.262357, 0.2298541, 
    0.1883335, 0.1509473, 0.1142129, 0.08566466, 0.06717503, 0.06131542, 
    0.04964566, 0.01520491, -0.04050589, -0.08826065, -0.1522737, -0.2137971, 
    -0.2553496, -0.3062615, -0.3363233, -0.3547173, -0.3953583, -0.3396943, 
    -0.3781703, -0.3546346, -0.3387657, -0.327405, -0.3299444, -0.3399863, 
    -0.3542774, -0.3714161, -0.3830843, -0.3870077, -0.3770456, -0.351541, 
    -0.3131785,
  -0.206799, -0.1682086, -0.1208301, -0.08909202, -0.0842905, -0.08235312, 
    -0.074736, -0.06842077, -0.06905539, -0.08311796, -0.11567, -0.1746061, 
    -0.2329879, -0.2669072, -0.260983, -0.2116828, -0.1442027, -0.07818651, 
    -0.02183867, 0.01942098, 0.04622775, 0.06668679, 0.08055398, 0.09468158, 
    0.1045449, 0.1034055, 0.07803094, 0.04285836, 0.02925181, 0.03406882, 
    0.04949856, 0.06497717, 0.0756216, 0.08169222, 0.08756828, 0.09290886, 
    0.09305334, 0.08895397, 0.08205271, 0.07832527, 0.07979012, 0.0951376, 
    0.04175282, 0.0336132, -0.01988626, -0.06604505, -0.03139257, 0.04987359, 
    0.1399777, 0.2245315, 0.2980014, 0.368721, 0.4411659, 0.5048053, 
    0.5417682, 0.5439, 0.5311234, 0.5340688, 0.4957075, 0.4207234, 0.3067913, 
    0.1911011, 0.0942421, 0.04012489, 0.007392406, -0.01716733, -0.04721296, 
    -0.07584251, -0.09527647, -0.08256459, -0.05069685, -0.02670527, 
    -0.01913548, -0.01737785, -0.03811359, -0.05354309, -0.115962, -0.177485, 
    -0.1690717, -0.1560354, -0.118633, -0.05315375, 0.01676786, 0.04295629, 
    0.04269589, 0.04798561, 0.03590876, 0.05280304, 0.07900763, 0.0970571, 
    0.07016945, 0.001794338, -0.0892539, -0.1731253, -0.220439, -0.2332153,
  -0.05829728, 0.0103066, 0.0489133, 0.04219136, -0.01291933, -0.09355092, 
    -0.1428349, -0.1597781, -0.1854136, -0.1920214, -0.1361127, -0.003430367, 
    0.1627331, 0.2898965, 0.3344278, 0.3670287, 0.3326201, 0.255244, 0.12043, 
    -0.0454877, -0.08736622, 0.04056287, 0.1847525, 0.263171, 0.2881383, 
    0.3423053, 0.3978879, 0.4063185, 0.3479693, 0.2660358, 0.1680703, 
    0.07412505, 0.01719117, -0.03022099, -0.06789994, -0.07076454, 
    -0.02935815, 0.03393936, 0.1228061, 0.2289255, 0.3199587, 0.3742881, 
    0.3723021, 0.3509488, 0.2473183, 0.1491895, 0.01683235, 0.03418279, 
    0.1461461, 0.2646523, 0.402917, 0.525622, 0.6352251, 0.7087929, 
    0.6987994, 0.6522988, 0.6065303, 0.4106483, 0.2910357, 0.1524777, 
    0.08227873, 0.003926039, -0.06718364, -0.2004844, -0.292135, -0.3139124, 
    -0.3110642, -0.2603326, -0.1570587, -0.06550694, 0.03825283, 0.1123247, 
    0.1401734, 0.1762252, 0.1247916, 0.02184558, -0.0930953, -0.14679, 
    -0.1632285, -0.2108197, -0.09405541, 0.01606822, 0.08153033, 0.1230993, 
    0.1839718, 0.2259479, 0.2356972, 0.2067096, 0.2182492, 0.1801467, 
    0.21348, 0.2250037, 0.1229527, 0.0391314, -0.06718373, -0.09477186,
  0.05944324, 0.1570344, 0.3373413, 0.358469, 0.2622933, 0.07620955, 
    -0.2054963, -0.4574652, -0.5601683, -0.6840286, -0.5602975, -0.3816853, 
    -0.1998825, -0.06397724, -0.0199182, -0.1366, -0.3722768, -0.4442821, 
    -0.430481, -0.2291632, -0.1215294, 0.05264044, 0.325671, 0.5568233, 
    0.7409706, 0.9496291, 1.012927, 0.852056, 0.5676146, 0.3139687, 
    0.1546907, 0.08286428, -0.004375219, -0.1241832, -0.2311974, -0.2750444, 
    -0.2509241, -0.2069283, -0.1744576, -0.1125112, -0.0250926, 0.02642107, 
    0.04251814, 0.03366375, -0.00369072, -0.05040264, -0.1162071, -0.1312146, 
    -0.02556634, 0.1151893, 0.2689489, 0.3966997, 0.4534055, 0.4122597, 
    0.3337929, 0.1875852, 0.08006569, 0.03426492, -0.000940159, -0.05974551, 
    -0.1538536, -0.2362592, -0.3391238, -0.4547977, -0.5227665, -0.52026, 
    -0.4152634, -0.2608852, -0.1696091, -0.02239227, 0.1170118, 0.2206739, 
    0.1565139, -0.03209281, -0.2012172, -0.3095992, -0.4806928, -0.4876589, 
    -0.490068, -0.4491012, -0.2719365, -0.1568323, -0.04023075, 0.05382824, 
    0.1047561, 0.1525754, 0.2131549, 0.2455117, 0.2827513, 0.3701373, 
    0.4903684, 0.2362506, 0.1574583, 0.07056046, -0.01900685, -0.02429628,
  0.2584021, 0.169958, 0.3704789, 0.5141478, 0.4918654, 0.5039907, 0.4439178, 
    0.5960164, 0.4369507, 0.3085985, 0.1052933, -0.1125453, -0.2497522, 
    -0.3429164, -0.413327, -0.3505316, -0.3382435, -0.06102943, 0.2441778, 
    0.4830608, 0.4256544, 0.3877151, 0.3036494, 0.2767286, 0.3556833, 
    0.4586639, 0.4780331, 0.363287, 0.195529, 0.03493357, -0.07706261, 
    -0.1493931, -0.2775683, -0.4567981, -0.5919867, -0.6232371, -0.4785757, 
    -0.2326446, 0.01333523, 0.1544161, 0.2473683, 0.1820688, 0.1774955, 
    0.1176648, 0.05474043, -0.06550694, -0.07857656, -0.02686882, 
    -0.04622078, 0.1100786, 0.3698766, 0.5624061, 0.6055539, 0.5075233, 
    0.3570024, 0.174011, 0.08571351, 0.03055388, -0.0131799, -0.1429324, 
    -0.3941857, -0.6320925, -0.8624311, -1.00802, -1.113082, -1.126282, 
    -0.9618451, -0.6631798, -0.3949018, -0.1816695, -0.1765751, -0.245553, 
    -0.4460737, -0.6236615, -0.8007123, -0.8607709, -0.8353152, -0.5978965, 
    -0.4998008, -0.331588, -0.09596002, 0.008874059, 0.07847065, 0.1114132, 
    0.1370317, 0.1855018, 0.2230995, 0.2850624, 0.3611855, 0.50933, 
    0.6492714, 0.7040564, 0.6945347, 0.5510129, 0.3708533, 0.2631385,
  -0.2029421, -0.3279096, -0.3643028, -0.4163051, -0.4786422, -0.5242478, 
    -0.5380824, -0.5078902, -0.4465294, -0.3873334, -0.3858688, -0.411552, 
    -0.4694948, -0.5147585, -0.5465621, -0.5740523, -0.4891243, -0.2581186, 
    0.029284, 0.2260609, 0.3274446, 0.2089224, -0.03080678, -0.1642702, 
    -0.1887493, -0.1996057, -0.09244418, 0.03432941, 0.02290368, -0.02725887, 
    -0.0770632, -0.1676883, -0.2287724, -0.4330528, -0.7746553, -0.6790009, 
    -0.2448864, -0.2855926, -0.2094531, -0.1428027, -0.119153, -0.2383268, 
    -0.4264941, -0.5782356, -0.6169395, -0.6622036, -0.6087041, -0.4347618, 
    -0.1671023, 0.1164751, 0.2914587, 0.3234086, 0.2562701, 0.1455114, 
    0.04977572, 0.01191759, 0.0122596, -0.01195908, -0.1894821, -0.4739221, 
    -0.7898404, -1.083313, -1.267786, -1.379814, -1.467835, -1.481832, 
    -1.361634, -1.146481, -0.9282677, -0.8593712, -0.9408978, -1.057353, 
    -1.172278, -1.230612, -1.230416, -1.183069, -1.05444, -0.837838, 
    -0.5884727, -0.2962364, -0.1948041, -0.2447716, -0.2650189, -0.2833457, 
    -0.1573368, -0.08450142, -0.05696249, -0.01671165, 0.08672261, 0.2672076, 
    0.4742714, 0.5951698, 0.6220903, 0.5170936, 0.2411659, -0.0422813,
  -1.029049, -1.152063, -1.248336, -1.397034, -1.564043, -1.715182, -1.81829, 
    -1.823157, -1.773401, -1.676315, -1.52747, -1.301119, -1.082744, 
    -1.025224, -1.216224, -1.471741, -1.607125, -1.582565, -1.489498, 
    -1.412659, -1.367884, -1.26165, -1.078333, -0.8888471, -0.7214643, 
    -0.5521934, -0.3650352, -0.2038373, -0.05452091, 0.04648822, 0.08087939, 
    0.08789444, -0.03874946, -0.3025515, -0.627877, -0.9413047, -1.122229, 
    -1.15343, -1.131962, -1.199768, -1.33372, -1.379863, -1.312854, 
    -1.142151, -0.9390099, -0.7883101, -0.6409789, -0.4611942, -0.2560514, 
    -0.1302372, -0.1782191, -0.3361782, -0.4400682, -0.4336712, -0.3721478, 
    -0.2727664, -0.2172487, -0.2255173, -0.3099897, -0.5063928, -0.763001, 
    -0.9214319, -1.0304, -1.114401, -1.206067, -1.246302, -1.178984, 
    -1.089303, -1.101152, -1.190214, -1.267802, -1.250078, -1.166386, 
    -1.090198, -1.042444, -1.010169, -0.9648399, -0.8063276, -0.5987266, 
    -0.4753706, -0.5190392, -0.7101036, -0.8489871, -0.8650678, -0.8478477, 
    -0.8184695, -0.7519819, -0.6481895, -0.4826296, -0.2964317, -0.1851687, 
    -0.1885541, -0.2773074, -0.4427045, -0.6356081, -0.8321902,
  -0.6192183, -0.60553, -0.6583946, -0.7662721, -0.9423957, -1.093779, 
    -1.166566, -1.101673, -0.9630339, -0.891484, -0.8864551, -0.8951952, 
    -0.8686652, -0.9097459, -1.012431, -1.060478, -0.9829715, -0.88538, 
    -0.8788049, -0.9794068, -1.066842, -1.008085, -0.7943324, -0.5659956, 
    -0.4328901, -0.3184371, -0.1305791, 0.1169958, 0.3160844, 0.4283402, 
    0.3898149, 0.2545774, 0.03991246, -0.2057745, -0.5015264, -0.8300745, 
    -0.9918587, -0.9505012, -0.8784311, -1.007793, -1.251673, -1.369056, 
    -1.339369, -1.260348, -1.232419, -1.196237, -1.11515, -1.001412, 
    -0.8614056, -0.7589967, -0.7761843, -0.8932416, -0.9128544, -0.735673, 
    -0.4929974, -0.3624473, -0.3633749, -0.4340944, -0.5688275, -0.7217573, 
    -0.9151164, -1.004553, -0.9777957, -1.01458, -1.152144, -1.209127, 
    -1.109697, -1.010234, -1.11707, -1.36847, -1.531783, -1.511031, 
    -1.344755, -1.158232, -1.067444, -1.030188, -0.9561322, -0.8057415, 
    -0.6381309, -0.5292606, -0.5261033, -0.6038374, -0.6999475, -0.7350713, 
    -0.7153609, -0.6450646, -0.5351362, -0.3867639, -0.2778284, -0.2067019, 
    -0.1869102, -0.2753379, -0.4218876, -0.5618453, -0.6385056, -0.6271286,
  -0.4877403, -0.6131477, -0.6716604, -0.714678, -0.7308729, -0.7261524, 
    -0.6837373, -0.5882621, -0.4937954, -0.4846487, -0.5623341, -0.6837537, 
    -0.8641896, -1.088441, -1.186732, -1.086878, -0.9449019, -0.8493941, 
    -0.7961876, -0.733232, -0.6461387, -0.5574832, -0.4970825, -0.4715779, 
    -0.4035282, -0.241338, -0.00624609, 0.2403359, 0.372318, 0.3609898, 
    0.212878, -0.02208376, -0.2830858, -0.5551562, -0.8325, -1.05369, 
    -1.134729, -1.08486, -1.117787, -1.336911, -1.559535, -1.618275, 
    -1.56419, -1.523515, -1.451657, -1.290442, -1.081963, -0.9445932, 
    -0.8938282, -0.8844039, -0.8877566, -0.8234012, -0.6319461, -0.3816206, 
    -0.2226524, -0.1628869, -0.185185, -0.3042443, -0.4879028, -0.6809044, 
    -0.8614056, -0.9846647, -1.012936, -0.9604784, -0.9283003, -0.8911908, 
    -0.8254683, -0.7935184, -0.9487916, -1.235478, -1.459501, -1.491647, 
    -1.340199, -1.09098, -0.8683884, -0.7247527, -0.5762012, -0.4360807, 
    -0.3701789, -0.3386192, -0.3077111, -0.3053672, -0.4261029, -0.578512, 
    -0.5947715, -0.468372, -0.302861, -0.1714644, -0.1244105, -0.1138799, 
    -0.09486949, -0.1234502, -0.2126266, -0.2947721, -0.3262825, -0.3657682,
  -0.2338021, -0.1362765, 0.01979494, 0.09617949, 0.08569765, 0.08527422, 
    0.09660244, 0.09311914, 0.01974678, -0.1372352, -0.3460579, -0.5312309, 
    -0.6533012, -0.6896453, -0.5804007, -0.4177699, -0.3539186, -0.3415978, 
    -0.2614546, -0.1449668, -0.04180932, 0.01977921, -0.0257287, -0.08044863, 
    0.008988142, 0.2437539, 0.4412959, 0.5072463, 0.4350941, 0.2702508, 
    0.08170891, -0.07751894, -0.2523227, -0.4742637, -0.6791139, -0.7663708, 
    -0.778903, -0.8302865, -0.9603972, -1.077275, -1.083233, -1.063831, 
    -1.055628, -0.9687467, -0.7891083, -0.6906381, -0.7270637, -0.7765756, 
    -0.7541142, -0.716207, -0.623271, -0.3565879, -0.01884389, 0.196162, 
    0.2016478, 0.167403, 0.1010942, -0.1390424, -0.4715624, -0.7390103, 
    -0.9184697, -1.003073, -0.9557419, -0.7280729, -0.5249968, -0.4959278, 
    -0.6263797, -0.7998986, -1.01222, -1.245879, -1.3193, -1.155237, 
    -0.8712528, -0.5109499, -0.2242641, -0.03824568, 0.03986311, 0.07986975, 
    0.0783565, -0.05925775, -0.1637006, -0.2454553, -0.3938601, -0.4842899, 
    -0.4044563, -0.2196741, -0.03393197, 0.1460322, 0.2536657, 0.2680374, 
    0.2036983, 0.06650758, -0.07626629, -0.1313438, -0.1494915, -0.2124479,
  0.3313344, 0.4245317, 0.446928, 0.338448, 0.2436566, 0.2776895, 0.2647991, 
    0.1977243, 0.08742166, -0.007727861, -0.06124377, -0.1639946, -0.2338016, 
    -0.2261357, -0.1897748, -0.2080202, -0.2372682, -0.1192994, 0.07624078, 
    0.1538284, 0.1615273, 0.1457392, 0.08105826, 0.02648497, 0.08740616, 
    0.1987178, 0.2594919, 0.2851431, 0.2979522, 0.275475, 0.2124543, 
    0.1144562, -0.01069021, -0.1108041, -0.1772757, -0.2139454, -0.2698374, 
    -0.4104137, -0.5630503, -0.5881481, -0.5054004, -0.4336395, -0.4871385, 
    -0.4650357, -0.279912, -0.2422166, -0.3950489, -0.4750124, -0.3484831, 
    -0.1272262, 0.1068234, 0.3423702, 0.4998083, 0.5498244, 0.5095085, 
    0.4669142, 0.2878778, -0.07387304, -0.4193814, -0.5635865, -0.6563601, 
    -0.6251755, -0.4387336, -0.2336388, -0.197685, -0.3648074, -0.647099, 
    -0.8614221, -0.9658979, -0.9695927, -0.7741172, -0.4422324, -0.1636355, 
    0.0649941, 0.3655474, 0.5520539, 0.5384471, 0.4523306, 0.3020382, 
    0.1290888, -0.00170517, -0.05629516, -0.1160281, -0.1563275, -0.05377269, 
    0.2013056, 0.4581579, 0.5472366, 0.4732132, 0.4119012, 0.3301305, 
    0.2310743, 0.253226, 0.3288774, 0.3199906, 0.2798052,
  0.5593128, 0.4471059, 0.3860545, 0.4090037, 0.5224314, 0.6504431, 
    0.6530796, 0.5714066, 0.3838251, 0.1795936, -0.01291943, -0.1761029, 
    -0.2214155, -0.1727505, -0.1681604, -0.1182258, -0.003056288, 0.1453487, 
    0.2364944, 0.1899613, 0.09936881, 0.02759123, -0.01404297, -0.005188465, 
    0.09547925, 0.2207396, 0.3520708, 0.498132, 0.630163, 0.6873891, 
    0.6672556, 0.6244986, 0.5643585, 0.5362659, 0.4972198, 0.4142447, 
    0.2557812, 0.08240867, 0.07339168, 0.1335976, 0.1005733, 0.04422557, 
    -0.05888319, -0.2151495, -0.203447, -0.1048793, -0.05875301, 0.04261422, 
    0.1212766, 0.2679888, 0.542354, 0.6572629, 0.6255732, 0.6260127, 
    0.5738481, 0.4476762, 0.2322626, -0.02081347, -0.2512822, -0.3650029, 
    -0.4011357, -0.3212039, -0.1540979, -0.06132436, -0.09250927, -0.2099411, 
    -0.4276984, -0.5889121, -0.5451295, -0.310364, -0.05914378, 0.09443688, 
    0.2087924, 0.431042, 0.7175816, 1.06431, 1.257165, 0.933337, 0.4801794, 
    0.2486528, 0.2329788, 0.2285354, 0.2289749, 0.2199582, 0.3375361, 
    0.5916377, 0.7890009, 0.757637, 0.6143101, 0.6331578, 0.6826695, 
    0.5905309, 0.6526237, 0.7388382, 0.6390498, 0.5910192,
  0.1731319, 0.2186561, 0.4314326, 0.5331581, 0.6584509, 0.6959674, 0.479968, 
    0.2398963, -0.04574847, -0.3835088, -0.5893846, -0.6817347, -0.541126, 
    -0.3214808, -0.183655, 0.04347718, 0.1172401, 0.04679734, 0.03035861, 
    -0.05077744, -0.1199344, -0.06775331, 0.08498108, 0.1935744, 0.3172725, 
    0.4709022, 0.609395, 0.8252641, 0.9969926, 0.9670776, 0.8743852, 
    0.7873082, 0.693607, 0.6155796, 0.5673701, 0.5401893, 0.5013219, 
    0.4664749, 0.4519731, 0.3704137, 0.1562539, -0.1386843, -0.2464643, 
    -0.2306277, -0.1320762, -0.008768946, 0.0615598, 0.2022173, 0.2978554, 
    0.3946653, 0.5927609, 0.6623411, 0.7009642, 0.7534706, 0.619828, 
    0.3176796, 0.1758339, 0.1501015, 0.009752989, -0.07559836, -0.01840436, 
    0.1103878, 0.2314978, 0.2435256, 0.1482133, 0.02158582, -0.1871876, 
    -0.3557259, -0.2026657, -0.01464498, 0.05281925, 0.1411657, 0.4546911, 
    1.004789, 1.443233, 1.994812, 2.207898, 1.137992, 0.2391315, 0.3298053, 
    0.7119992, 0.586869, 0.3275263, 0.1805539, 0.2839879, 0.4088576, 
    0.3497432, 0.3669958, 0.4568723, 0.5916543, 0.6820838, 0.5900916, 
    0.6020708, 0.571667, 0.3652867, 0.25155,
  0.4209348, 0.6407589, 0.8557819, 0.9490433, 1.09211, 1.038399, 0.7316933, 
    0.4627317, 0.02062559, -0.5233525, -0.5313438, -0.2940068, -0.01581651, 
    0.2256386, 0.4661171, 0.634623, 0.4471393, 0.2731321, 0.2520546, 
    0.1322141, -0.03621034, 0.005960878, 0.1798867, 0.2820514, 0.4671913, 
    0.7520058, 0.8758339, 1.013741, 1.105538, 1.057312, 0.9699257, 0.7810585, 
    0.6162636, 0.6299353, 0.7482297, 0.7135128, 0.5954628, 0.6233274, 
    0.5478066, 0.2679889, 0.129024, -0.1134402, -0.3305952, -0.2778119, 
    -0.1005332, 0.01663792, 0.01048553, 0.09212619, 0.2921425, 0.4660846, 
    0.5665566, 0.694063, 0.8565305, 0.824483, 0.4535032, 0.09642312, 
    0.05491921, 0.1055377, 0.07895892, 0.1668658, 0.2834023, 0.3542193, 
    0.4375038, 0.3311887, 0.06178769, -0.05369085, -0.1967084, -0.2231246, 
    0.04350948, 0.175134, 0.3812212, 0.7511919, 1.102234, 1.581107, 1.865254, 
    2.170918, 2.03415, 0.7924677, 0.1373736, 0.6851113, 0.9887246, 0.5266802, 
    0.1778519, -0.1625129, -0.2481408, -0.01150346, 0.04780602, 0.2204137, 
    0.5129433, 0.5891966, 0.5621295, 0.4369667, 0.3616901, 0.3189492, 
    0.2809444, 0.3292356,
  0.6259478, 0.7995639, 0.8932981, 1.113561, 1.063382, 0.7322628, 0.4068072, 
    0.3214068, -0.2055463, -0.6934859, -0.3528445, 0.04876661, 0.09516966, 
    0.2862506, 0.6311886, 0.7264848, 0.5597205, 0.4685745, 0.2460322, 
    -0.01643503, -0.04991496, 0.006351233, 0.2016964, 0.3254269, 0.4518266, 
    0.6422075, 0.7141963, 0.7940794, 0.8310909, 0.9519241, 0.9504595, 
    0.538985, 0.385095, 0.5023965, 0.6880084, 0.741817, 0.6375526, 0.7085648, 
    0.4455929, 0.0375852, -0.05751568, -0.2969855, -0.3157516, -0.06342387, 
    -0.00282836, 0.1176469, 0.2220576, 0.3229368, 0.4851435, 0.5532913, 
    0.6229692, 0.7479041, 0.6887082, 0.3288448, -0.00673449, -0.1772097, 
    -0.07507759, 0.1013059, 0.1915402, 0.3578977, 0.438513, 0.3989621, 
    0.3180051, 0.04824604, -0.1717572, -0.05263305, -0.00561142, 0.01312232, 
    0.237748, 0.4407102, 0.7094765, 0.95072, 1.20321, 1.590303, 1.694828, 
    1.886609, 1.392648, 0.2822953, 0.06523821, 0.6330279, 0.6589882, 
    0.1468623, -0.02717745, -0.21707, -0.42817, -0.1021612, 0.1434771, 
    0.3030312, 0.4649941, 0.4640338, 0.4148476, 0.3414101, 0.2260618, 
    0.168998, 0.3279824, 0.481677,
  0.7406614, 0.9217155, 0.9453979, 1.109266, 0.6824739, 0.3424355, 0.1146848, 
    -0.04903591, -0.2996055, -0.3192509, 0.05806065, 0.2239296, 0.113057, 
    0.5790566, 1.115124, 0.9627967, 0.5962274, 0.328112, -0.0804652, 
    -0.2161422, -0.04366505, -0.01555634, 0.02972364, 0.04442096, 0.1529498, 
    0.3700397, 0.4645703, 0.5591016, 0.6938996, 0.9006701, 0.6405306, 
    0.2305377, 0.3194049, 0.5190956, 0.4377968, 0.4011594, 0.4359245, 
    0.445235, 0.1603065, -0.110641, -0.02813745, -0.07221365, 0.1496124, 
    0.288089, 0.08014631, 0.1871123, 0.3191929, 0.2889357, 0.1881869, 
    0.06344795, 0.1227086, 0.1493363, -0.1618943, -0.4873825, -0.4909469, 
    -0.3898073, -0.2018191, -0.07525659, 0.02353901, 0.1468137, 0.1012408, 
    0.02843809, -0.1126589, -0.252226, -0.2239057, -0.1456016, -0.1189252, 
    0.07777077, 0.3682005, 0.5306354, 0.6589394, 0.7412471, 1.01379, 
    1.358125, 1.449954, 1.526501, 0.8503771, -0.06721622, -0.2364057, 
    0.008092761, 0.1543007, -0.03686166, 0.008190393, -0.03998637, 
    -0.3570114, -0.348987, -0.04622011, 0.1867063, 0.260746, 0.3418819, 
    0.2919145, 0.1317745, 0.1322628, 0.2196977, 0.4675329, 0.572872,
  0.7464221, 0.792923, 0.7182345, 0.5862517, 0.08589244, -0.03842413, 
    -0.07499623, -0.290198, -0.0782188, 0.3358762, 0.4680853, 0.4332571, 
    0.242305, 0.6378456, 0.8997432, 0.5625846, 0.1919961, -0.1272099, 
    -0.2921512, -0.185576, -0.05001235, -0.04831958, -0.05113554, 
    -0.06666303, 0.1101112, 0.4525261, 0.4962919, 0.3855824, 0.4479198, 
    0.4864125, 0.222595, 0.1202348, 0.1472206, 0.1691769, 0.06647491, 
    0.15378, 0.2551138, 0.2085643, -0.003837347, -0.190361, -0.0692029, 
    0.1681356, 0.2791872, -0.1689248, -0.3872366, -0.1484833, -0.2559702, 
    -0.3665173, -0.3347294, -0.3774865, -0.5526006, -0.6828414, -0.8519821, 
    -0.7851526, -0.4918092, -0.3107059, -0.08165312, -0.05432558, 
    -0.02397078, 0.01461971, -0.1434044, -0.06721622, -0.02747011, -0.055058, 
    0.0370481, 0.1173378, 0.2340045, 0.5183144, 0.6619667, 0.5340533, 
    0.5489457, 0.7407427, 1.037324, 1.203389, 1.241979, 1.11716, 0.3755403, 
    -0.006767005, -0.1772752, -0.2509893, -0.2155235, -0.1529584, 
    -0.03175071, 0.03652728, -0.1965619, -0.3279097, -0.09636658, 0.1470416, 
    0.1871293, 0.3016964, 0.3030635, 0.2007523, 0.3232456, 0.4878457, 
    0.6789262, 0.6790724,
  0.5149617, 0.3961468, 0.3151093, 0.3584337, 0.261218, 0.2241737, 0.198197, 
    0.138464, 0.2005404, 0.2504592, 0.3634968, 0.3570356, 0.03076553, 
    0.3262408, 0.683255, 0.344095, 0.1518104, 0.06418014, 0.07311583, 
    0.04160547, 0.02243233, 0.01131582, -0.04112577, -0.007857561, 0.2029815, 
    0.4225454, 0.4009147, 0.2475615, 0.1598337, 0.03367877, -0.04745746, 
    0.005977035, -0.1706831, -0.2254684, -0.1237919, -0.06824183, 
    -0.06215477, -0.1790328, -0.174736, -0.3494923, -0.3814263, -0.2155728, 
    -0.5056438, -0.8572712, -0.6298146, -0.6706188, -0.9258108, -0.8800094, 
    -0.8487271, -0.9563118, -1.169463, -1.145553, -1.014938, -0.6974082, 
    -0.2874799, -0.1943646, -0.02327091, 0.03719461, 0.07845438, 0.1108111, 
    0.1773964, 0.4273151, 0.4061236, 0.3423053, 0.394828, 0.5525266, 
    0.6781939, 0.6424191, 0.5591507, 0.5304402, 0.6378615, 0.7377639, 
    0.8625844, 0.7655957, 0.7452197, 0.5754604, 0.32253, 0.2467649, 
    -0.1658167, -0.2074507, -0.1857872, -0.1695111, -0.1348595, -0.06233339, 
    -0.0008099675, -0.05992508, -0.01287079, 0.2278193, 0.3390335, 0.3713902, 
    0.4242711, 0.5418332, 0.6846066, 0.729821, 0.7155631, 0.5875032,
  0.1498585, 0.001224995, 0.03800869, 0.3291543, 0.42183, 0.3201048, 
    0.2995318, 0.2218137, 0.1463414, 0.1157424, 0.2029493, 0.01124978, 
    -0.2819135, 0.003893375, 0.5609264, 0.444665, 0.213871, 0.07492208, 
    0.08922863, -0.1502566, -0.3100386, -0.2652144, -0.1316531, -0.01130795, 
    0.006660223, 0.06958342, -0.0002734661, -0.2926719, -0.6075809, 
    -0.6126919, -0.5678024, -0.6236781, -0.7597132, -0.5305954, -0.4538051, 
    -0.4602664, -0.5452275, -0.6876917, -0.6320276, -0.8921347, -0.7480917, 
    -0.9736123, -1.251055, -1.048775, -0.7338181, -1.105758, -1.34334, 
    -1.10986, -1.054033, -1.003691, -0.8490198, -0.6081342, -0.6167116, 
    -0.2606895, 0.2167031, 0.2422564, 0.3463092, 0.3956093, 0.4579954, 
    0.4783241, 0.547302, 0.6704953, 0.5708209, 0.6209022, 0.6684119, 
    0.694779, 0.6958368, 0.6246785, 0.5841672, 0.594974, 0.6288445, 0.531904, 
    0.5535517, 0.470057, 0.4960175, 0.4699111, 0.5012079, 0.1762571, 
    -0.3759404, -0.0928835, -0.02104115, -0.1171186, -0.1154909, 
    -0.005969465, -0.05600202, -0.1012006, 0.3658078, 0.5872433, 0.6131709, 
    0.7059609, 0.7125852, 0.7153351, 0.6349156, 0.558825, 0.4631217, 0.288805,
  -0.1758595, -0.1731892, -0.06150413, 0.1138709, -0.02025983, -0.170325, 
    -0.05543268, -0.1153286, 0.01598692, 0.07591498, -0.06342411, 
    -0.09177756, -0.08800101, 0.1704133, 0.6268258, 0.4947461, 0.05631864, 
    -0.3110315, -0.2800418, -0.5048954, -0.6764613, -0.4156866, -0.199508, 
    -0.30221, -0.4746382, -0.3154262, -0.2860316, -0.5637333, -0.7022912, 
    -0.5562786, -0.4224247, -0.3351038, -0.2876915, -0.5220176, -0.6512822, 
    -0.5491989, -0.6755823, -0.6452926, -0.6317836, -1.090996, -1.041159, 
    -1.415947, -1.307874, -0.8234175, -0.8665165, -1.127177, -1.387398, 
    -1.102584, -0.5313601, -0.119918, 0.1514036, 0.2759479, 0.07822649, 
    0.4015501, 0.6064655, 0.4384479, 0.4792844, 0.5767616, 0.5884966, 
    0.6080279, 0.5625523, 0.5689002, 0.5419143, 0.5432652, 0.5657592, 
    0.5905313, 0.5168333, 0.4870477, 0.4991243, 0.4666209, 0.4238148, 
    0.3361197, 0.3622284, 0.2947307, 0.2591834, 0.2152704, 0.006774545, 
    -0.03651989, -0.105351, 0.02062535, -0.01418895, -0.05896425, 
    -0.03399682, -0.05289352, -0.1306279, 0.1817257, 0.8299031, 0.8116413, 
    0.582149, 0.5926471, 0.4710162, 0.3558469, 0.2877636, 0.2097688, 
    0.09707332, -0.05364275,
  -0.3088186, -0.1885381, -0.09840131, 0.03657603, -0.15553, -0.5196249, 
    -0.4711715, -0.5456995, -0.2777146, -0.2519656, -0.2464483, 0.0294466, 
    0.1413119, 0.4761102, 0.7534218, 0.253145, -0.2069949, -0.4640587, 
    -0.3901981, -0.3850873, -0.3506961, -0.1691531, -0.1814905, -0.2516889, 
    -0.320683, -0.1416465, -0.01339135, -0.2078087, -0.2757123, -0.2375776, 
    -0.1249312, -0.1182253, -0.1992963, -0.2889447, -0.3264123, -0.4675417, 
    -0.7246382, -0.7699671, -0.504277, -0.6612432, -0.9465946, -1.032011, 
    -0.6334925, -0.2501752, -0.3756635, -0.5532188, -0.665198, -0.3998659, 
    0.07772194, 0.1627643, 0.2008828, 0.3889199, 0.3173216, 0.481791, 
    0.5253782, 0.4505572, 0.4690793, 0.5418496, 0.4470578, 0.3922237, 
    0.3609408, 0.3519564, 0.4046912, 0.4427609, 0.4533079, 0.4104369, 
    0.3546419, 0.3880239, 0.371048, 0.3070178, 0.2051787, 0.2147503, 
    0.2756214, 0.1809597, 0.07946277, 0.09180072, 0.01099014, -0.05575788, 
    0.0462929, -0.05826437, -0.02891868, -0.02839786, 0.006758422, 
    0.05143613, 0.2484413, 0.4888058, 0.6292356, 0.7613156, 0.6621457, 
    0.494258, 0.2960321, 0.04184937, -0.1408002, -0.2106569, -0.2367971, 
    -0.2699187,
  -0.3016567, -0.1599411, 0.03887105, 0.3027543, 0.2330604, -0.241793, 
    -0.3236127, -0.4370893, -0.2962691, -0.3798302, -0.3488569, 0.1417508, 
    0.5051959, 0.6113969, 0.5385129, 0.1889036, -0.05209577, -0.2124473, 
    -0.2157513, -0.004878998, 0.05835342, -0.02843037, -0.2010704, 
    -0.1966921, -0.2882448, -0.02445903, 0.3848509, 0.1469438, -0.1596153, 
    -0.2747359, 0.06505859, -0.04141903, -0.5478642, -0.559599, 0.033858, 
    0.2636594, 0.1332229, -0.0632937, -0.006229877, -0.06345645, -0.4968874, 
    -0.3098594, -0.2295861, -0.275045, -0.5368614, -0.7077436, -0.6050906, 
    -0.4264449, -0.2548628, -0.2510541, -0.2738405, -0.08085561, 0.04149151, 
    0.2380083, 0.3686397, 0.4518592, 0.4217161, 0.4529498, 0.4071002, 
    0.3940794, 0.4100624, 0.4266802, 0.393835, 0.4531612, 0.4598505, 
    0.4059933, 0.3860717, 0.3550494, 0.2126503, 0.1473501, 0.102119, 
    0.1300812, -0.03730154, -0.3009405, -0.3231897, -0.08004172, -0.05051699, 
    -0.09104437, -0.04760355, 0.011039, 0.07375056, 0.05003637, 0.04300515, 
    0.08076555, 0.2072467, 0.2572955, 0.3061236, 0.6120805, 0.3907589, 
    0.2588254, 0.209639, -0.09133768, -0.2555466, -0.2164353, -0.2507451, 
    -0.2494917,
  -0.1492639, 0.07982141, 0.2159707, 0.2186236, 0.1330603, 0.02614317, 
    0.04630918, 0.01675189, -0.1527468, -0.3577112, -0.1816206, 0.3602242, 
    0.700768, 0.5256549, 0.2170774, 0.04054749, -0.1550418, -0.2435346, 
    -0.1823855, -0.1664675, -0.2565717, -0.4795535, -0.6967409, -0.7315717, 
    -0.4741498, 0.1859087, 0.5966998, 0.008109316, -0.3058881, -0.505888, 
    -0.04535753, -0.116793, -0.1765912, -0.5950645, -0.2303673, -0.009761781, 
    -0.01272401, 0.05488652, 0.2089394, 0.1269894, -0.1608523, -0.06306589, 
    -0.1833135, -0.2311814, -0.3479294, -0.3819135, -0.272311, -0.2066531, 
    -0.1008749, 0.05791378, 0.1044471, 0.1090696, 0.1428099, 0.1991248, 
    0.2168005, 0.2664912, 0.3262892, 0.3221551, 0.310876, 0.3265986, 
    0.2593298, 0.245186, 0.184509, 0.2725787, 0.3109576, 0.4058795, 
    0.3512083, 0.2011594, 0.1359088, 0.05778372, 0.004805207, 0.03568095, 
    -0.1565067, -0.3293907, -0.2910606, -0.1366498, -0.05759707, -0.0240196, 
    -0.0119265, 0.02681029, 0.03991264, 0.07840556, 0.1076373, -0.01845348, 
    -0.006572008, 0.1070838, 0.2108595, 0.2967647, 0.0738157, 0.1004596, 
    0.07047909, -0.1242638, -0.1472294, -0.168372, -0.2461716, -0.1804323,
  0.1708372, 0.1689162, -0.04898703, -0.1213666, -0.03363872, -0.01215434, 
    0.02488992, 0.07545957, 0.0006386042, -0.3158002, -0.2554162, 0.374613, 
    0.5566933, 0.466345, 0.2540727, 0.04396546, 0.1140662, 0.170886, 
    0.2672727, 0.1042356, -0.126282, -0.4646122, -0.6334271, -0.5638796, 
    -0.2765912, 0.1151243, 0.4548216, -0.09429953, -0.8316695, -0.7824832, 
    -0.1439252, -0.004813865, -0.01925071, -0.1430951, -0.3017867, 
    -0.3752406, -0.4319626, 0.06922555, 0.1009315, -0.09986591, -0.10304, 
    0.01888371, 0.07482457, 0.2973666, 0.4808631, 0.6557817, 0.630326, 
    0.6838093, 0.7334347, 0.6466832, 0.6257524, 0.5237339, 0.3890173, 
    0.2644566, 0.1628616, 0.01889968, -0.136113, -0.29194, -0.357939, 
    -0.3415002, -0.3495405, -0.3375613, -0.3541141, -0.2305464, -0.1554812, 
    -0.04141868, -0.06552349, -0.09236269, -0.07331972, -0.1009076, 
    -0.122685, -0.05113547, -0.06313092, -0.1123334, -0.1442833, -0.03179954, 
    -0.0259077, 0.0274452, 0.05241272, 0.1103066, 0.08166051, -0.04665983, 
    -0.1088183, -0.01739407, 0.02392864, 0.09248352, 0.07513356, 0.1652706, 
    0.1130574, 0.1680374, 0.05509818, -0.1109011, -0.08440375, -0.01016891, 
    0.1229528, 0.1920285,
  0.2012728, 0.4035194, 0.1558794, 0.1339719, 0.2432328, 0.3533236, 
    0.2619179, 0.3127154, 0.5384639, 0.2359739, -0.2196577, 0.005097747, 
    0.272839, 0.4668818, 0.3534381, 0.07360375, 0.3202349, 0.3841993, 
    0.5126664, 0.5327675, 0.2911822, -0.2996547, -0.6771445, -0.8111943, 
    -0.7948692, -0.7811322, -0.002844453, 0.1576536, -0.5705854, -1.254554, 
    -0.8221157, -0.1494754, 0.1459674, -0.05191672, -0.4685184, -0.3440065, 
    -0.4019822, -0.2375126, -0.2275352, -0.2058229, -0.07314062, 0.06084347, 
    0.2168818, 0.3158076, 0.3457394, 0.4711292, 0.4972363, 0.5744171, 
    0.6705759, 0.7354848, 0.747822, 0.7416213, 0.7750037, 0.7036655, 
    0.5418491, 0.3238642, 0.02594781, -0.2810836, -0.4814088, -0.6114708, 
    -0.6875125, -0.7192183, -0.6987596, -0.623613, -0.4365523, -0.2577436, 
    -0.1904421, -0.1629682, -0.1950645, -0.06238222, -0.03822857, 
    -0.06238222, 0.1794634, 0.3645546, -0.07711196, 0.001192003, -0.02379173, 
    0.1614296, 0.1268105, -0.06077123, -0.02504563, 0.03753567, 0.2197137, 
    0.1419952, 0.1739776, 0.2251985, 0.2510121, 0.2972848, 0.2126501, 
    0.314034, 0.262406, -0.004000068, -0.2251589, -0.2537559, 0.0004594922, 
    0.03325582,
  -0.002974987, 0.08013082, -0.07099259, -0.2004356, -0.1771284, 0.2132686, 
    0.2727902, -0.0803347, 0.1036496, 0.5716183, 0.1550168, 0.09718752, 
    0.1937699, 0.09272814, 0.1114947, -0.03282511, 0.1233273, 0.3977902, 
    0.6619503, 0.7473179, 0.5282099, 0.09733415, -0.04696989, -0.466403, 
    -0.7149217, -1.208509, -0.5747036, 0.3803912, 0.3401244, -0.7643516, 
    -1.474964, -0.9862431, -0.3485315, -0.05330019, -0.3742802, -0.4810834, 
    -0.4144819, -0.2715621, -0.2387823, -0.2421184, -0.247571, -0.2401981, 
    -0.1171844, 0.0407095, 0.1289909, 0.1601434, 0.1863475, 0.1774282, 
    0.1816597, 0.2395878, 0.2737346, 0.3532104, 0.3923869, 0.4808474, 
    0.4360557, 0.3535199, 0.2333374, -0.05937099, -0.2914677, -0.3872852, 
    -0.4370413, -0.5698371, -0.5666637, -0.5543592, -0.4622691, -0.4219205, 
    -0.2373173, -0.1022263, -0.04146755, 0.08735722, -0.02421522, 
    -0.04099584, 0.002249599, 0.2659543, 0.02334368, -0.03971028, -0.1629355, 
    -0.1836388, -0.252878, -0.3268192, -0.1989708, -0.0008749962, 0.1004264, 
    0.1441438, 0.176517, 0.1484079, 0.2207713, 0.2527699, 0.2822294, 
    0.4645538, 0.6167841, 0.5429236, 0.3519242, 0.2585323, 0.3811232, 
    0.1478229,
  0.5890175, 0.3128293, -0.1522911, -0.6531374, -0.9470177, -0.8659956, 
    -0.7028934, -0.7339317, -1.012855, -0.635934, -0.4064415, -0.1592573, 
    0.03156281, -0.2007776, -0.221725, -0.07789329, 0.008239508, 0.248539, 
    0.6428092, 0.9529331, 0.6992714, 0.4618196, 0.5551624, -0.02991223, 
    -0.4730599, -1.015768, -0.932239, -0.1786746, -0.1212692, -0.5578086, 
    -1.210331, -1.399443, -1.124329, -0.6198205, -0.4190392, -0.4515264, 
    -0.4317183, -0.3144495, -0.2931113, -0.3250124, -0.338912, -0.3807905, 
    -0.3256798, -0.2805302, -0.197067, -0.1153777, -0.08953166, -0.0674448, 
    -0.04962254, -0.06243181, -0.05795622, 0.04922152, 0.1058135, 0.2520714, 
    0.2716513, 0.1658077, 0.1122766, -0.02970076, -0.245863, -0.3682261, 
    -0.3191681, -0.3569622, -0.3886027, -0.3700967, -0.2882609, -0.3061476, 
    -0.2698212, -0.3251922, -0.01264298, 0.3054889, 0.394356, 0.7737018, 
    0.4062862, -0.09065437, -0.2073851, -0.1942677, -0.3496382, -0.4630821, 
    -0.3964645, -0.2477664, -0.2156051, -0.102747, 0.004577398, 0.04282522, 
    0.08665681, 0.07658148, 0.1032596, 0.1745167, 0.2935424, 0.4611216, 
    0.878716, 1.092484, 0.9057981, 0.8478066, 1.021146, 0.9572303,
  0.4805536, 0.2978386, 0.06098998, -0.07712865, -0.3377243, -0.6016893, 
    -0.7693489, -0.4979622, -0.5619755, -0.6553679, -0.5817838, -0.2496057, 
    -0.07748637, -0.3001915, -0.1891725, -0.05452085, 0.05207092, 0.02702188, 
    0.547822, 0.9455924, 0.5846221, 0.8269242, 1.472888, 0.4802608, 
    -0.3963506, -0.2878218, -0.2307582, -0.3519819, -0.8516565, -1.356296, 
    -1.607907, -1.014205, -0.5798793, -0.8259565, -0.8684207, -0.5756962, 
    -0.5341109, -0.5432906, -0.4143846, -0.3333949, -0.384111, -0.4952599, 
    -0.4542443, -0.4087365, -0.4195275, -0.3373985, -0.2498171, -0.2105434, 
    -0.2151821, -0.1675751, -0.112448, 0.009752274, 0.1414907, 0.1947134, 
    0.2483265, 0.2216175, 0.111738, -0.01684284, -0.2261848, -0.4924939, 
    -0.6429658, -0.6549602, -0.6795697, -0.6757274, -0.5786419, -0.4086385, 
    -0.3349729, -0.5552053, -0.06536102, 0.2506386, 0.1918495, 0.1775591, 
    0.07904017, 0.1385127, -0.2418422, -0.3827437, -0.3809857, -0.4951296, 
    -0.636487, -0.5866335, -0.4760217, -0.3122849, -0.2004033, -0.1983523, 
    -0.1525025, -0.1369274, -0.1329069, -0.09955645, -0.04776478, 0.09266472, 
    0.2797413, 0.5101776, 0.2031455, 0.1452672, 0.3613312, 0.575557,
  0.1395543, 0.05932975, -0.1156703, -0.2237105, -0.3211064, -0.4119428, 
    -0.6297981, -0.7266238, -0.6994274, -0.597604, -0.5039024, -0.08505487, 
    -0.0988894, -0.561601, -0.2007611, 0.1039424, -0.2361128, -0.316972, 
    0.3160682, 0.5410193, 0.200362, 0.5599159, 1.454317, 0.9294472, 
    -0.361486, -0.5208299, -0.06304955, 0.1481807, -0.1906865, -0.8665655, 
    -1.547799, -0.9633102, -0.363017, -0.8117639, -1.048206, -0.7992474, 
    -0.6084435, -0.5508099, -0.5535117, -0.5261517, -0.4730268, -0.5038536, 
    -0.563603, -0.5300256, -0.5107062, -0.5351201, -0.5866663, -0.5722294, 
    -0.5019331, -0.3977175, -0.2414348, -0.05585551, 0.1487668, 0.2384968, 
    0.3204465, 0.211462, -0.01786733, -0.1674278, -0.3049114, -0.4257131, 
    -0.6071908, -0.7373178, -0.7976532, -0.7457151, -0.6924605, -0.4762321, 
    -0.1884389, -0.0801239, 0.05527729, 0.1111855, 0.04461646, -0.2486455, 
    -0.207711, 0.09987354, -0.2876264, -0.4206018, -0.3688764, -0.4704551, 
    -0.5804975, -0.5151329, -0.3617637, -0.3115522, -0.2421511, -0.1557256, 
    -0.1286426, -0.1574342, -0.1267219, -0.1023569, -0.1159778, -0.03646946, 
    -0.0162878, 0.2342014, 0.1683307, 0.07563853, 0.02236676, 0.02002335,
  -0.291435, 0.008678675, -0.1185509, -0.3117802, -0.3322554, -0.3314252, 
    -0.4392704, -0.5669235, -0.7285445, -0.7756639, -0.8144498, -0.3762008, 
    -0.3410606, -0.7033002, -0.1425907, 0.02775443, -0.5403932, -0.4728316, 
    -0.05347967, 0.1975299, 0.1237669, 0.2131548, 0.6721878, 1.357605, 
    1.12279, 0.09857106, -0.02576113, 0.2646351, 0.1205924, -0.3144331, 
    -0.8225226, -0.8049282, -0.4362103, -0.5097782, -0.6127241, -0.6524702, 
    -0.4929162, -0.4601361, -0.5568158, -0.5569786, -0.5289188, -0.4603477, 
    -0.4675255, -0.5359011, -0.571155, -0.5692996, -0.6498008, -0.719788, 
    -0.7269006, -0.6292281, -0.4048306, -0.1995571, -2.884865e-005, 
    0.05187559, 0.07978868, 0.07384777, -0.1180143, -0.3115196, -0.4382937, 
    -0.5594361, -0.6989224, -0.8241506, -0.9496551, -0.9583626, -0.9936323, 
    -0.7661896, -0.3301725, -0.009729505, 0.1542031, -0.01422143, 0.1247434, 
    0.3521197, 0.3841019, 0.3147823, -0.1277305, -0.2373659, -0.3166628, 
    -0.4714155, -0.6705202, -0.8106732, -0.7489871, -0.6012006, -0.4239382, 
    -0.3248008, -0.2573367, -0.2539187, -0.2655566, -0.2758424, -0.3054819, 
    -0.2578259, -0.3160105, -0.06391048, 0.2325573, 0.3576858, 0.05019927, 
    -0.3654747,
  -0.3336065, -0.3563116, -0.2357384, -0.3564415, -0.2788047, -0.2276492, 
    -0.2057416, -0.2577761, -0.6800581, -0.7333624, -0.5612429, -0.5693484, 
    -0.8158329, -0.8259729, -0.1928672, -0.2635053, -0.6664838, -0.7093225, 
    -0.2637331, 0.1347692, 0.08239245, 0.05319369, 0.08747128, 0.5663124, 
    0.9012728, 0.5779011, 0.1213093, 0.01328444, -0.008606195, 0.405212, 
    0.3517291, -0.1384241, -0.09376243, 0.1127317, 0.06504291, -0.06021756, 
    -0.002372444, -0.06412381, -0.2293583, -0.3263472, -0.4517053, 
    -0.4799443, -0.4563767, -0.4498498, -0.5425091, -0.6564742, -0.6863568, 
    -0.7501264, -0.8915163, -0.7949506, -0.5368452, -0.3166791, -0.01578391, 
    0.1498247, 0.1192418, 0.03527391, -0.2854129, -0.6228315, -0.7010542, 
    -0.6875938, -0.7125612, -0.8375618, -0.9386201, -0.995749, -1.027079, 
    -0.7037404, -0.4091599, -0.09480411, 0.0254758, -0.06457949, 0.2605993, 
    0.6764686, 0.6699095, 0.3181189, 0.08921278, -0.03513616, -0.2628216, 
    -0.5077761, -0.6469363, -0.742444, -0.7895143, -0.821871, -0.8240198, 
    -0.7527633, -0.5174929, -0.3747846, -0.3435671, -0.3179162, -0.3541471, 
    -0.2801719, -0.3234994, -0.470912, -0.09320784, 0.4262738, 0.5802445, 
    0.1515501,
  0.3701375, 0.2035357, 0.1035846, -0.1948041, -0.3711062, -0.4958946, 
    -0.3726037, -0.2046999, -0.482825, -0.5681115, -0.2597618, -0.2131472, 
    -0.5162885, -0.528349, -0.2948855, -0.4273725, -0.7748497, -1.146839, 
    -0.7102014, -0.01601207, 0.06300819, -0.2602503, -0.2109017, -0.1712203, 
    -0.1696901, -0.007842064, 0.160013, 0.1849158, 0.07729877, 0.4708369, 
    0.7482784, 0.421309, 0.2875527, 0.2834837, 0.3995479, 0.4210976, 
    0.3214068, 0.2418333, 0.2307652, 0.102917, -0.06549096, -0.2136357, 
    -0.389905, -0.3721478, -0.3702273, -0.5823042, -0.6898078, -0.714873, 
    -0.8402634, -0.844137, -0.6565228, -0.448043, -0.1650678, 0.1279498, 
    0.2034381, 0.08086322, -0.2023399, -0.5974408, -0.8927859, -0.9341108, 
    -0.8080367, -0.7763145, -0.8611786, -0.9081187, -0.6879365, -0.3855431, 
    -0.1248497, 0.1134153, 0.2738807, 0.4895872, 0.6506547, 0.6288449, 
    0.6171097, 0.4362013, 0.290287, 0.4246944, 0.3105831, -0.1777147, 
    -0.4824671, -0.5439579, -0.5466435, -0.6160609, -0.7184861, -0.7525682, 
    -0.7004032, -0.6626917, -0.528398, -0.4655235, -0.4940391, -0.4532351, 
    -0.3434371, -0.3382611, -0.5085244, -0.3751097, 0.02445054, 0.4996944,
  -0.07221293, -0.140312, -0.2948855, -0.4314579, -0.4292443, -0.436015, 
    -0.3339643, -0.1315391, -0.1587689, -0.4349409, -0.398043, -0.314726, 
    -0.3187464, -0.3561811, -0.2343386, -0.2785932, -0.4496544, -0.8614546, 
    -0.9893192, -0.5716596, -0.5137172, -0.7710094, -0.6705205, -0.09436488, 
    0.2514036, 0.1177771, 0.08442767, -0.08105084, -0.3954552, -0.1738731, 
    -0.05645812, -0.09547174, 0.02874708, 0.1259967, 0.1685746, 0.1961625, 
    0.07015359, 0.02171606, 0.2838255, 0.3675168, 0.2552605, 0.1117063, 
    -0.08596611, -0.2504847, -0.338115, -0.3364384, -0.3611133, -0.4327445, 
    -0.5694788, -0.7242315, -0.703805, -0.5191209, -0.3161263, -0.09753895, 
    0.09853876, -0.01890922, -0.2876428, -0.6351362, -0.9703901, -1.105384, 
    -0.9996544, -0.6926721, -0.5127244, -0.4814255, -0.2976201, -0.1685672, 
    -0.07546816, 0.1515989, 0.2505084, 0.4699414, 0.7219108, 0.7061234, 
    0.8399453, 0.7566609, 0.3540888, 0.4404659, 0.5517942, 0.3357297, 
    -0.08964479, -0.3554002, -0.286129, -0.1340783, -0.1410284, -0.2690237, 
    -0.4201629, -0.5201304, -0.476299, -0.3599248, -0.2541143, -0.2818647, 
    -0.4511517, -0.3998009, -0.3211064, -0.5090299, -0.4740196, -0.2010216,
  -0.1076459, -0.074736, -0.3270961, -0.476103, -0.3485638, -0.1005821, 
    0.1429237, 0.3051957, 0.2753456, 0.02609432, -0.08920512, 0.001745224, 
    -0.02465487, 0.1556842, 0.342468, 0.07200903, -0.1959597, -0.3830365, 
    -0.6208945, -0.3510866, -0.04171193, -0.336601, -0.5958784, -0.3637006, 
    0.1546751, 0.3526568, 0.46711, 0.08849669, -0.2745567, -0.2102989, 
    -0.29456, -0.3114383, -0.2024051, 0.002363861, 0.05306375, 0.06876981, 
    0.09865296, 0.09534892, 0.3104531, 0.6615924, 0.7747922, 0.6895052, 
    0.5648638, 0.313041, -0.02924418, -0.1545372, -0.1085737, -0.05979419, 
    0.007946014, -0.09929633, -0.3049116, -0.3879359, -0.2928185, -0.1314092, 
    -0.0650351, -0.1984501, -0.3812466, -0.5952114, -0.8091599, -1.000208, 
    -1.080042, -0.7665815, -0.1150841, 0.2506223, 0.1462604, -0.1152306, 
    0.05244526, 0.3830767, 0.06167376, 0.05382872, 0.7521197, 1.228405, 
    1.3231, 1.174695, 0.7941443, 0.5267616, 0.5617551, 0.6208697, 0.4669472, 
    0.1016639, -0.1534795, -0.1361129, 0.03524137, 0.2102089, 0.1622431, 
    -0.09143591, -0.1789846, -0.09587932, 0.04139376, -0.05513966, 
    -0.2185509, -0.3043419, -0.2526981, -0.1898238, -0.3549278, -0.3024701,
  0.3147172, 0.2620641, -0.1001917, -0.1376589, -0.02620071, 0.1485227, 
    0.3542193, 0.6321979, 0.766817, 0.5434772, 0.1848671, 0.2099485, 
    0.1391965, 0.132914, 0.4970742, 0.437162, 0.1508827, -0.1066043, 
    -0.2506635, 0.08546931, 0.6761432, 0.8147987, 0.4344928, 0.2080605, 
    0.1207232, 0.08520892, 0.1055703, -0.1328088, -0.278935, -0.1518679, 
    -0.0316205, -0.02253845, 0.07689178, 0.2639036, 0.3489622, 0.3343951, 
    0.3256549, 0.4025103, 0.5822955, 0.9882362, 1.116768, 1.026143, 
    0.9576858, 0.8724488, 0.6447954, 0.427315, 0.2967975, 0.2422075, 
    0.2714715, 0.3731158, 0.3537798, 0.10391, -0.2090783, -0.336585, 
    -0.4170537, -0.5404263, -0.6195765, -0.8040495, -0.9821744, -1.014857, 
    -0.9669722, -0.6171024, 0.1076208, 0.7762567, 0.7607297, 0.2094928, 
    0.306026, 0.5489134, 0.1253945, -0.258769, 0.2153359, 0.7960324, 
    1.082865, 1.248946, 1.001257, 0.8628945, 0.591817, 0.4595904, 0.3483111, 
    0.1115598, -0.1459597, -0.3190229, -0.161292, 0.2409866, 0.6395872, 
    0.6536171, 0.5691602, 0.679414, 0.705765, 0.421423, 0.07946324, 
    -0.109274, -0.1160282, 0.04056358, 0.0921424, 0.1490598,
  0.4428098, 0.5045773, 0.2119504, 0.04598366, 0.1072467, 0.115873, 
    0.06501037, 0.3587115, 0.8088906, 0.7177935, 0.2724973, 0.1019081, 
    0.2091347, 0.2384316, 0.30308, 0.3370318, 0.3378456, 0.2593625, 
    0.1311236, 0.2568398, 0.6407916, 0.7012084, 0.5064003, 0.2614132, 
    0.08102596, 0.05138731, 0.03971738, -0.06223577, -0.03897727, 0.1266314, 
    0.2964393, 0.3235061, 0.3553584, 0.5414751, 0.6468138, 0.503194, 
    0.3477252, 0.4568394, 0.6369665, 0.8780799, 1.22546, 1.356465, 1.336543, 
    1.389538, 1.333712, 1.158011, 1.117598, 1.137162, 0.9606324, 0.8399128, 
    0.9069211, 0.8261595, 0.3819537, -0.0901165, -0.37887, -0.5579228, 
    -0.8707647, -1.063115, -1.06279, -1.007207, -0.9363412, -0.6379035, 
    -0.0174768, 0.5969114, 0.8257524, 0.5101109, 0.3349322, 0.2685585, 
    0.120235, -0.0457319, 0.03953844, 0.1721555, 0.4100136, 0.5755898, 
    0.4775918, 0.3472044, 0.3191933, 0.2581744, 0.09886453, 0.04687884, 
    -0.1329877, -0.4419232, -0.5970341, -0.3399053, 0.2785683, 0.6415236, 
    0.7819538, 0.9878618, 1.189668, 1.078682, 0.625492, 0.1608595, 
    0.05635095, 0.2286983, 0.3270543, 0.2869505,
  0.5213737, 0.8661007, 0.6984739, 0.3842161, 0.2499387, 0.1637408, 
    0.05698621, 0.09790425, 0.2890012, 0.2752643, 0.03532286, -0.04675722, 
    0.2130247, 0.4577349, 0.4577186, 0.2827349, 0.2209348, 0.311983, 
    0.2163124, 0.1071816, 0.3560748, 0.7070676, 0.7038773, 0.4410032, 
    0.3888059, 0.4097207, 0.2878457, 0.1111041, 0.1227089, 0.1743202, 
    0.1892126, 0.2697628, 0.3220899, 0.3741573, 0.3714554, 0.3487667, 
    0.4196165, 0.4142455, 0.1464067, 0.194079, 0.8085486, 1.160225, 1.231514, 
    1.329057, 1.399304, 1.308532, 1.287129, 1.472042, 1.464538, 1.315238, 
    1.326697, 1.346553, 1.005391, 0.5142617, 0.1268103, -0.22734, -0.7056117, 
    -0.9598436, -0.9138312, -0.8018355, -0.7155564, -0.26318, 0.2081416, 
    0.4904494, 0.383044, 0.3027381, 0.1418495, -0.03090437, 0.08844784, 
    0.3534544, 0.2910032, 0.1113157, 0.2041705, 0.4182981, 0.5266151, 
    0.4663938, 0.3553749, 0.244063, 0.1655312, 0.1422076, -0.03295541, 
    -0.3725549, -0.6094363, -0.7431116, -0.4448694, -0.06277293, 0.2593788, 
    0.5956907, 0.823311, 0.9064652, 0.8275099, 0.5381055, 0.2602898, 
    0.1221715, 0.08649445, 0.1956251,
  0.1703, 0.2394081, 0.4903846, 0.708858, 0.8531126, 0.8593463, 0.7369179, 
    0.5267454, 0.416996, 0.341817, 0.1658567, 0.03415097, 0.1569374, 
    0.4043494, 0.5487668, 0.4216998, 0.232442, 0.1661496, 0.155619, 
    0.1320025, 0.2553098, 0.5453, 0.6446325, 0.4655309, 0.3486692, 0.2683469, 
    0.189636, 0.1675169, 0.1923541, 0.08903366, -0.02190375, 0.03605497, 
    0.2322139, 0.2698278, 0.04961324, 0.03948927, 0.2321488, 0.283793, 
    0.01798892, -0.4035776, 0.1146846, 0.4559606, 0.599727, 0.8307004, 
    1.067696, 1.097302, 1.093802, 1.311006, 1.580993, 1.683484, 1.698099, 
    1.605391, 1.280586, 0.8327832, 0.3840204, -0.1070765, -0.677861, 
    -0.8828743, -0.6339157, -0.2626266, -0.06837201, 0.1147172, 0.2279333, 
    0.05425179, -0.03350866, 0.01808649, 0.01860738, -0.06938092, 
    -0.04376243, 0.1259804, 0.1617877, 0.09445369, 0.1335649, 0.3096064, 
    0.5414424, 0.4531126, 0.4065631, 0.2460162, 0.2180539, 0.2644569, 
    0.1048702, -0.2514125, -0.7890753, -0.6875125, -0.664368, -0.5093874, 
    -0.1244754, 0.2948605, 0.4831418, 0.4874387, 0.3738808, 0.2193073, 
    0.1511592, 0.2350135, 0.2686725, 0.2378293,
  -0.3726851, -0.2909306, 0.07231832, 0.5159218, 0.8241249, 1.064913, 
    1.007279, 0.9826536, 0.6631712, 0.4821165, 0.3689165, 0.2976764, 
    0.3052936, 0.3772499, 0.4448442, 0.3822141, 0.2280312, 0.05775118, 
    -0.09452742, -0.170976, -0.1446739, 0.02412486, 0.2654006, 0.4106479, 
    0.4446322, 0.3512732, 0.2789426, 0.2520871, 0.2460487, 0.1575071, 
    0.023067, -0.0412885, 0.03504622, 0.113887, 0.03569698, -0.00618124, 
    0.1046585, 0.1304889, 0.01434255, -0.3046355, -0.3002083, -0.006587982, 
    0.2240593, 0.2936394, 0.3227413, 0.4938507, 0.6308134, 0.8421423, 
    1.206319, 1.560567, 1.794454, 1.706335, 1.446309, 1.007312, 0.5403359, 
    0.03644586, -0.4437463, -0.5981247, -0.3331833, 0.001533508, 0.3012079, 
    0.1183467, 0.05286813, -0.04428339, -0.03432232, 0.07554097, 0.2310423, 
    0.2556516, 0.2161822, 0.2415729, 0.2763547, 0.2816933, 0.1640825, 
    0.03709674, 0.04580426, 0.1874062, 0.2027383, 0.2104693, 0.277315, 
    0.4000361, 0.2010615, -0.1384242, -0.2896286, -0.1436487, 0.007018566, 
    0.003437877, 0.02331102, 0.1959022, 0.4118528, 0.5301145, 0.4264198, 
    0.1975949, 0.04775769, 0.05044323, 0.05931371, -0.1385217,
  -0.7916138, -0.5031213, 0.05960655, 0.2523152, 0.4522337, 0.6338418, 
    0.7556516, 0.7738158, 0.6456093, 0.5522988, 0.5367063, 0.4948769, 
    0.3706581, 0.2939817, 0.2539101, 0.26794, 0.2577024, 0.1515989, 
    -0.04612245, -0.1817833, -0.2575157, -0.247864, -0.1753054, -0.09849882, 
    -0.006815851, 0.06403375, 0.03765029, -0.01638615, -0.0341596, 
    -0.04164672, -0.08523379, -0.113196, -0.05317, 0.02303445, 0.029789, 
    0.02098364, 0.03839898, 0.03109086, 0.08130264, 0.1653354, 0.2010124, 
    0.1270864, 0.02158523, -0.02120376, -0.06903934, -0.0554657, -0.05455399, 
    -0.6090789, -0.5130992, -0.09537458, 0.420218, 0.8097203, 1.272725, 
    0.9553424, 0.4828652, 0.08320697, -0.1701622, -0.2808067, -0.1720504, 
    -0.1511358, -0.06910455, -0.03692675, -0.01850224, 0.02923554, 
    0.04547912, 0.07853574, 0.1406614, 0.2089719, 0.2768756, 0.3725787, 
    0.4439654, 0.4793331, 0.3176469, 0.1231644, -0.01988578, -0.09091449, 
    -0.17428, -0.1873171, -0.0503056, 0.08113933, 0.05736017, -0.2200645, 
    -0.3067833, -0.2615522, -0.1104457, 0.1400754, -0.01083684, -0.2800584, 
    -0.3646449, -0.2257611, -0.005969435, 0.1937538, 0.1822304, 0.004707634, 
    -0.2971804, -0.6831341,
  -0.7612592, -0.7719851, -0.6179488, -0.1695274, -0.001493573, 0.1407102, 
    0.2153359, 0.264164, 0.2864133, 0.3203163, 0.421358, 0.4712115, 
    0.4083534, 0.2908404, 0.2279498, 0.2156614, 0.1856484, 0.09001036, 
    -0.02559838, -0.1429975, -0.2083295, -0.1823692, -0.1533816, -0.1382123, 
    -0.1228151, -0.1138145, -0.1057904, -0.1273074, -0.1565717, -0.2345827, 
    -0.3512169, -0.4444623, -0.4547814, -0.3668256, -0.2255658, -0.1103965, 
    -0.06252871, -0.04672467, -0.04019797, -0.04067004, -0.01716769, 
    -0.05885029, -0.1442344, -0.2953579, -0.4119104, -0.4451624, -0.4733691, 
    -0.4724576, -0.3837032, -0.096416, 0.3504596, 0.7685251, 1.113708, 
    1.11208, 0.8237669, 0.4889199, 0.2254107, 0.09769265, 0.1207233, 
    0.1369179, 0.1679725, 0.2188027, 0.2485064, 0.2531288, 0.2167193, 
    0.1698443, 0.1363808, 0.2378619, 0.4706581, 0.6931028, 0.833858, 
    0.8201861, 0.6749386, 0.4985063, 0.339587, 0.2361202, 0.07912165, 
    -0.01703715, -0.04571557, -0.03031874, -0.03572226, -0.1798141, 
    -0.3193484, -0.3835086, -0.2637331, -0.09451151, -0.07789326, -0.4752903, 
    -0.5218711, -0.6349897, -0.7035449, -0.2629359, 0.05353522, 0.03118849, 
    -0.2113732, -0.5473269,
  0.003502965, -0.2061974, -0.4437299, -0.5779096, -0.6161583, -0.3196414, 
    -0.2398236, -0.1129519, 0.05220109, 0.2111041, 0.3833372, 0.5325885, 
    0.6148313, 0.587406, 0.5052285, 0.3757688, 0.2035357, -0.02616805, 
    -0.26956, -0.3962202, -0.3689415, -0.2861615, -0.1927534, -0.1515914, 
    -0.1334599, -0.1001917, -0.08282506, -0.03972602, -0.02522402, 
    -0.1015424, -0.2746543, -0.4682417, -0.6094037, -0.6392052, -0.5324831, 
    -0.4737267, -0.405107, -0.342851, -0.3083783, -0.2646446, -0.2487755, 
    -0.2568647, -0.2812299, -0.332646, -0.3898399, -0.4282351, -0.4765751, 
    -0.4929651, -0.5217903, -0.3667285, -0.1809378, 0.07029915, 0.3755894, 
    0.5190467, 0.5337605, 0.4384803, 0.3830278, 0.3195189, 0.3175005, 
    0.3161985, 0.3319536, 0.3333372, 0.3433795, 0.3199583, 0.2509967, 
    0.1926145, 0.1945677, 0.2796425, 0.4705279, 0.6330116, 0.7799844, 
    0.770235, 0.6256386, 0.4660518, 0.4445187, 0.3609085, 0.2730342, 
    0.150785, 0.02895856, 0.02018619, -0.02003199, -0.03201109, -0.08534801, 
    -0.2743452, -0.3680954, -0.4299279, -0.4045212, -0.4960415, -0.6135063, 
    -0.5829887, -0.6184213, -0.4850879, -0.3539674, -0.4234176, 0.1043491, 
    0.1734085,
  0.4596553, 0.5609086, 0.4730669, 0.27961, 0.07926813, -0.06915306, 
    -0.1222292, -0.06057558, 0.09564187, 0.2809284, 0.3645709, 0.5017779, 
    0.5532753, 0.49058, 0.3919147, 0.2473183, 0.09723687, -0.0368126, 
    -0.1266727, -0.2511355, -0.2830528, -0.2929812, -0.3039024, -0.305693, 
    -0.2845665, -0.2241664, -0.1296024, 0.0112831, 0.1301145, 0.1653847, 
    0.1099811, -0.00800398, -0.1753217, -0.3011843, -0.4021771, -0.4049278, 
    -0.3610313, -0.4152305, -0.5193809, -0.4776655, -0.3261192, -0.266142, 
    -0.2455854, -0.2797488, -0.3364708, -0.3926231, -0.4458784, -0.4823205, 
    -0.500387, -0.5249799, -0.510592, -0.4300745, -0.3137496, -0.1864873, 
    -0.07183897, 0.0366087, 0.1093137, 0.1408727, 0.145528, 0.1700069, 
    0.1973996, 0.2576047, 0.3503131, 0.3494342, 0.3664427, 0.4019895, 
    0.4460325, 0.5310097, 0.6083372, 0.7230833, 0.7111529, 0.6497272, 
    0.6499225, 0.5397499, 0.4608437, 0.3055538, 0.2713578, 0.2327183, 
    0.1629918, 0.08901733, 0.07705462, 0.01325226, -0.09003544, -0.2067673, 
    -0.2872686, -0.3659306, -0.3976198, -0.2950648, -0.3027956, -0.471514, 
    -0.5965302, -0.5194631, -0.4489224, -0.2442183, -0.1001263, -0.06021762,
  0.06242251, 0.06447315, 0.1717484, 0.1914912, -0.009517789, -0.04298121, 
    -0.06431913, -0.01340759, 0.07858443, 0.1686398, 0.292647, 0.3069048, 
    0.2886593, 0.2034054, 0.117175, -0.02128524, -0.07670522, -0.1519819, 
    -0.199573, -0.2160769, -0.2269331, -0.1904584, -0.1829064, -0.2094851, 
    -0.2074506, -0.1592898, -0.1266075, -0.07524031, -0.02969994, 
    0.004951764, 0.02710346, -0.03191347, -0.1009564, -0.2131309, -0.3035606, 
    -0.3348432, -0.3557742, -0.3838503, -0.3960248, -0.4021609, -0.3665001, 
    -0.3418418, -0.3219688, -0.3210411, -0.3479454, -0.3761355, -0.400045, 
    -0.4248823, -0.4647586, -0.4979454, -0.5201461, -0.5345992, -0.511731, 
    -0.4671673, -0.4063437, -0.3518515, -0.2881148, -0.2020795, -0.1147425, 
    -0.06041312, 0.004463196, 0.05898821, 0.1286334, 0.2497434, 0.3892128, 
    0.3805865, 0.4238157, 0.4732949, 0.5096555, 0.5425657, 0.5704953, 
    0.5521035, 0.5109576, 0.340401, 0.3213092, 0.2451861, 0.1813027, 
    0.0526894, -0.01195905, -0.0227989, -0.1069137, -0.1972133, -0.2542605, 
    -0.211113, -0.1713508, -0.1140751, -0.01215436, 0.1119665, 0.1944046, 
    0.1609733, 0.02052736, -0.05011082, -0.08160424, -0.08305287, 
    -0.05924082, -0.005920649,
  0.09230494, 0.06994164, 0.07096708, 0.0879432, -0.04566687, -0.03728461, 
    -0.003202677, 0.002803326, 0.0511269, 0.07344127, 0.08423209, 0.09419322, 
    0.08623409, 0.05560267, 0.01961637, -0.02621686, -0.07735622, -0.1320112, 
    -0.1828087, -0.2099572, -0.2180951, -0.219381, -0.2164024, -0.1757775, 
    -0.09229758, -0.04999615, -0.02025983, 0.01956764, 0.03086323, 0.0372597, 
    0.01766336, -0.009891987, -0.04584576, -0.09314394, -0.1572064, 
    -0.1914838, -0.2069786, -0.2233035, -0.2412885, -0.2449669, -0.2486452, 
    -0.2457971, -0.2501915, -0.2576134, -0.2833295, -0.3240847, -0.3726524, 
    -0.4255821, -0.4640749, -0.522392, -0.5676231, -0.5915815, -0.5938275, 
    -0.5636355, -0.5281538, -0.4711388, -0.4110802, -0.3073692, -0.2084271, 
    -0.1191368, -0.0481407, 0.03572971, 0.1247923, 0.2014849, 0.278438, 
    0.3484738, 0.4324906, 0.5034705, 0.5529497, 0.6037146, 0.6158078, 
    0.5415891, 0.4816932, 0.297888, 0.2481484, 0.1765663, 0.0890336, 
    0.02659857, -0.07597315, -0.1373825, -0.1702437, -0.2005332, -0.1615198, 
    -0.1174444, -0.05448854, 0.03003311, 0.1384153, 0.2378456, 0.3553098, 
    0.3841507, 0.3320186, 0.2378778, 0.2335811, 0.1986364, 0.1458368, 
    0.1050979,
  0.4043821, 0.3753294, 0.3432655, 0.29058, 0.2659056, 0.2247434, 0.1794472, 
    0.1423703, 0.101843, 0.05513078, 0.0009641051, -0.05619735, -0.1184857, 
    -0.1755658, -0.2179161, -0.2419071, -0.248808, -0.26331, -0.268144, 
    -0.2592084, -0.2458132, -0.2335737, -0.2137168, -0.186487, -0.1650841, 
    -0.1328738, -0.1026166, -0.09293236, -0.07740501, -0.07333599, 
    -0.07494733, -0.08324811, -0.09994733, -0.130709, -0.1623822, -0.1953575, 
    -0.2132611, -0.223515, -0.2380007, -0.2465619, -0.2563438, -0.2611452, 
    -0.2636355, -0.2698367, -0.2847455, -0.3058881, -0.3302696, -0.3546348, 
    -0.3798302, -0.3975548, -0.4086062, -0.4166628, -0.4204389, -0.4197553, 
    -0.4108523, -0.386959, -0.3530561, -0.3043582, -0.2542768, -0.2086225, 
    -0.1523237, -0.1091433, -0.06269151, -0.007466912, 0.05828834, 0.1249225, 
    0.1834999, 0.2356809, 0.2779335, 0.3066933, 0.3034544, 0.3023801, 
    0.2694374, 0.2119668, 0.1648638, 0.1417031, 0.1244992, 0.09264696, 
    0.06852591, 0.0675329, 0.07568741, 0.06631243, 0.07331115, 0.07109755, 
    0.08065164, 0.09901101, 0.1409706, 0.1838743, 0.2310422, 0.3334674, 
    0.3879921, 0.4258339, 0.4392291, 0.43975, 0.4437864, 0.4250038,
  0.3996458, 0.399955, 0.3976113, 0.3908893, 0.3790078, 0.3633014, 0.3433306, 
    0.3214719, 0.296472, 0.2663287, 0.2424518, 0.2216835, 0.1928587, 
    0.1683307, 0.1357298, 0.1005247, 0.06476621, 0.03102598, 0.0008339137, 
    -0.02139915, -0.04740826, -0.07406842, -0.0967735, -0.1088991, 
    -0.1155886, -0.1350873, -0.1508588, -0.1611452, -0.1742963, -0.1819297, 
    -0.1856732, -0.191793, -0.18289, -0.1874148, -0.2029584, -0.2151005, 
    -0.2361941, -0.2490196, -0.2583132, -0.2677696, -0.2845339, -0.3015423, 
    -0.3081016, -0.3129356, -0.3222455, -0.334127, -0.3396446, -0.3465945, 
    -0.3501752, -0.3628379, -0.369088, -0.3720177, -0.3733197, -0.3776329, 
    -0.3753217, -0.377991, -0.3775352, -0.3732221, -0.3636843, -0.3563113, 
    -0.3386844, -0.3212364, -0.2997358, -0.2859662, -0.2624962, -0.2388308, 
    -0.2122521, -0.1924116, -0.1725873, -0.1507286, -0.1364545, -0.1230756, 
    -0.1058393, -0.09294862, -0.07856061, -0.05928978, -0.04257428, 
    -0.02698183, -0.007873751, 0.01348041, 0.03349994, 0.05753966, 
    0.08236062, 0.1109576, 0.138985, 0.1686236, 0.2019407, 0.2355507, 
    0.2647825, 0.2953489, 0.3229368, 0.3460976, 0.3728717, 0.3911497, 
    0.3988157, 0.4046588,
  0.003294468, -0.01947546, -0.04146385, -0.06446171, -0.08739471, 
    -0.1103773, -0.1338305, -0.1568122, -0.1807542, -0.2046638, -0.2270761, 
    -0.2494073, -0.2717705, -0.2937753, -0.315048, -0.3345304, -0.351506, 
    -0.3656979, -0.3779869, -0.389201, -0.4001876, -0.410816, -0.4208258, 
    -0.4290614, -0.4346114, -0.4362878, -0.4325601, -0.4222901, -0.4051027, 
    -0.3801684, -0.3482671, -0.3101001, -0.2657156, -0.2156835, -0.1626883, 
    -0.1069102, -0.04890156, 0.008324623, 0.06496429, 0.1192288, 0.169425, 
    0.2157149, 0.2572842, 0.2928309, 0.3216715, 0.3441825, 0.3649664, 
    0.3739171, 0.364542, 0.3541093, 0.3483477, 0.3283267, 0.3061919, 
    0.3471594, 0.3113198, 0.3207107, 0.3445716, 0.3466702, 0.2885327, 
    0.1649489, 0.1793532, 0.2555575, 0.1687088, 0.1592522, 0.1348708, 
    0.1152906, 0.1016512, 0.09636116, 0.09405041, 0.0836978, 0.08858156, 
    0.1012931, 0.1195059, 0.1334057, 0.1743727, 0.1983962, 0.2196856, 
    0.2830319, 0.2777586, 0.3015046, 0.3167219, 0.3264878, 0.3294833, 
    0.3267655, 0.3188558, 0.3043861, 0.2849199, 0.2610915, 0.2342523, 
    0.204614, 0.1733483, 0.1422606, 0.1118729, 0.08208752, 0.05366969, 
    0.02730274,
  -0.04152822, -0.03868055, -0.03443241, -0.03363562, -0.03741074, 
    -0.04621649, -0.05653572, -0.07037115, -0.08514881, -0.107496, -0.137867, 
    -0.1719003, -0.2055588, -0.2372158, -0.2667234, -0.2899005, -0.3020103, 
    -0.3035077, -0.2989993, -0.2892337, -0.2875087, -0.2959397, -0.3204026, 
    -0.3563237, -0.3947186, -0.4250245, -0.4393802, -0.433326, -0.4080002, 
    -0.3654711, -0.3081465, -0.2373142, -0.1566987, -0.07043505, 0.01457357, 
    0.0932703, 0.1634178, 0.2253313, 0.2769423, 0.3187075, 0.3639555, 
    0.352644, 0.3224354, 0.3237877, 0.3187084, 0.2433825, 0.2911043, 
    0.2734284, 0.2385325, 0.1913805, 0.2523024, 0.1887772, 0.1817944, 
    0.2032793, 0.1846437, 0.2689047, 0.2729248, 0.251505, 0.2394607, 
    0.1848058, 0.1432214, 0.08098149, 0.006144285, -0.06791234, -0.1058836, 
    -0.1208742, -0.1310463, -0.1471438, -0.1673589, -0.195663, -0.2285565, 
    -0.2239828, -0.1820078, -0.1260834, -0.03270721, 0.06068468, 0.1352782, 
    0.221508, 0.2596593, 0.2678785, 0.3019767, 0.3004959, 0.240063, 
    0.2319252, 0.2091874, 0.1794021, 0.1633866, 0.1408936, 0.1121008, 
    0.08156681, 0.04916, 0.01660872, -0.008065224, -0.0244875, -0.03422022, 
    -0.0406661,
  -0.01262236, -0.05707264, -0.1009536, -0.1357512, -0.1600835, -0.176831, 
    -0.1970136, -0.2061447, -0.2163824, -0.2350997, -0.2546955, -0.2688396, 
    -0.2834072, -0.3054771, -0.3351655, -0.3481536, -0.3286057, -0.2860115, 
    -0.2347417, -0.1872152, -0.1573491, -0.1508877, -0.1501389, -0.1669846, 
    -0.2084072, -0.292017, -0.392912, -0.4463787, -0.4393642, -0.385653, 
    -0.3050218, -0.2125084, -0.1272709, -0.0627203, -0.01973581, 0.01024437, 
    0.02871799, 0.03392649, 0.0263586, 0.0135169, 0.0007400513, -0.02626181, 
    -0.06610632, -0.06415224, -0.09100819, -0.1591561, -0.1842041, 
    -0.1633384, -0.09224439, 0.007364988, 0.1265541, 0.2532957, 0.3850175, 
    0.5267327, 0.665535, 0.751668, 0.7437418, 0.7973869, 0.7180574, 
    0.5888901, 0.4149323, 0.2087317, -0.01133728, -0.1952891, -0.3511155, 
    -0.4799404, -0.6024333, -0.6981369, -0.7625737, -0.7888265, -0.787395, 
    -0.7500577, -0.6553149, -0.4774494, -0.3566179, -0.2228451, -0.06914902, 
    -0.01327419, 0.06107521, 0.1324773, 0.1792879, 0.1881106, 0.1750407, 
    0.1507076, 0.1616612, 0.1784906, 0.1913977, 0.1782305, 0.1470134, 
    0.04444098, 0.06061935, 0.032722, 0.03417015, 0.03952551, 0.0362215, 
    0.02411222,
  -0.1513593, -0.1804121, -0.1870854, -0.1823492, -0.1940029, -0.2448654, 
    -0.33383, -0.4178145, -0.4765551, -0.510931, -0.4653897, -0.3360605, 
    -0.1584888, 0.02406311, 0.1382718, 0.1873121, 0.1538968, 0.09019303, 
    0.03480649, -0.01478738, -0.02062988, -0.01058841, 0.004141331, 
    0.01047277, 0.000333786, -0.05218971, -0.1558191, -0.2202882, -0.1796632, 
    -0.07793832, 0.03565264, 0.1105387, 0.1470134, 0.1717691, 0.1908121, 
    0.198755, 0.1953368, 0.2057369, 0.2271724, 0.2653067, 0.3097076, 
    0.3085036, 0.3536534, 0.3584709, 0.3507071, 0.3401108, 0.2162175, 
    0.2299066, 0.2909257, 0.3266354, 0.3897865, 0.4665769, 0.5814856, 
    0.7030511, 0.8105381, 0.8896074, 0.9270101, 0.9015867, 0.7597737, 
    0.4984455, 0.2929931, 0.1115639, -0.04719299, -0.2388108, -0.4432702, 
    -0.6396891, -0.7556887, -0.8779058, -0.9145432, -0.8351326, -0.7002044, 
    -0.5556569, -0.4128184, -0.2809658, -0.23982, -0.2319589, -0.2298918, 
    -0.2581952, -0.2704351, -0.2552004, -0.1796956, -0.002449751, 0.1084715, 
    0.2411376, 0.336759, 0.3900304, 0.3974847, 0.3581294, 0.2947994, 
    0.1963948, 0.1038327, 0.1163006, 0.07603312, 0.05529737, -0.006095886, 
    -0.09950376,
  -0.1649826, -0.1806073, -0.1019135, -0.09794235, -0.09686756, -0.1645594, 
    -0.3163023, -0.4741955, -0.535573, -0.6303482, -0.5409927, -0.3854909, 
    -0.1933517, -0.007235289, 0.09322023, 0.0775795, -0.002156258, 
    -0.0644455, -0.1541591, -0.1363044, -0.02806863, 0.07556176, 0.1246982, 
    0.125155, 0.09728944, 0.05314898, -0.01871014, -0.1053805, -0.13134, 
    -0.06778288, 0.04051781, 0.08949304, 0.07334709, 0.06221437, 0.07997084, 
    0.1051831, 0.1384511, 0.1897535, 0.2017336, 0.1780505, 0.1292233, 
    0.1001873, 0.08216906, 0.0577054, 0.0138588, 0.1408763, 0.2258697, 
    0.3655026, 0.4357502, 0.4284748, 0.4447182, 0.477335, 0.544018, 
    0.6076735, 0.6789951, 0.7417067, 0.7677647, 0.7480382, 0.6683181, 
    0.5687575, 0.4634678, 0.3367101, 0.1495845, -0.0008063912, -0.1002365, 
    -0.1457115, -0.1633385, -0.1842043, -0.2154706, -0.276636, -0.06825387, 
    -0.09390485, -0.1273034, -0.2952233, -0.52605, -0.7032639, -0.7287521, 
    -0.7802658, -0.8644127, -0.9210371, -0.7370038, -0.6526936, -0.4722414, 
    -0.2236412, 0.02393365, 0.2120845, 0.3270746, 0.3619867, 0.3361403, 
    0.2981195, 0.3050694, 0.06535602, 0.02556092, -0.02548057, -0.08545709, 
    -0.1505136,
  0.5416585, 0.3533119, 0.3969971, 0.6123126, 0.6486566, 0.7199936, 0.751163, 
    0.863956, 1.070613, 1.066365, 0.7893958, 0.4363197, 0.06867671, 
    -0.2341394, -0.3025322, -0.1745205, -0.218955, -0.04530716, 0.2102451, 
    0.3264885, 0.2094314, 0.1915121, 0.08998215, -0.03583241, -0.1456304, 
    -0.2596288, -0.3391209, -0.3772736, -0.3779221, -0.3028407, -0.1650805, 
    -0.002776146, 0.1342525, 0.1589437, 0.1311264, 0.01073265, -0.08890963, 
    -0.09748602, -0.08925009, 0.03789854, 0.1041908, 0.07754564, 0.05350685, 
    0.0195713, -0.02816677, 0.1975007, 0.3951082, 0.5343339, 0.6353595, 
    0.6347246, 0.5419347, 0.5023676, 0.4930902, 0.4971103, 0.5591546, 
    0.5295323, 0.4562902, 0.4295486, 0.3962479, 0.2896723, 0.1697015, 
    0.007282928, -0.185816, -0.403622, -0.5366136, -0.6123948, -0.6767503, 
    -0.7703212, -0.9215908, -1.071379, -1.170175, -1.10385, -1.17273, 
    -1.178654, -1.193336, -1.18829, -1.19358, -1.065634, -0.9271082, 
    -0.8932377, -0.6970625, -0.6290775, -0.4632085, -0.2052171, 0.07923931, 
    0.271378, 0.3843663, 0.4142979, 0.4102615, 0.4199294, 0.3996658, 
    0.3464759, 0.3610433, 0.3914144, 0.4214599, 0.4346273,
  0.2190506, 0.07715601, -0.01052296, -0.03236461, -0.01296401, -0.00633955, 
    0.06823778, 0.2192295, 0.385278, 0.4111897, 0.1473061, -0.3147223, 
    -0.7590908, -0.8792404, -0.6741132, -0.4823494, -0.3228278, -0.1338472, 
    0.09894943, 0.2830801, 0.3426018, 0.2365472, 0.05492282, -0.1177654, 
    -0.2864342, -0.3632734, -0.4571867, -0.4695239, -0.4527433, -0.3980391, 
    -0.2632078, -0.1696045, -0.01931143, -0.09525633, -0.3801684, -0.4646246, 
    -0.277678, -0.2583261, -0.1801193, -0.1282959, -0.1464274, -0.1322348, 
    -0.04556441, -0.0364337, 0.137166, 0.2623289, 0.4954015, 0.6354405, 
    0.5573807, 0.2812414, 0.07245243, -0.06029499, -0.09745312, -0.0929935, 
    -0.1232669, -0.1652917, -0.1994224, -0.2204349, -0.2407311, -0.3490645, 
    -0.4865321, -0.6458257, -0.84301, -1.094605, -1.330868, -1.505819, 
    -1.652857, -1.828899, -2.054208, -2.240162, -2.292033, -2.271721, 
    -2.208309, -2.09677, -1.961434, -1.794719, -1.572128, -1.318287, 
    -1.132496, -1.051913, -0.7703538, -0.712053, -0.5198004, -0.2477464, 
    0.0828526, 0.3072993, 0.434936, 0.4871658, 0.5191157, 0.5793859, 
    0.5964758, 0.6445228, 0.7033935, 0.66062, 0.593595, 0.419897,
  -0.8415778, -0.9862554, -0.9971766, -0.8800216, -0.874683, -0.9641199, 
    -1.073999, -1.133683, -1.210327, -1.271249, -1.333488, -1.324618, 
    -1.213843, -1.11687, -1.086679, -1.086776, -1.042896, -0.8993083, 
    -0.738143, -0.5834719, -0.4948487, -0.4947184, -0.5650799, -0.7081465, 
    -0.7753338, -0.774097, -0.7396728, -0.7993246, -0.8898356, -0.8630782, 
    -0.648137, -0.3430751, -0.1354417, -0.09304261, -0.1493577, -0.2518642, 
    -0.3955979, -0.5716397, -0.7531822, -0.8822838, -0.9659425, -0.9779377, 
    -0.8792565, -0.6655197, -0.4156988, -0.2437422, -0.2097735, -0.2907305, 
    -0.4312416, -0.5847901, -0.6830974, -0.7152265, -0.7269289, -0.7471273, 
    -0.8651935, -0.9737221, -1.016919, -1.005005, -1.041854, -1.116203, 
    -1.120484, -1.099813, -1.187232, -1.402612, -1.590927, -1.587753, 
    -1.483879, -1.481421, -1.621184, -1.792506, -1.863729, -1.869295, 
    -1.861613, -1.857219, -1.911418, -1.973869, -1.950871, -1.776229, 
    -1.498202, -1.212314, -0.9754646, -0.8061773, -0.7086349, -0.5899665, 
    -0.46329, -0.3629319, -0.2527757, -0.1046962, 0.05606222, 0.1865961, 
    0.2811109, 0.3260491, 0.2440178, 0.06467226, -0.2408941, -0.5699143,
  -0.7092859, -0.5700766, -0.4166913, -0.4140217, -0.5783129, -0.7248621, 
    -0.7510178, -0.7128017, -0.6775646, -0.6897547, -0.6662197, -0.5467534, 
    -0.4527595, -0.4663012, -0.5983486, -0.7366295, -0.7632245, -0.6756915, 
    -0.621102, -0.7154379, -0.9078049, -1.04677, -1.079127, -1.081535, 
    -1.048104, -0.9465746, -0.7920659, -0.699471, -0.6816975, -0.6470785, 
    -0.5112708, -0.3594325, -0.2765713, -0.2669034, -0.3449957, -0.4478121, 
    -0.6182065, -0.8463144, -1.003215, -1.055705, -1.032855, -0.9679127, 
    -0.8916919, -0.8232672, -0.7640228, -0.7771571, -0.8435144, -0.9261317, 
    -1.017196, -1.114999, -1.217407, -1.3559, -1.581096, -1.779566, -1.87815, 
    -1.868108, -1.724488, -1.602727, -1.583407, -1.56163, -1.452694, 
    -1.271021, -1.2337, -1.390568, -1.38606, -1.1226, -0.9161868, -1.071346, 
    -1.349976, -1.537964, -1.603866, -1.63466, -1.642001, -1.680249, 
    -1.786466, -1.85424, -1.729126, -1.439949, -1.140503, -0.9106039, 
    -0.711499, -0.5424235, -0.4832766, -0.5027592, -0.5518804, -0.5481369, 
    -0.4767665, -0.3766038, -0.2750087, -0.1487555, -0.01039286, 0.001488656, 
    -0.1380784, -0.3934169, -0.6307378, -0.7426844,
  -0.3798418, -0.3753991, -0.457968, -0.6503994, -0.845046, -0.941659, 
    -0.9054937, -0.7394943, -0.5871835, -0.4809332, -0.4342537, -0.4610114, 
    -0.5446382, -0.5942149, -0.5583425, -0.4916103, -0.4960372, -0.5720463, 
    -0.7110598, -0.8962001, -1.058748, -1.117522, -1.071574, -0.9624594, 
    -0.8419842, -0.7324952, -0.6591065, -0.6138102, -0.5908444, -0.587769, 
    -0.5566003, -0.5860765, -0.7116299, -0.8633561, -0.9608655, -1.060182, 
    -1.179452, -1.1899, -1.107561, -1.008717, -0.9662032, -0.9718347, 
    -0.9672937, -0.8991139, -0.8416758, -0.9076424, -1.0747, -1.237151, 
    -1.394523, -1.525171, -1.579387, -1.684335, -1.943873, -2.069491, 
    -1.897681, -1.641138, -1.503508, -1.467717, -1.434107, -1.374553, 
    -1.253915, -1.117326, -1.066187, -1.028508, -0.776945, -0.4586018, 
    -0.4634525, -0.7733808, -0.9838952, -1.005265, -1.026099, -1.210686, 
    -1.443107, -1.662183, -1.833277, -1.744116, -1.331276, -0.8639255, 
    -0.6646245, -0.6362226, -0.5995362, -0.477222, -0.3839931, -0.3524494, 
    -0.3479898, -0.2917559, -0.1717693, -0.02925634, 0.09265113, 0.1642328, 
    0.1654537, 0.03566849, -0.1715418, -0.3253989, -0.3773521, -0.3803632,
  -0.1297777, -0.2300549, -0.4251065, -0.5612564, -0.5464778, -0.4441338, 
    -0.3028078, -0.1782475, -0.0755949, -0.04393816, -0.1180587, -0.214787, 
    -0.2381434, -0.2189212, -0.2497001, -0.3864996, -0.5824308, -0.7585211, 
    -0.8715088, -0.8991296, -0.8484133, -0.7263429, -0.6430745, -0.6592857, 
    -0.6695068, -0.6487224, -0.6129473, -0.5232012, -0.43606, -0.4620206, 
    -0.580966, -0.702239, -0.8234463, -0.8634844, -0.8349533, -0.8529549, 
    -0.9514728, -1.011727, -1.014917, -0.9893966, -0.9089928, -0.8176031, 
    -0.7524507, -0.6927662, -0.7177174, -0.940048, -1.1434, -1.209367, 
    -1.305542, -1.404615, -1.36381, -1.355201, -1.503899, -1.504241, 
    -1.218726, -1.022144, -1.111125, -1.225708, -1.14187, -0.9952885, 
    -0.8399012, -0.6773033, -0.5168049, -0.3444254, -0.08827305, 0.05694175, 
    0.02927256, -0.06382656, -0.1278725, -0.3094318, -0.6329505, -0.9812584, 
    -1.273153, -1.472323, -1.44983, -1.111582, -0.5726333, -0.2635016, 
    -0.2270918, -0.3222572, -0.3012612, -0.1702561, -0.06174374, -0.06384254, 
    -0.07572412, -0.04452312, 0.02219236, 0.09802222, 0.1037519, 0.06997859, 
    0.01652813, -0.05067575, -0.09875512, -0.08119321, -0.07085752, 
    -0.08594561,
  0.1014233, -0.03811097, -0.1923101, -0.2529883, -0.2105241, -0.1283951, 
    -0.04514313, 0.02949953, 0.04361057, 0.01473713, -0.03908777, -0.1195402, 
    -0.1562757, -0.1901941, -0.308521, -0.4599857, -0.5021405, -0.4690514, 
    -0.459725, -0.4663984, -0.4330159, -0.3977789, -0.4797448, -0.7208741, 
    -0.8991621, -0.8483965, -0.6996338, -0.5598392, -0.5047615, -0.6611581, 
    -0.8593524, -0.8720789, -0.8144617, -0.7739997, -0.7392178, -0.766366, 
    -0.7797613, -0.719296, -0.6502371, -0.5616961, -0.4228935, -0.3411059, 
    -0.4179289, -0.5829837, -0.7327397, -0.8119879, -0.7896245, -0.706714, 
    -0.7393965, -0.7654871, -0.6679611, -0.598202, -0.6043869, -0.5791753, 
    -0.5880296, -0.696916, -0.8109298, -0.7860273, -0.6426517, -0.4441652, 
    -0.1849365, 0.05327964, 0.2020915, 0.3075278, 0.4762776, 0.5838294, 
    0.5905681, 0.5604081, 0.3249106, -0.1728432, -0.5643148, -0.7544355, 
    -0.9707932, -1.169214, -0.9707117, -0.467782, -0.05920458, 0.09794092, 
    0.07368898, 0.004012108, -0.05000806, 0.01380944, 0.06737375, 0.05471206, 
    0.06651187, 0.1047444, 0.1736246, 0.2453041, 0.2416583, 0.1881914, 
    0.1933672, 0.1921791, 0.1960202, 0.2097574, 0.1885011, 0.15118,
  0.302367, 0.0703361, -0.02388597, 0.02606535, 0.09061623, 0.21018, 
    0.3681879, 0.4482496, 0.3754797, 0.2619054, 0.08646607, -0.1494226, 
    -0.2570727, -0.3222091, -0.4511151, -0.4813884, -0.4865316, -0.4816651, 
    -0.428589, -0.37203, -0.3521244, -0.4632246, -0.6516525, -0.7562094, 
    -0.6907473, -0.4377358, -0.2515712, -0.2699957, -0.3176517, -0.3689868, 
    -0.3620694, -0.2629163, -0.2652602, -0.3330822, -0.3004165, -0.1831474, 
    -0.06796169, 0.004076481, 0.04742002, 0.05378342, -0.03967333, 
    -0.1373458, -0.2166748, -0.3215088, -0.303833, -0.2316325, -0.1476647, 
    -0.1703534, -0.1600349, -0.1084234, -0.05181533, -0.1126389, -0.1199142, 
    -0.1885338, -0.4685633, -0.6564212, -0.4656821, -0.2201582, -0.05596542, 
    0.1723875, 0.4662188, 0.6736407, 0.6721759, 0.7114991, 0.8728598, 
    0.9384195, 0.882804, 0.7704179, 0.507869, 0.1415286, -0.08604383, 
    -0.219898, -0.3874435, -0.4381921, -0.1307371, 0.3126864, 0.5572667, 
    0.5434158, 0.4113848, 0.2749107, 0.1758385, 0.2826414, 0.400301, 
    0.3759199, 0.3671144, 0.3808513, 0.3699785, 0.4745196, 0.5380775, 
    0.4613849, 0.3687253, 0.2930417, 0.3148354, 0.3883708, 0.4138261, 
    0.4245846,
  0.2354083, 0.08345556, 0.1359451, 0.2077067, 0.3621011, 0.6026773, 
    0.5875568, 0.3404212, 0.08924913, -0.3324144, -0.7570562, -0.9112225, 
    -0.7700768, -0.7219645, -0.7511477, -0.648039, -0.4966556, -0.2805912, 
    -0.07303917, -0.04380757, -0.1103114, -0.202857, -0.1913497, 
    -0.0006432533, 0.1290932, 0.2049884, 0.1327721, -0.008976221, 
    0.009578466, 0.04269993, 0.009024858, -0.07766104, -0.2194095, 
    -0.1939378, 0.0541904, 0.2839429, 0.4125564, 0.5185299, 0.5445552, 
    0.3694737, 0.09089351, -0.000643611, 0.00630635, -0.02297422, 0.01037537, 
    0.01302837, 0.01924598, 0.1609613, 0.2693109, 0.2107334, 0.1999424, 
    0.2098708, 0.2238358, 0.1255935, -0.2102138, -0.2775153, -0.01545471, 
    0.2152909, 0.450545, 0.7198972, 0.9669025, 1.142277, 1.182772, 1.28492, 
    1.272909, 1.085018, 1.0038, 0.904126, 0.6499426, 0.3321533, 0.1534095, 
    0.09772921, 0.09714317, 0.1985595, 0.5369384, 1.037476, 1.401001, 
    1.097013, 0.4449627, 0.2324297, 0.4912679, 0.7014083, 0.7731364, 
    0.6492269, 0.4904703, 0.4636314, 0.4441978, 0.5411214, 0.5555743, 
    0.3930417, 0.32714, 0.3774656, 0.5232501, 0.6367429, 0.5629965, 0.4271562,
  0.2234614, 0.2250729, 0.4467526, 0.7952875, 1.185001, 1.298445, 0.8218829, 
    0.3954021, -0.03687382, -0.7601485, -0.873446, -0.3709393, -0.01861191, 
    0.004516602, 0.03332478, 0.271264, 0.3786371, 0.4740635, 0.5986403, 
    0.5522375, 0.4930252, 0.4902907, 0.5065342, 0.4916905, 0.2657302, 
    0.06996197, -0.02712462, 0.02850688, 0.2478916, 0.3768793, 0.4083411, 
    0.3407469, 0.3144772, 0.5475013, 0.8402421, 0.9098868, 0.8561924, 
    0.8922441, 0.7741127, 0.3518797, 0.1734615, 0.1861892, -0.01441288, 
    -0.1781499, -0.1628829, -0.08407432, 0.09196723, 0.3739495, 0.5169182, 
    0.4912837, 0.6015537, 0.6369379, 0.4992263, 0.2858311, 0.1183669, 
    0.2597894, 0.4978428, 0.5948154, 0.8571365, 1.039428, 1.093481, 1.201099, 
    1.248624, 1.20297, 0.8570554, 0.4852943, 0.461336, 0.5108155, 0.460441, 
    0.3634518, 0.3602291, 0.4191979, 0.4659586, 0.6550537, 0.9855871, 
    1.473999, 1.725349, 0.892342, 0.1317134, 0.143074, 0.6835525, 0.7504475, 
    0.7484945, 0.5253174, 0.2923423, 0.344686, 0.3727947, 0.3994385, 
    0.3854408, 0.3617591, 0.4208085, 0.473494, 0.5204666, 0.4660397, 
    0.3914466, 0.3283443,
  0.3401442, 0.4307531, 0.6129636, 1.047436, 1.140388, 0.6204015, 0.3238196, 
    0.3076575, -0.1481689, -0.8245363, -0.3148845, 0.3861892, 0.3883539, 
    0.3260655, 0.5106358, 0.7530349, 0.777384, 0.7032303, 0.7218175, 
    0.6767167, 0.5857989, 0.4541909, 0.3231035, 0.2017822, 0.04299319, 
    0.01623511, 0.09689939, 0.3566813, 0.631193, 0.8415772, 0.9983799, 
    0.7526771, 0.639282, 0.7240801, 0.7071859, 0.7015704, 0.7144282, 
    0.6154209, 0.3054112, 0.05371846, 0.1872799, 0.09585786, -0.2903565, 
    -0.4383708, -0.4053792, -0.08474147, 0.4146889, 0.7086666, 0.8483475, 
    0.8401935, 0.7077877, 0.492358, 0.4618891, 0.5541905, 0.5090083, 
    0.6135654, 0.7932531, 0.7782628, 0.8847407, 0.9546299, 0.9461502, 
    0.9920487, 0.8608476, 0.5605872, 0.1773031, 0.07668424, 0.3321531, 
    0.5738685, 0.7028239, 0.7050215, 0.6055256, 0.4342361, 0.473087, 
    0.8506587, 1.202205, 1.530932, 1.285652, 0.4330804, -0.07626188, 
    0.2455969, 0.7922928, 0.5755943, 0.4681723, 0.4291583, 0.219914, 
    0.2397376, 0.2001058, 0.1922767, 0.2820062, 0.4297439, 0.4590245, 
    0.411889, 0.3688227, 0.228572, 0.2854242, 0.3264562,
  0.4325112, 0.6309648, 0.7608471, 0.9992745, 0.5607502, -0.04100776, 
    -0.06094527, -0.05147302, -0.2236903, -0.1817633, 0.5509029, 0.7919999, 
    0.4972895, 0.5992588, 0.7931554, 0.8570718, 0.7851154, 0.6934001, 
    0.6190515, 0.4059167, 0.2596762, 0.198755, 0.2045002, 0.2197838, 
    0.1623774, 0.1589105, 0.3617103, 0.7211502, 0.93505, 1.116772, 1.108911, 
    0.6363845, 0.503751, 0.6038975, 0.4701573, 0.5289626, 0.5808019, 
    0.492505, 0.3396891, 0.1915767, 0.3025798, 0.242537, -0.08711815, 
    -0.2948492, -0.3134363, 0.05493975, 0.5352619, 0.6315506, 0.6381267, 
    0.4857829, 0.2584556, 0.3151613, 0.5194252, 0.6376542, 0.6016519, 
    0.6038818, 0.648413, 0.4707923, 0.4416581, 0.5714106, 0.6050531, 
    0.512182, 0.2719476, 0.1121005, 0.05962682, 0.2776119, 0.6324297, 
    0.8415931, 0.7965408, 0.5154861, 0.3951085, 0.2756587, 0.3983966, 
    0.8429115, 1.102351, 1.228035, 0.6609938, -0.04572797, -0.2633384, 
    0.0417558, 0.5285395, 0.4168704, 0.3667728, 0.3204993, -0.0174886, 
    -0.2035401, -0.06962132, 0.05414165, 0.1051345, 0.2632889, 0.3070879, 
    0.3110754, 0.3810463, 0.2709063, 0.3243895, 0.3317299,
  0.5177321, 0.5387602, 0.3915277, 0.2312412, -0.1284105, -0.2163491, 
    -0.1008707, -0.1719651, -0.05127827, 0.4199948, 0.9478915, 0.7469966, 
    0.4067465, 0.4503168, 0.5021074, 0.5080156, 0.3897049, 0.2767003, 
    0.3486569, 0.1659582, 0.06161261, 0.1386628, 0.1951571, 0.1998446, 
    0.1888583, 0.3521068, 0.6974356, 0.8322339, 0.8252513, 0.8174229, 
    0.5929118, 0.1724198, 0.1073318, 0.2072181, 0.230509, 0.4620523, 
    0.5342362, 0.3608475, 0.2491455, 0.2082926, 0.3443758, 0.3320708, 
    -0.09322262, -0.5056572, -0.3905528, 0.005247831, 0.3198643, 0.4141839, 
    0.3681388, 0.3853264, 0.51381, 0.6189535, 0.5600338, 0.4960854, 
    0.4821694, 0.3571042, 0.2406167, 0.147127, 0.2148353, 0.3822667, 
    0.298917, 0.1686762, 0.08583109, 0.1112706, 0.3017002, 0.6375076, 
    0.7146397, 0.6311761, 0.5510167, 0.3315668, 0.2886149, 0.2311114, 
    0.3969316, 0.6785719, 0.7650619, 0.7238193, 0.08924913, -0.09258682, 
    -0.1080325, -0.1482991, 0.2093501, 0.1698321, 0.1081132, 0.261352, 
    0.01460716, -0.2091722, -0.115243, 0.04686689, 0.1009359, 0.2316002, 
    0.256405, 0.2905028, 0.4021893, 0.3088462, 0.3327549, 0.3743565,
  0.2413969, 0.01950645, -0.2092047, -0.2625902, -0.09869033, 0.1586831, 
    0.2634027, 0.2961338, 0.3628656, 0.5534747, 0.8016994, 0.6560295, 
    0.2118729, 0.3158931, 0.511775, 0.4175532, 0.449796, 0.4249585, 
    0.5054431, 0.3432686, 0.05611062, -0.01394153, 0.1487703, 0.2355707, 
    0.2132883, 0.4137115, 0.5815015, 0.4257073, 0.3267815, 0.3198645, 
    0.1129636, -0.1297122, -0.008309603, 0.1655188, 0.1526449, 0.2154379, 
    0.298559, 0.1916904, 0.1823001, 0.1724193, 0.1450267, 0.03472424, 
    -0.3564219, -0.6874442, -0.5294037, -0.1516204, 0.1668694, 0.1825919, 
    0.1412346, 0.4636633, 0.5543537, 0.2856039, 0.1697022, 0.09162593, 
    -0.07333171, -0.2643963, -0.2119551, -0.0307703, 0.106697, 0.06511176, 
    -0.09917866, 0.005883157, 0.2015212, 0.3130447, 0.4065505, 0.5244379, 
    0.447729, 0.3021887, 0.2973386, 0.2720294, 0.2831624, 0.3016191, 
    0.5012119, 0.480655, 0.3993893, 0.4063067, 0.1505609, 0.2733636, 
    -0.004630566, -0.006632686, 0.2550206, 0.152742, 0.1289626, 0.2082758, 
    0.08866316, -0.09154463, -0.1423261, 0.003800154, 0.09227705, 0.1508539, 
    0.2332437, 0.330102, 0.4023514, 0.3134677, 0.2238355, 0.2469311,
  -0.1009531, -0.3718996, -0.3635349, -0.1078048, 0.1471104, 0.2296787, 
    0.2644118, 0.282641, 0.3209712, 0.3365151, 0.4965248, 0.3610263, 
    -0.1397058, 0.2287672, 0.6211166, 0.5295486, 0.5585675, 0.5927801, 
    0.5907133, 0.2596426, -0.04685116, -0.06286716, 0.2214589, 0.205101, 
    0.1004629, 0.2409904, 0.1957266, -0.05759358, -0.1737065, -0.1976645, 
    -0.2608968, -0.3067627, -0.2914963, -0.1657796, -0.1593668, -0.01008368, 
    -0.004810333, -0.321054, -0.1410568, -0.1121674, -0.2479739, -0.458847, 
    -0.6684661, -0.7782326, -0.6020925, -0.3049402, -0.139869, -0.1278408, 
    0.03781748, 0.3489662, 0.2468503, -0.1108971, -0.288957, -0.4886315, 
    -0.5161218, -0.3109788, -0.1526942, -0.09992731, 0.02897885, 0.03026474, 
    0.08749124, 0.2606196, 0.290421, 0.3582758, 0.3776445, 0.3225826, 
    0.3582761, 0.4260986, 0.3992429, 0.3702228, 0.4001215, 0.4215729, 
    0.5344143, 0.3926182, 0.3742104, 0.484756, 0.5198485, 0.2707758, 
    -0.1475016, 0.04286236, 0.2914138, 0.1193272, 0.1676833, 0.127156, 
    -0.0602293, -0.1883879, -0.05674696, 0.07399821, 0.121557, 0.2718987, 
    0.4530022, 0.4562738, 0.37976, 0.3027096, 0.2348547, 0.1438546,
  -0.4332285, -0.4727631, -0.3776946, -0.1245532, 0.05629009, 0.1878821, 
    0.2394284, 0.09859216, 0.2528239, 0.3168373, 0.2511473, 0.2240148, 
    -0.1342049, 0.2192135, 0.573802, 0.5691309, 0.5524974, 0.4793856, 
    0.4191315, -0.008521318, -0.1236253, -0.09610248, -0.03645134, 
    -0.1251063, -0.2711351, -0.260637, -0.3810954, -0.627108, -0.6173425, 
    -0.5547931, -0.5453854, -0.4042073, -0.3922604, -0.6540287, -0.5537193, 
    -0.1889899, -0.2381113, -0.327076, -0.02295732, -0.1421642, -0.4812918, 
    -0.6699467, -0.8910568, -0.7792244, -0.5010993, -0.4606693, -0.5246015, 
    -0.3102783, -0.0593183, 0.1644933, 0.1866612, -0.05920476, -0.311109, 
    -0.4060959, -0.1973395, 0.07577258, 0.1025141, 0.07352644, 0.1997635, 
    0.1944573, 0.2080806, 0.1894121, 0.1418536, 0.2282145, 0.3172282, 
    0.386499, 0.4428625, 0.442065, 0.4283929, 0.4367588, 0.4244366, 
    0.4311109, 0.3957438, 0.3143454, 0.2523503, 0.2192464, 0.05878049, 
    -0.04559755, -0.05508679, 0.1410235, 0.06013137, -0.0235275, 0.0439043, 
    -0.07357585, -0.1812255, -0.1042082, 0.01017952, -0.002905846, 0.1646883, 
    0.3968334, 0.3039951, 0.1910882, 0.1895418, 0.05389786, -0.06438112, 
    -0.2375584,
  -0.5085702, -0.551311, -0.5476978, -0.2992432, -0.1063888, -0.001912594, 
    0.01898599, -0.03900576, 0.1251057, -0.008211493, -0.03143764, 
    0.06919765, -0.0559659, 0.4447498, 0.4666743, 0.2229562, 0.227351, 
    -0.0550375, -0.2869387, -0.4281006, -0.5107827, -0.6082599, -0.6410403, 
    -0.6879153, -0.8773519, -0.6569908, -0.4916753, -0.611711, -0.5024498, 
    -0.6111249, -0.5881426, -0.592863, -0.6074463, -0.6594808, -0.5246508, 
    -0.6510501, -0.7112556, -0.5058193, -0.08508301, -0.1444423, -0.9507253, 
    -0.9403245, -0.9122152, -0.5281168, -0.3420167, -0.4932377, -0.3610925, 
    -0.0542078, -0.009709239, 0.2952387, 0.2902257, -0.03422081, -0.1737228, 
    -0.1443606, 0.01926225, 0.1920976, 0.2542558, 0.1550697, 0.140112, 
    0.1231524, 0.1411868, 0.1052655, 0.2061443, 0.3205976, 0.3849847, 
    0.4371333, 0.4134676, 0.3426182, 0.3031001, 0.2568426, 0.1511135, 
    0.1883378, 0.1553302, 0.1604733, 0.06563258, -0.01065329, -0.04610234, 
    -0.07004455, 0.04987752, 0.05030096, -0.06490132, 0.002286434, 
    -0.05565619, -0.1377683, -0.02954912, 0.02712369, 0.08591223, 0.04143, 
    0.1193433, 0.102612, 0.02611399, -0.06797767, -0.1419199, -0.321363, 
    -0.3993902, -0.4377203,
  -0.6549406, -0.5751224, -0.3061278, 0.04834807, 0.1164467, -0.2370201, 
    -0.2448163, -0.2368079, -0.1323001, -0.1982828, -0.1718676, 0.3201904, 
    0.413322, 0.5236731, 0.5997963, 0.431746, 0.3308022, 0.02313614, 
    -0.2864827, -0.4026937, -0.6781496, -0.7076741, -0.6022869, -0.8511476, 
    -0.9482992, -0.3479579, -0.1624111, -0.1340904, -0.1057863, -0.5012937, 
    -0.1689534, -0.1104736, -0.2854737, -0.5852785, -0.4571695, -0.2013593, 
    -0.01691914, -0.1429772, -0.03436747, -0.2092859, -1.421607, -0.9658612, 
    -0.6019779, -0.3149664, -0.3598395, -0.3332281, -0.0575771, 0.04598737, 
    0.04146266, 0.287589, 0.2792882, 0.1776769, 0.2715896, 0.2555577, 0.3281, 
    0.3843662, 0.3833083, 0.3519281, 0.3697993, 0.3775141, 0.3708896, 
    0.3110266, 0.2743896, 0.2806234, 0.3218832, 0.2475662, 0.2019281, 
    0.1991935, 0.1343009, 0.08960724, 0.01942492, -0.0806241, -0.1370203, 
    -0.2809007, -0.3170168, -0.06768453, -0.04081279, -0.1345789, -0.1235927, 
    -0.09165913, -0.0002689958, -0.0004319251, -0.06189026, -0.1019617, 
    -0.119849, -0.1231362, -0.05251455, 0.197664, 0.08207202, -0.06333828, 
    0.03052568, -0.344914, -0.6070397, -0.5269458, -0.6094491, -0.5837817,
  -0.3146728, -0.1539141, 0.02930462, 0.1567784, 0.1690668, -0.02871968, 
    -0.05046447, -0.08718322, -0.2615805, -0.2538664, -0.2053473, 0.5520096, 
    1.134203, 1.10297, 0.861547, 0.7090415, 0.3895097, 0.08199, -0.1961349, 
    -0.4971435, -0.5505294, -0.3114178, -0.3686934, -0.6224527, -0.4950445, 
    0.01752138, 0.03690553, -0.04802306, -0.3080002, -0.7999921, -0.03197467, 
    -0.03855026, -0.07761276, -0.7017171, -0.4504639, -0.0006435076, 
    -0.004142851, -0.02828023, -0.1645432, -0.7737877, -1.287704, -0.5163172, 
    -0.2833258, -0.201734, -0.4102137, -0.3196212, -0.1573489, -0.003768086, 
    0.1261312, 0.1669515, 0.1796958, 0.2004967, 0.2875084, 0.2772056, 
    0.3008705, 0.3350505, 0.3449788, 0.3771241, 0.3875241, 0.4059485, 
    0.3940017, 0.3634191, 0.3149652, 0.2849685, 0.1771886, 0.075203, 
    0.02728653, -0.04750168, -0.04239118, -0.153231, -0.2044191, -0.2264892, 
    -0.2247318, -0.334969, -0.2872809, -0.004386991, -0.005428672, 
    -0.08335835, -0.1396084, -0.1586351, -0.09546775, 0.06849714, 0.1435134, 
    -0.0873785, -0.1577724, -0.09719299, 0.07723734, 0.365014, 0.2615635, 
    0.1812088, 0.1377192, -0.2628014, -0.2444907, -0.004223347, -0.1171632, 
    -0.1408772,
  -0.1402264, 0.06778157, 0.05972433, -0.01771708, 0.09960064, 0.1390538, 
    0.1306716, 0.1079014, -0.03890812, -0.1858478, -0.1494224, 0.3252187, 
    0.8115473, 1.296167, 1.122158, 0.6864988, 0.4399654, -0.005038042, 
    -0.1881435, -0.373739, -0.2630942, -0.1559823, -0.2890389, -0.3496504, 
    -0.3421627, 0.02985779, 0.3414626, -0.06942606, -1.169247, -1.29257, 
    -0.3846116, -0.06055562, -0.1001552, -0.6141037, -0.4159918, -0.2738042, 
    -0.3125573, 0.01162863, -0.2225509, -0.5276779, -0.3507086, -0.07458538, 
    -0.0006270409, 0.1282793, 0.07015765, 0.04230952, 0.07456839, 0.2096596, 
    0.2539631, 0.1836667, 0.147306, 0.02349436, -0.02204585, -0.06250823, 
    -0.1207438, -0.1124108, -0.116138, -0.1587, -0.1959721, -0.1565353, 
    -0.1114182, -0.09911358, -0.1119391, -0.09878803, -0.1182542, 
    -0.06431532, -0.04366064, -0.1111249, -0.09748566, -0.1461185, 
    -0.06390828, -0.03291875, -0.04982954, 0.08465958, 0.1583246, -0.1319749, 
    -0.2737391, -0.1382249, -0.01538959, 0.01516053, -0.04393778, -0.0583909, 
    -0.1005619, 0.05189538, 0.131958, 0.2517986, 0.2795815, 0.3092368, 
    0.2747639, 0.2809809, 0.103458, -0.1400313, -0.05474472, 0.03094864, 
    -0.0538168, -0.07543135,
  0.1767008, 0.2776282, 0.1462153, 0.04064882, 0.04940546, 0.1613358, 
    0.1788648, 0.2656162, 0.3026769, -0.03576721, -0.1087161, 0.3184481, 
    0.5451565, 1.062296, 1.221444, 0.6567631, 0.4375076, 0.06691834, 
    0.00782004, -0.08596253, 0.01058733, -0.07665277, -0.1968517, -0.4487724, 
    -0.6126554, -0.4760988, -0.1180914, 0.009545296, -0.5227457, -1.153524, 
    -0.8921148, -0.30079, -0.3610926, -0.3363851, -0.4430751, -0.2649664, 
    -0.1455979, 0.0510492, 0.00798279, 0.0459224, 0.1715084, 0.09034002, 
    0.2881589, 0.3662353, 0.4632894, 0.4657145, 0.3538327, 0.3209717, 
    0.3077714, 0.3941641, 0.3779378, 0.3704834, 0.2672281, 0.155021, 
    0.03500128, -0.08526206, -0.1836506, -0.2360274, -0.2608966, -0.3581787, 
    -0.4174889, -0.4507409, -0.4165777, -0.3655361, -0.2392991, -0.1721116, 
    -0.1071863, -0.04161018, -0.1224533, -0.06862837, -0.05534714, 
    -0.03337449, -0.02131405, 0.1007075, 0.3022869, 0.02005962, -0.005998313, 
    0.1019776, -0.0581142, -0.1703376, -0.2434978, -0.1923263, -0.003719807, 
    0.2214756, 0.313875, 0.3646557, 0.31656, 0.2842848, 0.2636142, 0.2781656, 
    0.1727293, -0.1016526, -0.2008877, 0.01540482, 0.1009841, 0.08255994,
  -0.07622886, 0.02862144, 0.1584063, 0.2863196, 0.2667233, 0.6080813, 
    0.6410725, 0.4995195, 0.6882241, 0.6050371, 0.06123817, 0.1117918, 
    0.7717032, 0.820385, 1.209936, 0.9482985, 0.566007, 0.3488845, 0.1898682, 
    -0.03959167, 0.06862736, -0.04016161, -0.1570878, -0.4615483, -0.8260345, 
    -1.381601, -1.165829, 0.09543407, 0.5544187, -0.582772, -1.352173, 
    -1.281454, -1.125513, -0.253622, -0.6526615, -0.7002853, -0.38593, 
    -0.1416266, 0.07171977, 0.07071078, 0.1148353, 0.01276851, 0.3037355, 
    0.3225503, 0.392195, 0.4777093, 0.485359, 0.4308181, 0.357511, 0.3473384, 
    0.2333083, 0.244132, 0.1818762, 0.228621, 0.2030025, 0.1729403, 
    0.1292396, -0.02883339, -0.1108811, -0.1237879, -0.1164315, -0.2690845, 
    -0.2960374, -0.2823818, -0.2352786, -0.2698812, -0.208716, -0.104387, 
    -0.1437913, -0.07554586, -0.2235276, -0.01296449, -0.04151249, 
    -0.4112384, -0.1496342, -0.2354741, -0.3893803, -0.5562419, -0.6990645, 
    -0.5967369, -0.5750902, -0.333293, -0.09644413, 0.1651928, 0.2169023, 
    0.24545, 0.3269444, 0.3477452, 0.3383536, 0.357218, 0.4139731, 0.1272215, 
    -0.180591, 0.02813292, 0.1666909, -0.02108574,
  0.5002031, 0.3971273, 0.1673417, 0.1199131, -0.1235765, -0.1963141, 
    -0.2045009, -0.1441005, -0.3406988, -0.1913336, -0.4069261, -0.4437424, 
    0.1367757, 0.22771, 0.7250404, 0.9969141, 0.5655349, 0.3432367, 
    0.3147057, 0.20979, 0.2310622, 0.4371338, 0.3169994, -0.1680598, 
    -0.6150312, -1.341903, -1.076473, -0.1053307, 0.1400793, -0.07276237, 
    -0.516561, -1.55258, -1.867375, -0.893775, -1.178182, -1.324878, 
    -0.8481857, -0.4168707, -0.1930752, -0.1416265, -0.03208864, -0.1626874, 
    0.0809654, 0.2382567, 0.2011147, 0.1999266, 0.2536044, 0.2014885, 
    0.107657, 0.002253771, -0.07136297, -0.1350834, -0.1875575, -0.1504478, 
    -0.1665611, -0.1285405, -0.05752802, -0.03423691, -0.04737186, 
    -0.04497957, 0.01904964, -0.008505821, -0.06779957, -0.08617449, 
    -0.123023, -0.209579, -0.2600999, -0.3120198, -0.1379155, -0.1095953, 
    -0.2106533, 0.1037185, 0.06490028, -0.2312427, -0.174439, -0.544426, 
    -0.8561771, -0.8275473, -0.7160566, -0.703687, -0.7396082, -0.5189699, 
    -0.3231044, -0.1374114, 0.01698351, 0.1002517, 0.1832266, 0.2458081, 
    0.3683667, 0.4995189, 0.7823315, 0.7440178, 0.6570063, 0.6803465, 
    0.8497311, 0.7779702,
  0.7247797, 0.6759353, 0.4150465, 0.3571203, 0.1500728, -0.2304934, 
    -0.5642664, -0.4726162, -0.6147225, -0.7249439, -0.6109626, -0.5684652, 
    -0.0224534, -0.08594625, 0.1362875, 0.3875403, 0.3832443, 0.3232822, 
    0.3911539, 0.3233969, 0.4283612, 1.280721, 1.365127, -0.001653194, 
    -0.6580658, -0.6804612, -0.3092526, -0.2161868, -0.1842535, 0.4676673, 
    0.3766029, -0.8118735, -1.099862, -0.959188, -1.516463, -1.484449, 
    -1.089445, -0.7915288, -0.4416103, -0.1716722, -0.2696214, -0.3920007, 
    -0.174455, -0.03882647, -0.01426601, 0.03057432, -0.01804209, 
    -0.06488514, -0.04418182, -0.1605394, -0.2550378, -0.3598881, -0.3316495, 
    -0.2855394, -0.2015712, -0.2365649, -0.258033, -0.1934497, -0.2496994, 
    -0.2538824, -0.2962332, -0.2452731, -0.3241467, -0.3163991, -0.3430748, 
    -0.3108811, -0.3169694, -0.4472907, 0.004157901, 0.0003005043, 
    -0.05354065, 0.1499424, 0.06947386, 0.4169026, 0.3711993, 0.003669649, 
    -0.3244552, -0.6819097, -1.008244, -1.023332, -0.8322839, -0.6265059, 
    -0.4190025, -0.3101318, -0.1567309, -0.06301355, 0.02950001, 0.05944681, 
    0.09676933, 0.183064, 0.2627354, 0.34091, 0.1551831, 0.3158125, 
    0.8475341, 0.9373937,
  0.1722084, 0.2026768, 0.2189366, 0.4132893, 0.2233801, -0.06366426, 
    -0.3198164, -0.5716393, -0.5695727, -0.3674567, -0.2115159, -0.3761477, 
    -0.1205654, -0.2155522, 0.065063, 0.2456293, 0.0856359, 0.2625563, 
    0.3482987, 0.3496822, 0.2364496, 1.208553, 1.770271, 0.3119855, 
    -0.6998634, -0.4193441, -0.1408777, -0.01875842, 0.08854949, 0.5473713, 
    0.5454831, 0.2762936, 0.2411371, -0.3458905, -1.364364, -1.533635, 
    -1.136141, -0.829452, -0.6142014, -0.3478765, -0.3223883, -0.3411546, 
    -0.3453864, -0.2276291, -0.09375858, -0.09842968, -0.2145915, -0.3118083, 
    -0.3038985, -0.3644772, -0.3847413, -0.5168054, -0.5225182, -0.4191487, 
    -0.2098551, -0.2427491, -0.3080971, -0.1955328, -0.1700933, -0.08173108, 
    -0.1899338, -0.249439, -0.3619885, -0.3044362, -0.3427334, -0.2355723, 
    -0.06112576, -0.1747971, 0.2136469, 0.2392329, 0.02160603, 0.005102515, 
    0.337475, 0.6237869, 0.1595616, -0.1432704, -0.4380947, -0.6942959, 
    -0.8293707, -0.8729904, -0.8304613, -0.8094162, -0.5520756, -0.3255781, 
    -0.11674, -0.03366756, -0.007512093, -0.00481081, -0.06239557, 
    -0.1133552, -0.1901798, -0.2761173, -0.4432049, -0.3240485, 0.1421139, 
    0.2975671,
  0.1170492, 0.0335362, -0.08440002, 0.01380974, -0.2002853, -0.6391199, 
    -0.5510665, -0.6083744, -0.9789801, -0.8018641, -0.3879158, -0.4452881, 
    -0.4386154, -0.3653893, 0.2070228, 0.246443, 0.1211019, 0.2782627, 
    0.3670648, 0.4181069, 0.1823156, 0.6394444, 1.124747, 0.7477448, 
    0.1683669, 0.07264817, -0.05007386, 0.02176881, 0.3831618, 0.3979082, 
    0.3904862, 0.5769122, 0.4813226, 0.3864334, -0.3087161, -0.9801517, 
    -0.9951257, -0.749862, -0.7517663, -0.6797445, -0.403931, -0.220549, 
    -0.2342372, -0.07007709, -0.0126064, -0.0355556, -0.08840394, -0.2472743, 
    -0.4069584, -0.6157146, -0.6186445, -0.6636149, -0.7922605, -0.9045981, 
    -0.6853762, -0.4783124, -0.5335859, -0.4634197, -0.3239174, -0.2239671, 
    -0.1825123, -0.1450446, -0.2577891, -0.2709565, -0.4275804, -0.3124437, 
    0.1293695, -0.01145065, -0.01016499, -0.0120855, -0.1262293, 0.1617752, 
    0.9973875, 1.15424, 0.4530511, 0.1281489, -0.3129481, -0.564901, 
    -0.7232832, -0.9859624, -1.036972, -0.9673426, -0.6643317, -0.397014, 
    -0.1253827, 0.0383873, 0.07281089, 0.06301188, -0.1020269, -0.2606864, 
    -0.4187598, -0.369379, -0.1696057, -0.2679615, -0.1872311, 0.06677246,
  -0.1053308, -0.08620644, -0.176913, -0.1142828, -0.06991434, -0.5455818, 
    -0.537297, -0.4887619, -1.093254, -1.007788, -0.4036869, -0.4464442, 
    -0.7853436, -0.5996504, 0.02173638, 0.05174907, 0.001749071, 0.1975013, 
    0.2896888, 0.2361731, 0.3077064, 0.6408443, 0.6430739, 0.1845292, 
    -0.2379806, -0.04885292, -0.1345623, -0.3578539, 0.09618306, 0.6526931, 
    0.6861081, 0.598885, 0.5659581, 0.6098223, 0.5120193, -0.007251382, 
    -0.3906336, -0.5480553, -0.6334229, -0.7911866, -0.6750406, -0.3726481, 
    -0.2092853, -0.0357995, 0.002514482, 0.08405733, 0.03612411, -0.1475185, 
    -0.2501064, -0.5467373, -0.7272874, -0.7823328, -0.8678635, -1.024878, 
    -1.023511, -0.8279871, -0.7893316, -0.7165121, -0.5435306, -0.4154215, 
    -0.2354579, -0.1392341, -0.2574964, -0.3319917, -0.4141035, -0.1613858, 
    0.08905387, 0.02652121, -0.1927822, -0.2913498, -0.1294355, 0.4868891, 
    1.237963, 0.9504634, 0.6701248, 0.7465575, 0.1317298, -0.5663661, 
    -0.7311283, -0.794084, -1.041154, -1.170841, -0.9880294, -0.7282964, 
    -0.3350022, -0.0688237, 0.05546033, 0.05993652, -0.1225512, -0.2691169, 
    -0.5679288, -0.9079685, -0.5896888, -0.2906828, 0.0005941391, 0.08063905,
  0.2557533, 0.3428786, 0.1465082, -0.1342697, -0.3559656, -0.6177981, 
    -0.537378, -0.5284427, -0.967684, -0.8819903, -0.3657146, -0.3736576, 
    -0.5969651, -0.3557217, -0.009709284, -0.09986225, -0.3916264, 
    -0.3916425, 0.1672282, 0.4550861, 0.3354082, 0.154272, 0.0114007, 
    -0.1347255, -0.7044843, -0.7218022, -0.3553141, -0.4115313, -0.08653216, 
    0.5088135, 0.6751055, 0.6187739, 0.5613846, 0.4481684, 0.5570226, 
    0.5310785, 0.163045, -0.1468017, -0.1264899, -0.4129803, -0.6204674, 
    -0.4911866, -0.4095135, -0.2702229, -0.1205971, 0.04771328, 0.1325276, 
    0.02399909, -0.1498942, -0.3854085, -0.5263105, -0.7825606, -1.076132, 
    -1.166659, -1.229533, -1.165145, -0.9667567, -0.8334234, -0.8341884, 
    -0.8429609, -0.7250082, -0.493938, -0.3974857, -0.4667082, -0.152369, 
    0.1579665, 0.1390863, 0.06136823, 0.1275473, 0.245044, 0.05749512, 
    0.1193435, 0.476766, 0.4187415, 0.5646074, 1.132788, 0.9411702, 
    0.08254409, -0.4303629, -0.697665, -0.9370689, -1.010555, -0.9232504, 
    -0.813957, -0.5367105, -0.3159589, -0.14218, -0.000317812, -0.1402427, 
    -0.3643315, -0.6295173, -0.9790132, -1.206666, -1.10429, -0.4546638, 
    0.1556718,
  -0.2773844, -0.2006429, -0.1455, -0.2010828, -0.5890874, -0.8658615, 
    -0.5292079, -0.3513597, -0.5669521, -0.567652, -0.4635665, -0.2294192, 
    -0.1535732, -0.3124435, -0.3925706, -0.3649012, -0.4572515, -0.7533453, 
    -0.4319421, 0.07901156, -0.003914595, -0.2457275, 0.1026448, 0.4549718, 
    0.3957107, 0.3424228, 0.2317946, -0.1000576, 0.02910911, 0.2876704, 
    0.4445228, 0.5044186, 0.4490961, 0.298624, 0.5456129, 0.7274327, 
    0.5407304, 0.2725664, 0.4789143, 0.4688884, 0.1899812, 0.182169, 
    0.2246819, 0.2749422, 0.2924554, 0.2888746, 0.3599358, 0.3687901, 
    0.1357985, -0.1250246, -0.2239828, -0.4551191, -0.8076416, -1.043303, 
    -1.198397, -1.236938, -1.05647, -0.858846, -0.8193283, -0.8251553, 
    -0.8743088, -0.8114994, -0.6608324, -0.4685144, -0.1005127, 0.379988, 
    0.300919, 0.1416743, 0.3415607, 0.7114499, 0.5674231, 0.2208743, 
    0.2621822, 0.3596596, 0.3558512, 0.6915935, 0.9743246, 0.8617431, 
    0.329761, -0.3513589, -0.7445078, -0.7350183, -0.5882087, -0.4704838, 
    -0.36622, -0.3007243, -0.1658772, -0.05345911, -0.009090773, -0.1957118, 
    -0.599862, -0.9222577, -1.217261, -1.482041, -1.03772, -0.4646893,
  -0.5281826, -0.4940513, -0.2664306, -0.06988174, -0.3791917, -0.834335, 
    -0.7282311, -0.5068601, -0.4821051, -0.5347744, -0.4881272, -0.2770595, 
    -0.1619385, -0.3236091, -0.4782639, -0.5027917, -0.3788663, -0.623251, 
    -0.6626878, -0.2090582, 0.02036893, -0.000741154, 0.2286536, 0.2106685, 
    0.2457922, 0.5309486, 0.4639075, 0.1214593, 0.07679793, 0.08740985, 
    0.2927972, 0.4265539, 0.346557, 0.1194248, 0.04538514, 0.2655674, 
    0.4678462, 0.3777421, 0.4703367, 0.701896, 0.6168702, 0.5532472, 
    0.6470616, 0.8298905, 1.039396, 1.115226, 1.024438, 0.8869054, 0.7747636, 
    0.530997, 0.284936, 0.0360589, -0.2933187, -0.5855227, -0.8849692, 
    -1.090129, -1.007544, -0.8243247, -0.7685955, -0.7836185, -0.8379644, 
    -0.8900311, -0.7167728, -0.3952556, -0.2007731, -0.0817796, 0.007071331, 
    0.01468867, 0.08376426, 0.4687251, 0.8185787, 0.6927487, 0.54672, 
    0.5402914, 0.4273189, 0.3748124, 0.535164, 0.7279214, 0.7243896, 
    0.3539473, -0.1356366, -0.4423919, -0.3652921, -0.05422425, 0.1596918, 
    0.1867588, 0.2036858, 0.09291196, 0.1388429, 0.1253818, -0.2731858, 
    -0.7118735, -0.9996989, -1.058944, -1.018645, -0.6491135,
  0.06538832, -0.229598, -0.2945235, -0.1127201, -0.1340418, -0.2912034, 
    -0.4780198, -0.3838628, -0.1882249, -0.1901943, -0.2218512, -0.2172939, 
    -0.2067633, -0.08684143, -0.1179937, 0.0007888675, -0.005558729, 
    -0.2236089, -0.2719977, 0.08723092, 0.2772211, 0.3527584, 0.2367753, 
    0.1298578, 0.1285394, 0.2202549, 0.1575433, 0.04919374, 0.1636469, 
    0.2216221, 0.3265863, 0.4648351, 0.5222244, 0.4653396, 0.2339268, 
    0.197029, 0.3330479, 0.3616286, 0.363289, 0.4419673, 0.487166, 0.4835366, 
    0.5628824, 0.7430906, 1.049666, 1.399959, 1.613566, 1.565584, 1.356225, 
    1.119295, 0.9679928, 0.7377031, 0.3397696, 0.03628683, -0.2517664, 
    -0.6267176, -0.7924891, -0.6493411, -0.587378, -0.5333092, -0.4116615, 
    -0.4168544, -0.386288, -0.2019781, -0.09732318, -0.07824749, 0.004988, 
    0.01836693, -0.07806863, 0.1277094, 0.5474033, 0.7781814, 0.8452063, 
    0.8355708, 0.6736242, 0.5559646, 0.4913976, 0.4276119, 0.4023842, 
    0.3306231, 0.09839678, -0.1430256, -0.1797934, 0.07282662, 0.4017653, 
    0.7287023, 1.010473, 0.8930905, 0.6334066, 0.4721271, 0.3126215, 
    -0.1236253, -0.7167078, -0.8468673, -0.5283615, -0.0575771,
  0.3665928, 0.1812903, -0.1200283, -0.12343, 0.05287211, 0.04434365, 
    -0.1948816, -0.1302496, 0.06206822, 0.05825949, -0.01346904, 0.06577902, 
    0.1046299, 0.1032301, 0.2309809, 0.471134, 0.5670977, 0.3601319, 
    0.1640378, 0.3709385, 0.6917068, 0.6278884, 0.3342199, 0.1386966, 
    0.04911292, 0.07723749, 0.03729594, -0.04156131, -0.01343608, 0.1218339, 
    0.2614008, 0.1891356, 0.1513913, 0.258764, 0.2788975, 0.299682, 
    0.3311762, 0.2799067, 0.1634029, 0.261531, 0.5551996, 0.7220779, 
    0.8332272, 0.9883379, 1.167781, 1.335229, 1.634904, 1.933813, 1.958666, 
    1.70411, 1.483716, 1.238029, 0.9120843, 0.6083896, 0.321964, -0.1560962, 
    -0.4408779, -0.459986, -0.4049077, -0.2856369, -0.09133339, -0.03435051, 
    -0.04455566, -0.02855682, 0.06371212, 0.1640375, 0.1847894, 0.1023676, 
    -0.02416241, 0.09787554, 0.2789463, 0.4419509, 0.6464919, 0.5697992, 
    0.444376, 0.337475, 0.431111, 0.4239821, 0.2042231, 0.0194577, 
    -0.1470464, -0.3038656, -0.3639572, -0.208374, 0.06237745, 0.4325597, 
    0.8922603, 1.212247, 1.170304, 0.9334224, 0.7868241, 0.4945551, 
    -0.01490134, -0.315894, -0.0824793, 0.2399978,
  0.4660887, 0.571557, 0.2541254, -0.08168191, -0.09460509, -0.02650613, 
    -0.04165913, 0.08431751, 0.2491289, 0.1687577, -0.03633687, -0.06053934, 
    0.05637147, 0.2096104, 0.3266514, 0.4183182, 0.4183019, 0.3726151, 
    0.2959385, 0.2753985, 0.4215734, 0.5959058, 0.6685138, 0.5284095, 
    0.4533442, 0.4219639, 0.4674066, 0.2920161, 0.102335, 0.1169673, 
    0.254809, 0.1555254, -0.003979445, -0.03215349, 0.06747186, 0.1886468, 
    0.2653558, 0.1410233, -0.1527425, -0.1868411, 0.1284745, 0.3888588, 
    0.5380121, 0.8506912, 1.336596, 1.556583, 1.554077, 1.721736, 1.92102, 
    1.900366, 1.759269, 1.531665, 1.229728, 0.9514725, 0.6942623, 0.3806229, 
    0.01009846, -0.1441329, -0.04423046, 0.1318274, 0.2490962, 0.2700932, 
    0.1943438, 0.2246985, 0.2089596, 0.05935019, -0.07645731, -0.1792731, 
    -0.1356533, 0.006176174, 0.06626725, 0.07803489, 0.1586501, 0.2091872, 
    0.11866, 0.009040743, 0.09777769, 0.1908278, 0.1792393, 0.04195088, 
    -0.05524951, -0.3416917, -0.5172774, -0.5548098, -0.3983967, -0.07551265, 
    0.4636312, 0.9679607, 1.122388, 1.026505, 0.8795328, 0.6530513, 
    0.3376215, 0.03718203, -0.04816937, 0.09020942,
  0.3520421, 0.3257888, 0.2980544, 0.1522862, 0.003392965, -0.156275, 
    -0.234107, -0.07670145, 0.117781, 0.1006423, -0.1009365, -0.2630458, 
    -0.2396734, -0.03156799, 0.1745518, 0.2203363, 0.06143332, -0.01524311, 
    0.07648866, 0.1869215, 0.2110103, 0.2643142, 0.4051995, 0.4621172, 
    0.478035, 0.4346105, 0.3760492, 0.3810297, 0.352693, 0.3052812, 
    0.2468991, 0.2328529, 0.1753008, 0.1239499, 0.001114607, -0.006877065, 
    0.05479276, -0.1521889, -0.6232991, -0.7801187, -0.6452554, -0.3801678, 
    -0.1671307, -0.009562373, 0.4667722, 0.9989662, 1.212866, 1.284155, 
    1.324487, 1.377123, 1.412638, 1.343042, 1.09729, 0.8539469, 0.7340251, 
    0.6166906, 0.3975496, 0.2133701, 0.2935786, 0.483357, 0.5016351, 
    0.4654381, 0.4339272, 0.1696041, 0.01416773, -0.1286056, -0.2105394, 
    -0.2796637, -0.2652431, -0.1826259, -0.07567605, -0.02175349, 0.06809026, 
    0.1703855, 0.1775469, 0.05856878, -0.02243713, 0.08900492, 0.199861, 
    0.3075923, 0.2898678, 0.128377, -0.3885666, -0.6831468, -0.7029709, 
    -0.4001387, 0.1613686, 0.7114011, 1.05782, 1.101863, 0.9703526, 
    0.7533118, 0.5653236, 0.4273677, 0.3361567, 0.3386793,
  0.1706294, 0.1452875, 0.201391, 0.2430739, -0.01561747, -0.4501064, 
    -0.5041102, -0.2886643, -0.07486226, -0.1070563, -0.2300055, -0.2993252, 
    -0.3520107, -0.3486416, -0.154859, 0.06784607, 0.09240663, -0.0395107, 
    -0.1246832, 0.01475364, 0.1666091, 0.175154, 0.07788855, 0.004353642, 
    -0.004402995, 0.008943439, 0.03306448, 0.08505011, 0.1350173, 0.1357986, 
    0.03763774, 0.01047307, 0.1876541, 0.3408606, 0.2328363, 0.02696067, 
    -0.1306891, -0.2970626, -0.6116129, -0.9048746, -0.9310961, -0.6946045, 
    -0.5450603, -0.4212807, -0.3159266, -0.03643441, 0.2986732, 0.5294354, 
    0.6528236, 0.6624594, 0.7578694, 0.7525307, 0.6846429, 0.5700434, 
    0.6145586, 0.6633544, 0.7239013, 0.6370686, 0.5725017, 0.5259358, 
    0.6316977, 0.6699297, 0.4018145, 0.2786213, 0.1434971, 0.1286696, 
    0.1660232, 0.1646885, 0.1062738, 0.06693462, 0.1568435, 0.3240801, 
    0.3939857, 0.4018959, 0.3282794, 0.1514725, 0.001911938, 0.05952901, 
    0.2690346, 0.5216875, 0.6407142, 0.3739662, 0.01091278, -0.2658451, 
    -0.3538336, -0.210409, 0.08762147, 0.444555, 0.7583082, 0.9526607, 
    0.9424717, 0.6916091, 0.417781, 0.311173, 0.3337966, 0.2731685,
  0.2785395, 0.3238195, 0.3798252, 0.189184, -0.1888433, -0.5361741, 
    -0.4782639, -0.2785569, -0.1691168, -0.2611578, -0.334693, -0.325139, 
    -0.309107, -0.3209234, -0.2802334, -0.09680236, 0.06450947, 0.07396585, 
    0.02346134, 0.08550555, 0.2396399, 0.2980057, 0.1865472, 0.05529726, 
    0.0141353, 0.02163851, 0.01493269, 0.02624458, 0.06086367, 0.07320088, 
    0.0229242, 0.0217686, 0.120613, 0.2895094, 0.3174555, 0.1420323, 
    -0.06981669, -0.1652106, -0.326083, -0.5405846, -0.7242923, -0.8463953, 
    -0.7121176, -0.525578, -0.4611409, -0.4166753, -0.3280692, -0.7145276, 
    -0.497226, -0.3264897, -0.1970627, -0.1733643, 0.2301673, 0.2744704, 
    0.2771397, 0.3151443, 0.3467197, 0.338289, 0.2763753, 0.2588623, 
    0.3664629, 0.3824137, 0.3812419, 0.2632239, 0.1966221, 0.2434971, 
    0.3235915, 0.3492588, 0.334708, 0.3606033, 0.4767493, 0.5300372, 
    0.5964597, 0.4517822, 0.2308836, 0.04631317, -0.2176194, -0.141122, 
    0.185522, 0.5330157, 0.6835039, 0.4482662, 0.1054437, -0.1429938, 
    -0.1069747, 0.1598228, 0.2510822, 0.2585531, 0.3895909, 0.5682367, 
    0.6566482, 0.5362868, 0.3152582, 0.2548741, 0.2485102, 0.2874424,
  0.4799066, 0.5535883, 0.5192621, 0.422615, 0.1061763, -0.1612555, 
    -0.1899339, -0.2637132, -0.2672451, -0.3253017, -0.3250413, -0.3504969, 
    -0.3398199, -0.3677495, -0.4032476, -0.3387132, -0.1878018, -0.04460478, 
    0.0802325, 0.273999, 0.3675209, 0.3843828, 0.2932694, 0.1521397, 
    0.05401143, -0.01493385, -0.07592019, -0.1433681, -0.1601162, -0.1655361, 
    -0.2096765, -0.1411381, -0.03381401, 0.03994894, -0.001001582, 
    -0.1117763, -0.1643805, -0.2185634, -0.2215908, -0.2442796, -0.3958909, 
    -0.5571213, -0.6335862, -0.5765713, -0.4890063, -0.4440839, -0.409302, 
    -0.4060147, -0.4001069, -0.3651128, -0.3506436, -0.2216558, -0.02954912, 
    0.2067622, 0.3275954, 0.3480544, 0.3042556, 0.3003494, 0.3942296, 
    0.466837, 0.5127518, 0.5730706, 0.5659744, 0.5327061, 0.4205479, 
    0.2967686, 0.2449294, 0.2351312, 0.3218663, 0.4486567, 0.5203204, 
    0.5428137, 0.4871334, 0.3155841, 0.1434813, 0.01556778, -0.06696832, 
    -0.1045334, 0.06646264, 0.4045976, 0.6065182, 0.4953038, 0.162182, 
    -0.1777592, -0.281568, -0.2568607, -0.1527264, 0.06273508, 0.0945549, 
    0.2047114, 0.3028402, 0.396199, 0.3834062, 0.3677324, 0.3746171, 0.38907,
  0.7065181, 0.6504471, 0.5928299, 0.4822667, 0.3701247, 0.3338292, 
    0.2607009, 0.1597243, 0.0630772, -0.05878153, -0.235523, -0.3415775, 
    -0.3796961, -0.4518315, -0.4984948, -0.42286, -0.2946863, -0.1237872, 
    0.09227669, 0.2968993, 0.4396076, 0.4680911, 0.4106523, 0.2969151, 
    0.1891351, 0.08360127, 0.0006748736, -0.09219623, -0.1117926, -0.161581, 
    -0.1511642, -0.0586344, -0.009724855, 0.01931095, -0.02624571, 
    -0.1084235, -0.2025804, -0.1832933, -0.1328375, -0.04652567, -0.02655496, 
    -0.03096578, -0.1195726, -0.1718349, -0.2602301, -0.3146246, -0.392294, 
    -0.475106, -0.5310147, -0.3909595, -0.3292408, -0.2038178, 0.0448482, 
    0.2130613, 0.3785563, 0.4383379, 0.3894613, 0.3106852, 0.1719486, 
    0.3013591, 0.3638099, 0.4661209, 0.5621822, 0.5725336, 0.459057, 
    0.2584548, 0.1064203, 0.06265402, 0.132348, 0.2683507, 0.2739661, 
    0.2894123, 0.2278562, 0.1607827, 0.0009520054, -0.003605366, -0.1233971, 
    -0.1017175, -8.583069e-006, 0.1307042, 0.3047927, 0.2541583, 0.1655517, 
    -0.009317994, -0.09652507, -0.1808354, -0.20398, -0.2387128, -0.2966719, 
    -0.2129481, -0.1142988, 0.1323321, 0.1894778, 0.4847088, 0.7845947, 
    0.7692949,
  0.9016032, 0.8493244, 0.7731038, 0.7167232, 0.663712, 0.6358638, 0.5883052, 
    0.4606846, 0.2299554, 0.01284951, -0.2040125, -0.4043542, -0.5399174, 
    -0.5374923, -0.4983483, -0.5330815, -0.252287, -0.05054545, 0.1938723, 
    0.3675537, 0.4804608, 0.5152584, 0.4940507, 0.421736, 0.309236, 
    0.2055089, 0.1629469, 0.1732985, 0.1880935, 0.2174066, 0.2120032, 
    0.1825433, 0.08796328, 0.001179457, -0.08796448, -0.04226134, 
    -0.03939676, -0.02837788, 0.02440532, 0.06992941, 0.1235752, 0.1356032, 
    0.09857523, 0.02865337, -0.05332905, -0.1582444, -0.2683193, -0.3633714, 
    -0.4049399, -0.3978275, -0.3732179, -0.2989013, -0.1578207, -0.02108586, 
    0.07867014, 0.1539307, 0.2302327, 0.2856039, 0.3285726, 0.3754964, 
    0.4084555, 0.4288, 0.4236567, 0.5398188, 0.4959874, 0.4238519, 0.3406325, 
    0.2418371, 0.179386, 0.2113847, 0.09237421, 0.04095829, 0.03272259, 
    -0.06957221, -0.1068443, -0.09211457, -0.01856315, 0.08426905, 0.11171, 
    0.09696394, 0.04112081, -0.01420122, -0.08809435, -0.06485188, 
    0.004435301, 0.01262212, -0.03705287, -0.08290261, -0.2000574, 
    -0.3703698, -0.5020102, -0.2106528, 0.09367704, 0.4000407, 0.4333253, 
    0.7214435,
  0.3653075, 0.5226969, 0.7103918, 0.7079667, 0.638061, 0.4922439, 0.4148026, 
    0.3123938, 0.2215248, 0.08713353, -0.1180584, -0.2650635, -0.4320557, 
    -0.535311, -0.590145, -0.575464, -0.4757081, -0.3528402, -0.1657797, 
    0.02928865, 0.1955645, 0.3126218, 0.3782305, 0.402742, 0.390193, 
    0.3999913, 0.3927973, 0.3798741, 0.3706456, 0.3327224, 0.2558669, 
    0.1730219, 0.08750755, 0.02224059, -0.02481343, -0.06244364, -0.0833258, 
    -0.0892503, -0.1130621, -0.1434169, -0.1511806, -0.1661383, -0.1713629, 
    -0.1763597, -0.1936122, -0.2278408, -0.2831305, -0.3364671, -0.3562424, 
    -0.3677497, -0.3619066, -0.3333258, -0.3231043, -0.3126062, -0.2909266, 
    -0.2444096, -0.1680098, -0.06748903, 0.0390867, 0.1607664, 0.2771401, 
    0.3699622, 0.4418534, 0.4906816, 0.4834386, 0.5230385, 0.4904701, 
    0.4351315, 0.3242917, 0.2170162, 0.09789193, 0.01182407, -0.03438359, 
    -0.07069546, -0.05564022, 0.03719848, 0.02336365, -0.01257384, 
    -0.03702046, -0.07635966, -0.1337326, -0.1907308, -0.2088623, -0.1515867, 
    -0.04523945, 0.05469519, 0.1242588, 0.16796, 0.1582108, 0.1112058, 
    0.0696367, 0.03405738, 0.123836, 0.2089922, 0.3159747, 0.3468828,
  0.2565669, 0.2487707, 0.2738031, 0.3028397, 0.2857334, 0.2659418, 
    0.2286859, 0.1752843, 0.1196203, 0.02622837, -0.08142132, -0.1827071, 
    -0.2836348, -0.3731856, -0.4620199, -0.5081626, -0.5082277, -0.4639731, 
    -0.3854089, -0.2939213, -0.1788334, -0.0463953, 0.09431112, 0.214005, 
    0.2822829, 0.3382074, 0.3857172, 0.4005121, 0.3870192, 0.3658929, 
    0.3286696, 0.2656651, 0.19532, 0.1318923, 0.07062927, 0.01166117, 
    -0.05231991, -0.1091232, -0.1618413, -0.2140061, -0.247079, -0.2909917, 
    -0.3245203, -0.3564539, -0.3840907, -0.4028246, -0.4182054, -0.4207281, 
    -0.4142503, -0.4086188, -0.3871018, -0.3612718, -0.3268154, -0.3024013, 
    -0.2845302, -0.2533778, -0.2019457, -0.1474044, -0.06817263, 0.02417761, 
    0.1328365, 0.2217851, 0.3161535, 0.3826085, 0.4350501, 0.4590573, 
    0.4420325, 0.3786212, 0.3045651, 0.2266517, 0.1181881, 0.1118728, 
    0.04050249, -0.006812125, -0.03920145, -0.06711486, -0.09501183, 
    -0.1261479, -0.1611249, -0.1830325, -0.1846601, -0.1775962, -0.1350179, 
    -0.05489123, 0.04790795, 0.1434808, 0.2220127, 0.2859125, 0.345369, 
    0.37963, 0.3779048, 0.3538164, 0.3464597, 0.3153725, 0.2787025, 0.2653561,
  0.2688715, 0.265242, 0.2551671, 0.2223709, 0.1994706, 0.15852, 0.1127355, 
    0.05663204, -0.003849745, -0.06483603, -0.1241297, -0.1898686, 
    -0.2340743, -0.2807866, -0.3208256, -0.3378504, -0.3393966, -0.3139734, 
    -0.2724532, -0.2169031, -0.1587, -0.09663954, -0.03081927, 0.03024843, 
    0.08571716, 0.1247797, 0.1652419, 0.1975336, 0.2064691, 0.2127679, 
    0.2261794, 0.2216547, 0.2038649, 0.174275, 0.1612218, 0.1500564, 
    0.1277419, 0.08736122, 0.04738724, -0.007251561, -0.06016487, -0.1189865, 
    -0.1773849, -0.2302658, -0.2845464, -0.3348394, -0.3744065, -0.4009201, 
    -0.4297125, -0.4413499, -0.4472093, -0.4332119, -0.4110764, -0.3794847, 
    -0.3353115, -0.2766852, -0.2253506, -0.1659267, -0.1094326, -0.03073788, 
    0.05358845, 0.1162511, 0.1671464, 0.2097735, 0.2524329, 0.2726315, 
    0.2778724, 0.2681719, 0.2435789, 0.2033281, 0.150317, 0.1026443, 
    0.05521601, 0.00295347, -0.04620016, -0.08160053, -0.1119391, -0.1206957, 
    -0.1244716, -0.1269943, -0.1175704, -0.1033777, -0.07191634, -0.04120341, 
    0.001277059, 0.05537863, 0.09811951, 0.1340245, 0.1835036, 0.2206618, 
    0.2444412, 0.2605057, 0.2634354, 0.2734614, 0.2711503, 0.2701085,
  0.2229567, 0.2047927, 0.19685, 0.1792718, 0.1656488, 0.150333, 0.1329828, 
    0.123445, 0.1036859, 0.08680767, 0.06201926, 0.04465273, 0.02103618, 
    0.00231871, -0.007918894, -0.01247618, -0.01774962, -0.02126525, 
    -0.02126525, -0.01818909, -0.01548725, -0.008879185, -0.002157179, 
    0.004190477, 0.01820415, 0.02775819, 0.03716573, 0.04239035, 0.04642682, 
    0.05375102, 0.05659935, 0.05589944, 0.05778748, 0.05432069, 0.04598731, 
    0.04086035, 0.03086686, 0.007120073, -0.01052302, -0.02634335, 
    -0.04668838, -0.06278539, -0.0775314, -0.09292859, -0.1174728, 
    -0.1451095, -0.1641851, -0.1762457, -0.1890387, -0.2034918, -0.2103603, 
    -0.2132086, -0.2122809, -0.2033453, -0.1865484, -0.1653733, -0.1451097, 
    -0.1205817, -0.1032802, -0.07670146, -0.04496318, -0.01807514, 
    0.01146591, 0.03374785, 0.05350709, 0.0720129, 0.08169717, 0.08970499, 
    0.1020097, 0.1182205, 0.122322, 0.1290602, 0.1361078, 0.129988, 
    0.1256586, 0.1226638, 0.1225498, 0.1252842, 0.1288975, 0.1303624, 
    0.1270258, 0.1259678, 0.1333083, 0.1409581, 0.1477777, 0.155281, 
    0.1567946, 0.1686762, 0.1829991, 0.1923903, 0.2001866, 0.2131098, 
    0.2212315, 0.2221266, 0.2233473, 0.2255121,
  0.5780702, 0.6049261, 0.6249294, 0.6372995, 0.6423612, 0.6392851, 
    0.6287055, 0.6111441, 0.5866323, 0.5567493, 0.522944, 0.4875922, 0.45154, 
    0.4157166, 0.3797631, 0.3443954, 0.3091416, 0.2731547, 0.2352486, 
    0.1937933, 0.1483181, 0.09851342, 0.04385839, -0.01530501, -0.07957888, 
    -0.1475313, -0.2194066, -0.2939188, -0.3705952, -0.4483783, -0.5241265, 
    -0.5963926, -0.662961, -0.7222385, -0.7748265, -0.8184137, -0.8526416, 
    -0.8776584, -0.8930717, -0.8998752, -0.8993382, -0.8929424, -0.8821344, 
    -0.8676977, -0.8510313, -0.8336964, -0.8107805, -0.7938366, -0.7741103, 
    -0.7419324, -0.7160378, -0.6696177, -0.6650929, -0.6857147, -0.6196995, 
    -0.6332579, -0.6162653, -0.5746965, -0.4893126, -0.4327536, -0.4511456, 
    -0.4052308, -0.3710835, -0.3062396, -0.2473688, -0.187001, -0.1196833, 
    -0.04972887, 0.02103925, 0.07977962, 0.1372831, 0.1866155, 0.2280049, 
    0.3287866, 0.249929, 0.2678652, 0.2675238, 0.3385034, 0.2829533, 
    0.2761173, 0.2638454, 0.2524521, 0.2419214, 0.2351019, 0.232156, 
    0.2354766, 0.2452419, 0.2620062, 0.285167, 0.3145778, 0.3495553, 
    0.3885193, 0.4288843, 0.4697371, 0.5089951, 0.5453396,
  0.1844025, 0.2417431, 0.2982206, 0.3421826, 0.3728623, 0.389122, 0.3881946, 
    0.3712997, 0.3426864, 0.3065863, 0.2656031, 0.2259548, 0.191921, 
    0.1654561, 0.1506286, 0.1479437, 0.1538357, 0.163878, 0.1796006, 
    0.1961373, 0.2069607, 0.2067165, 0.1913031, 0.1546331, 0.09630013, 
    0.01627064, -0.08368039, -0.198411, -0.3203676, -0.4413958, -0.5533423, 
    -0.6463428, -0.7148819, -0.7553596, -0.7674212, -0.7538791, -0.7155485, 
    -0.6549864, -0.5758848, -0.4887438, -0.4134989, -0.2867575, -0.1509981, 
    -0.1060925, -0.0676651, -0.02816296, -0.0510149, -0.05820799, 
    -0.08480358, -0.1118383, -0.1567926, -0.2018285, -0.2080622, -0.2344947, 
    -0.2376519, -0.2097063, -0.2016168, -0.1844944, -0.1630264, -0.1338758, 
    -0.1111057, -0.07658434, -0.02228808, 0.03342485, 0.07746792, 0.1396587, 
    0.1724555, 0.1992786, 0.2460882, 0.3095648, 0.4024522, 0.488585, 
    0.5645616, 0.6336043, 0.6199813, 0.5734811, 0.5591903, 0.5160756, 
    0.5514917, 0.2979107, 0.2685814, 0.2377706, 0.06934667, 0.05186617, 
    -0.02218968, -0.07580306, -0.112017, -0.13399, -0.1403382, -0.1298397, 
    -0.1032286, -0.06550074, -0.02603006, 0.02411604, 0.08034945, 0.1351838,
  -0.1019912, -0.06196833, -0.008111238, 0.05790424, 0.1291606, 0.1883084, 
    0.2276474, 0.2736436, 0.332221, 0.3942004, 0.467833, 0.5315211, 
    0.5742946, 0.6021914, 0.6213818, 0.6371207, 0.6442981, 0.6296, 0.5940211, 
    0.5464139, 0.4909777, 0.4228786, 0.332921, 0.2321396, 0.1393011, 
    0.07763118, 0.02362764, -0.07039928, -0.216363, -0.3808653, -0.5343323, 
    -0.6523492, -0.7212296, -0.7462456, -0.7335341, -0.6902237, -0.6110725, 
    -0.5125542, -0.4031959, -0.293056, -0.2087622, -0.05109549, 0.01436663, 
    0.1186466, 0.1178486, 0.1771429, 0.1968045, 0.2313097, 0.2705187, 
    0.2903917, 0.2830511, 0.2592393, 0.2197701, 0.174783, 0.1444281, 
    0.1184028, 0.07336688, 0.0425396, 0.02450609, 0.0208931, 0.0362258, 
    0.06046057, 0.1077266, 0.1808386, 0.2497988, 0.3074486, 0.352598, 
    0.3881294, 0.4375596, 0.477778, 0.5054793, 0.5117292, 0.4990344, 
    0.4599071, 0.4211864, 0.3713646, 0.3528757, 0.533051, 0.4279079, 
    0.3591578, 0.3118923, 0.2790146, 0.1611764, 0.1246365, 0.08243262, 
    0.04029387, -0.006336689, -0.03517795, -0.07686114, -0.1555727, 
    -0.1278212, -0.1360245, -0.1187224, -0.1134009, -0.1124077, -0.1168995,
  -0.2373101, -0.254335, -0.2160537, -0.1478896, -0.07269436, -0.01709509, 
    0.008490562, 0.00344491, -0.002837658, 0.01809359, 0.07125139, 0.1516552, 
    0.2317657, 0.2873492, 0.3286896, 0.374474, 0.3311305, 0.2737901, 
    0.2581325, 0.2168239, 0.1498318, 0.08091879, -0.01795816, -0.12551, 
    -0.1899471, -0.1747776, -0.128163, -0.1535536, -0.2376847, -0.3201396, 
    -0.3675672, -0.3938531, -0.4226454, -0.4645562, -0.5032607, -0.5098363, 
    -0.4810113, -0.4197652, -0.3569555, -0.31511, -0.2851934, -0.2036834, 
    -0.1042042, 0.0355258, 0.2061954, 0.449506, 0.3838649, 0.454747, 
    0.4587996, 0.4180607, 0.3214298, 0.2128689, 0.1287868, 0.027192, 
    -0.02383363, -0.003342122, -0.04106987, 0.03956151, 0.0635525, 
    0.07374132, 0.03941512, 0.008132696, 0.01934671, 0.09472104, 0.2018501, 
    0.2851182, 0.3405054, 0.3944278, 0.4375596, 0.4536886, 0.4579697, 
    0.4306583, 0.3444285, 0.2517357, 0.1949978, 0.1626897, 0.09782958, 
    0.05881548, 0.0368433, 0.06099701, 0.1159775, 0.1336045, 0.1218696, 
    0.08113086, 0.04180771, 0.01412208, -0.00588116, -0.01585829, 
    -0.03153217, -0.03713119, 0.06290126, 0.09688568, 0.08710313, 0.04439545, 
    -0.06095934, -0.1683811,
  -0.1594617, -0.1465549, -0.06610203, 0.03830862, 0.08436918, 0.05866957, 
    0.008881569, -0.04526901, 0.08080292, 0.05053043, 0.1774683, 0.263732, 
    0.3056421, 0.368484, 0.5414009, 0.7507272, 0.8170519, 0.7540145, 
    0.6484003, 0.3307073, 0.189236, 0.0739367, -0.06548429, -0.1985731, 
    -0.2797256, -0.2769425, -0.3658423, -0.519537, -0.6156306, -0.6169648, 
    -0.5892797, -0.598948, -0.6210668, -0.668772, -0.7410383, -0.7570534, 
    -0.6606665, -0.4832082, -0.316103, -0.2291398, -0.1779351, -0.1698451, 
    -0.1029191, 0.06407309, 0.2590933, 0.4103947, 0.4399521, 0.4482691, 
    0.3419547, 0.1682236, -0.005880952, -0.1319227, -0.2295628, -0.269374, 
    -0.2548232, -0.1586155, -0.04240462, 0.0149847, 0.09130311, 0.1657495, 
    0.2079372, 0.1951603, 0.196967, 0.2172959, 0.206277, 0.1887967, 0.168354, 
    0.1560818, 0.1576443, 0.08596456, 0.07061625, 0.05484474, -0.03210163, 
    -0.1340061, -0.2365777, -0.3155491, -0.3984756, -0.3956924, -0.3679091, 
    -0.3333549, -0.1957086, -0.04876852, 0.06724715, 0.1367786, 0.1359972, 
    0.1057888, 0.05066179, 0.07027441, 0.1389756, 0.2181098, 0.31352, 
    0.1862251, 0.1254665, 0.05847448, -0.0470922, -0.1289117,
  0.3916125, 0.3229926, 0.4267035, 0.5392685, 0.524327, 0.5492296, 0.5771756, 
    0.6223092, 0.7376413, 0.7037544, 0.467751, 0.2250923, 0.122472, 0.104665, 
    0.2081819, 0.392426, 0.1596117, 0.05757809, 0.2411404, 0.1692009, 
    0.08952856, 0.02338326, -0.08078337, -0.2151592, -0.3325739, -0.4314828, 
    -0.5381241, -0.6256723, -0.6447968, -0.5849504, -0.4896541, -0.4002829, 
    -0.2988992, -0.3868704, -0.4869523, -0.6200895, -0.5494356, -0.40593, 
    -0.1909237, -0.2299695, -0.2648821, -0.3098526, -0.2354708, -0.1412816, 
    -0.07471275, -0.01885343, 0.02611685, 0.02146244, -0.02052951, 
    -0.03058815, -0.05272365, -0.08721256, -0.1080459, -0.08097881, 
    -0.01172429, 0.09364682, 0.183165, 0.2973089, 0.3746201, 0.4239365, 
    0.4501084, 0.414057, 0.3807562, 0.3207464, 0.2487901, 0.1502061, 
    0.06968848, -0.001828447, -0.05013575, -0.1130752, -0.07298729, 
    -0.04766178, -0.04103743, -0.1048721, -0.1630589, -0.2198949, -0.275917, 
    -0.2878148, -0.2669326, -0.297141, -0.2421116, -0.1340876, -0.0711644, 
    -0.07583562, -0.1587132, -0.2616917, -0.3571833, -0.3470107, -0.2782608, 
    -0.15829, -0.02650291, 0.08012158, 0.1696399, 0.2361763, 0.2534614, 
    0.2686307,
  0.5282497, 0.4383083, 0.4302681, 0.4039499, 0.3570094, 0.3303005, 
    0.3097274, 0.3335557, 0.4401636, 0.4876413, 0.3749295, 0.1152451, 
    -0.1078018, -0.1463596, -0.01231015, 0.1696715, 0.2994082, 0.405561, 
    0.5179462, 0.5858338, 0.5858669, 0.4803979, 0.3402288, 0.1989691, 
    0.1225698, 0.1129825, 0.04406953, -0.02479434, -0.09487915, -0.1006725, 
    -0.06665587, -0.1046931, -0.1875706, -0.2064025, -0.4459531, -0.4026911, 
    -0.4294491, -0.3762264, -0.2761123, -0.1674047, -0.1032119, -0.01506078, 
    0.1141547, 0.2232857, 0.2332466, 0.1210719, -0.00759016, -0.04863831, 
    -0.01167536, 0.07766366, 0.2320745, 0.3697373, 0.2889104, 0.2507433, 
    0.2075142, 0.2677678, 0.3586695, 0.4116807, 0.4437445, 0.4299749, 
    0.4190049, 0.3477484, 0.2413519, 0.1171006, -0.06512597, -0.2370661, 
    -0.4044651, -0.5488011, -0.6793351, -0.7035701, -0.6796116, -0.6306368, 
    -0.6002169, -0.7034721, -0.8351291, -0.8917859, -0.7527885, -0.586838, 
    -0.5201715, -0.4646215, -0.3687718, -0.3864151, -0.3542699, -0.3398493, 
    -0.36996, -0.4087458, -0.3578669, -0.2442438, -0.1086318, 0.03420672, 
    0.172488, 0.3592719, 0.545714, 0.7016222, 0.7269314, 0.6514919,
  0.2349066, 0.08622494, 0.007058278, -0.005295247, -0.05719954, -0.2375869, 
    -0.4336318, -0.5667859, -0.6504285, -0.7189019, -0.8177952, -0.9280815, 
    -0.8857638, -0.7645075, -0.5401422, -0.3201226, -0.1291395, -0.007476211, 
    0.05769312, -0.01820219, -0.07375216, -0.1146702, -0.1686903, -0.1506237, 
    -0.050933, 0.02527142, 0.003900766, -0.13482, -0.2938854, -0.4745336, 
    -0.6733941, -0.755572, -0.8140029, -0.8956923, -0.9183648, -0.8905818, 
    -0.875754, -0.8282931, -0.7266008, -0.5122457, -0.3458881, -0.2598362, 
    -0.08330655, 0.09379315, 0.1361434, 0.0921495, -0.003488779, -0.06305909, 
    -0.004790783, 0.1581318, 0.3640081, 0.5257107, 0.5643013, 0.5051377, 
    0.3982854, 0.3058865, 0.1798122, -0.02048063, -0.203635, -0.2743382, 
    -0.1780166, -0.07258043, -0.1400771, -0.4036188, -0.7039279, -0.9062878, 
    -1.070334, -1.183453, -1.243251, -1.208632, -1.116379, -1.055637, 
    -1.057216, -1.148687, -1.295432, -1.386887, -1.341916, -1.158794, 
    -0.9624076, -0.8262586, -0.719618, -0.6866101, -0.584006, -0.4715549, 
    -0.4746638, -0.4388239, -0.2329645, -0.01940657, 0.1738714, 0.3310492, 
    0.4703884, 0.6522569, 0.7518176, 0.7096788, 0.5529078, 0.4171331,
  0.08409274, -0.1581272, -0.351747, -0.4178118, -0.5257542, -0.7462621, 
    -0.9314027, -1.026569, -1.052382, -1.148297, -1.267242, -1.341786, 
    -1.36192, -1.395969, -1.48508, -1.599794, -1.730556, -1.838205, -1.89771, 
    -1.886399, -1.759429, -1.591216, -1.406646, -1.206565, -1.028065, 
    -0.8991591, -0.8784398, -0.8902398, -0.8741753, -0.8402236, -0.8316133, 
    -0.9350476, -1.05772, -1.060504, -0.8686256, -0.6579485, -0.60466, 
    -0.7308154, -0.8446827, -0.8002496, -0.6476126, -0.5516486, -0.5025115, 
    -0.4131403, -0.2794986, -0.2007222, -0.2240131, -0.278863, -0.2806208, 
    -0.1438375, 0.09572959, 0.279031, 0.3346951, 0.2884548, 0.1889923, 
    0.04226339, -0.1174697, -0.2757379, -0.3904189, -0.3943253, -0.2674697, 
    -0.2135309, -0.471555, -0.8584853, -1.050819, -1.079091, -1.17966, 
    -1.336936, -1.422222, -1.434852, -1.372271, -1.258518, -1.103407, 
    -1.041916, -1.116835, -1.202903, -1.130523, -0.962424, -0.8397844, 
    -0.7689834, -0.6432347, -0.5011449, -0.4420303, -0.494374, -0.4841362, 
    -0.4279839, -0.3654353, -0.3101618, -0.2447321, -0.1396377, 0.08064225, 
    0.346251, 0.4678493, 0.4374132, 0.3582953, 0.2530056,
  -0.2352432, -0.3834691, -0.3102107, -0.1796932, -0.3105199, -0.6718969, 
    -0.891151, -0.8498583, -0.8094292, -0.8900604, -0.9701061, -0.945025, 
    -0.9726453, -1.075006, -1.193056, -1.288255, -1.364329, -1.444146, 
    -1.515777, -1.534071, -1.447987, -1.290337, -1.152593, -1.025396, 
    -0.8858126, -0.8012424, -0.7514215, -0.6887912, -0.5254773, -0.3485243, 
    -0.3291397, -0.5420954, -0.7831767, -0.7785382, -0.5411029, -0.3668671, 
    -0.4568892, -0.6888719, -0.8482318, -0.8414111, -0.7291393, -0.66646, 
    -0.6770887, -0.5933323, -0.4801822, -0.5736063, -0.7430398, -0.8279197, 
    -0.8234594, -0.6986378, -0.4578993, -0.2829969, -0.2882052, -0.2522516, 
    -0.1650609, -0.2340713, -0.4401259, -0.5676488, -0.6164607, -0.651682, 
    -0.6817439, -0.8099501, -1.160438, -1.468918, -1.488108, -1.405409, 
    -1.507248, -1.66506, -1.654839, -1.505572, -1.342193, -1.133616, 
    -0.9119034, -0.8614638, -0.9881411, -1.067617, -0.9552789, -0.7012098, 
    -0.5367243, -0.5046768, -0.4695213, -0.3429744, -0.2470434, -0.2309952, 
    -0.2819228, -0.2907444, -0.290956, -0.3042859, -0.2226127, 0.01435006, 
    0.2745876, 0.393712, 0.3998317, 0.3121688, 0.1721951, -0.01445854,
  -0.1792698, -0.04985905, 0.02657318, -0.1018448, -0.4207249, -0.7325735, 
    -0.7660041, -0.6444058, -0.6586471, -0.7366743, -0.6791391, -0.5753303, 
    -0.6416879, -0.8391814, -1.040614, -1.194472, -1.29968, -1.325624, 
    -1.291135, -1.252496, -1.16856, -1.000705, -0.815321, -0.6409234, 
    -0.4517143, -0.2960829, -0.2017957, -0.1213108, -0.02777243, -0.03504801, 
    -0.2031312, -0.3960347, -0.4829326, -0.4277558, -0.3685107, -0.4527068, 
    -0.6404839, -0.756988, -0.8050675, -0.8038468, -0.7216516, -0.6952844, 
    -0.7942433, -0.7511773, -0.6129448, -0.7297099, -0.9193254, -0.952984, 
    -0.9945694, -0.984543, -0.7575738, -0.4832574, -0.4413141, -0.4758357, 
    -0.4367406, -0.4665909, -0.5584528, -0.6661514, -0.7804254, -0.898801, 
    -0.95842, -1.094471, -1.327984, -1.43648, -1.345464, -1.260259, 
    -1.370562, -1.506662, -1.382476, -1.11161, -0.8536676, -0.6358621, 
    -0.4803445, -0.4737041, -0.5974827, -0.6187062, -0.4715385, -0.2697492, 
    -0.126682, -0.1339738, -0.2048399, -0.1873429, -0.1785212, -0.2791724, 
    -0.4163306, -0.3999568, -0.2129124, -0.01509333, 0.1226022, 0.253266, 
    0.2996039, 0.2240831, 0.1347439, 0.05113387, -0.07065976, -0.1939509,
  0.183816, 0.2174096, -0.03099513, -0.3482966, -0.5405321, -0.5056038, 
    -0.3649468, -0.2308645, -0.1801481, -0.09456873, 0.004878044, 
    -0.07695866, -0.361659, -0.6342664, -0.8725154, -1.029416, -1.096165, 
    -1.069537, -0.9675186, -0.8679582, -0.7659883, -0.6211642, -0.5012585, 
    -0.431532, -0.3383679, -0.2513399, -0.2224665, -0.2148004, -0.2058649, 
    -0.2524476, -0.3341694, -0.3412986, -0.2827201, -0.3167858, -0.4690638, 
    -0.5769739, -0.5571661, -0.5220909, -0.5443244, -0.5224977, -0.4389215, 
    -0.4722381, -0.6395569, -0.5766175, -0.3753479, -0.5192928, -0.9151423, 
    -1.175184, -1.226649, -1.033794, -0.6685115, -0.4067764, -0.3534398, 
    -0.3511286, -0.3210993, -0.2252496, -0.2243056, -0.497206, -0.8445041, 
    -0.9986056, -1.058469, -1.216802, -1.354042, -1.345839, -1.228977, 
    -1.148101, -1.178782, -1.186822, -0.9702206, -0.5908747, -0.3282776, 
    -0.2823792, -0.2974014, -0.316184, -0.3662002, -0.2638402, -0.0844779, 
    0.01819086, 0.07302499, 0.04937553, -0.04185128, -0.08757091, -0.1020236, 
    -0.2187881, -0.2796769, -0.1447971, 0.04903424, 0.1626085, 0.1435004, 
    0.07123482, 0.006700277, -0.0508517, -0.07645404, -0.1140517, -0.1693249, 
    -0.07025313,
  0.2538025, 0.01426792, -0.2093322, -0.2624085, -0.2496972, -0.1694884, 
    -0.04639292, 0.1062443, 0.212234, 0.1141381, -0.1577203, -0.5447652, 
    -0.8590558, -1.053636, -1.228212, -1.314556, -1.199501, -1.005556, 
    -0.7972871, -0.6910698, -0.6724664, -0.6520725, -0.6603894, -0.652756, 
    -0.5768282, -0.447678, -0.329188, -0.2233129, -0.03044248, 0.1961529, 
    0.325417, 0.376687, 0.2891545, 0.07813597, -0.04427528, 0.003087521, 
    0.01645041, -0.1080613, -0.1936245, -0.1737361, -0.1898172, -0.3152244, 
    -0.4455297, -0.4208876, -0.4163954, -0.6043347, -0.8427625, -1.124794, 
    -1.06983, -0.61301, -0.155751, 0.01238054, 0.1677842, 0.3208278, 
    0.274555, 0.1680283, -0.01299381, -0.4055556, -0.6796115, -0.8144585, 
    -0.9822807, -1.074745, -0.9507867, -0.7772352, -0.6877656, -0.5911676, 
    -0.4908097, -0.3787653, -0.1732483, 0.02823281, -0.001356602, -0.1179743, 
    -0.0619359, 0.006602526, 0.103575, 0.3528755, 0.5454535, 0.3625269, 
    0.1411886, 0.09623504, 0.003689051, 0.01524496, 0.07675219, 0.01312935, 
    -0.01856017, 0.01955831, -0.03887272, -0.1396701, -0.2149304, -0.2585015, 
    -0.2391004, -0.1855848, -0.07930243, 0.04294705, 0.1370387, 0.2634218,
  -0.2010472, -0.2700419, -0.1330464, -0.08185816, -0.06540322, 0.09872437, 
    0.1672301, 0.1383891, 0.1105082, -0.3018618, -0.7357483, -0.9171283, 
    -1.006663, -1.116884, -1.221799, -1.136448, -0.8874077, -0.5816461, 
    -0.3700737, -0.4171278, -0.482004, -0.5045626, -0.5261772, -0.3707734, 
    -0.08942586, 0.2131294, 0.4837185, 0.7045842, 0.9051861, 0.8724223, 
    0.6420515, 0.4705179, 0.2894795, 0.1521261, 0.1971455, 0.1952574, 
    0.09349966, 0.07232618, 0.08741379, 0.05782318, -0.04554629, -0.07970917, 
    -0.09432516, -0.2037327, -0.4145238, -0.6208878, -0.7468154, -0.8411515, 
    -0.7663466, -0.4312392, -0.03493391, 0.336404, 0.7226996, 0.8486599, 
    0.6047634, 0.4384711, 0.2544866, -0.0564183, -0.2952527, -0.5568414, 
    -0.7861056, -0.6745822, -0.465679, -0.3520888, -0.1951878, -0.02866757, 
    0.08588326, 0.1286399, 0.1115987, 0.02890062, 0.07489681, 0.2164168, 
    0.3680446, 0.4634874, 0.5741806, 0.7501082, 0.7407823, 0.388715, 
    0.06942844, 0.04983175, 0.05948353, 0.1477814, 0.2892524, 0.1866157, 
    -0.09437382, -0.214898, -0.3122938, -0.3546114, -0.3785372, -0.3372613, 
    -0.1724663, -0.0743382, 0.04424906, 0.2074002, 0.2015895, 0.001752138,
  0.09483504, 0.3874295, 0.5061308, 0.4335395, 0.4861436, 0.7728618, 
    0.6606221, 0.4373963, 0.2172139, -0.4261775, -0.7256565, -0.5977921, 
    -0.6434138, -0.7537003, -0.7925504, -0.4785372, -0.10051, 0.05080843, 
    0.09758562, -0.04619694, -0.1192275, -0.08968653, 0.01840267, 0.3205186, 
    0.6201605, 0.8274847, 0.9289658, 0.9313585, 0.9144639, 0.7473904, 
    0.6168728, 0.667979, 0.5618429, 0.4850526, 0.5897732, 0.5049262, 
    0.3404889, 0.3097601, 0.3264918, 0.3066995, 0.3140407, 0.3307562, 
    0.04024535, -0.2490614, -0.5637099, -0.8504449, -0.9744034, -0.8424535, 
    -0.3895887, 0.1704209, 0.749311, 1.257872, 1.524636, 1.360265, 0.9954697, 
    0.7998969, 0.5605576, 0.2039008, 0.001052439, -0.2048883, -0.1684299, 
    0.09522557, 0.2185817, 0.3340766, 0.4559188, 0.3645453, 0.233279, 
    0.2495058, 0.3071558, 0.3857365, 0.5906355, 0.6838975, 0.5775009, 
    0.5845486, 0.7406846, 0.9233344, 0.9722278, 0.4768175, 0.1278266, 
    0.1049098, 0.3088487, 0.3657497, 0.292117, 0.03697371, -0.3713758, 
    -0.6100314, -0.574924, -0.3854383, -0.3214082, -0.2386936, 0.00990665, 
    0.139643, 0.1383247, 0.116531, 0.06130636, -0.02223861,
  0.64949, 0.773676, 0.6652777, 0.7411077, 0.8965603, 0.8156685, 0.5808375, 
    0.3401475, -0.02966034, -0.4702691, -0.4200575, -0.165077, -0.2551325, 
    -0.2185925, -0.06110555, 0.4055772, 0.6850205, 0.5629828, 0.4480252, 
    0.3330675, 0.1727486, 0.1579537, 0.2834096, 0.4701443, 0.499311, 
    0.5097765, 0.600841, 0.6353463, 0.6162546, 0.6796658, 0.7439887, 
    0.6183051, 0.4852152, 0.4599879, 0.489382, 0.3688095, 0.3449001, 
    0.364529, 0.4063584, 0.3422959, 0.3101672, 0.0772078, -0.3722223, 
    -0.6783583, -0.9710504, -1.034446, -0.7635146, -0.3516169, 0.2907823, 
    0.991173, 1.470226, 1.683946, 1.61767, 1.442768, 1.147456, 0.8398871, 
    0.5370713, 0.3823675, 0.34171, 0.2549261, 0.3299098, 0.4328232, 
    0.4452094, 0.4889594, 0.271072, 0.02183688, 0.01631951, 0.2064397, 
    0.5047145, 0.7327418, 0.8940043, 0.7974554, 0.6807236, 0.7861598, 
    0.8401474, 1.177159, 1.266092, 0.443696, -0.1334691, 0.05958104, 
    0.5036077, 0.3269966, 0.07416439, -0.01110566, -0.3460178, -0.4570203, 
    -0.2078341, 0.09384227, 0.06757258, 0.04755307, 0.08669695, 0.05258235, 
    0.07766373, 0.06050879, 0.171609, 0.3808375,
  0.7369738, 0.9129989, 1.028331, 1.138568, 0.893061, 0.4967719, 0.2100368, 
    -0.1678928, -0.210292, -0.2777887, -0.06748599, 0.1461046, -0.0322158, 
    -0.1337132, 0.06946062, 0.5058703, 0.5954211, 0.4163681, 0.3220484, 
    0.1195095, -0.06901646, 0.009157419, 0.107091, 0.1036723, 0.137738, 
    0.1736917, 0.2404728, 0.3857365, 0.5227966, 0.7822535, 0.7613553, 
    0.4067165, 0.4541612, 0.6241807, 0.460574, 0.2813097, 0.2742132, 
    0.4213488, 0.4473742, 0.291759, 0.08279073, -0.1800842, -0.4375548, 
    -0.5299208, -0.6918679, -0.6285536, -0.2947807, 0.0931586, 0.7918891, 
    1.310574, 1.332384, 1.299311, 1.262071, 1.194868, 0.9907661, 0.6988716, 
    0.5506781, 0.6017849, 0.6315374, 0.5686796, 0.5024846, 0.3418076, 
    0.181863, 0.06124127, -0.1126518, 0.03508568, 0.3490342, 0.6881614, 
    1.170877, 1.311241, 1.369786, 1.128185, 0.8585883, 0.9403427, 0.9239039, 
    1.195454, 0.8163195, -0.168918, -0.4020886, -0.04806858, 0.365359, 
    0.2133245, 0.1336533, 0.0672636, -0.2071993, -0.1070204, 0.2477484, 
    0.33004, 0.07219499, 0.07898211, 0.04600686, -0.1387424, -0.01533741, 
    0.06332457, 0.2438909, 0.4856553,
  0.8666117, 1.008018, 1.170845, 0.8906527, 0.2418239, 0.1568625, 0.0763129, 
    -0.1859919, -0.05400944, 0.01850033, 0.0644958, 0.2058697, 0.1249459, 
    -0.2188206, 0.06150186, 0.5007918, 0.5077093, 0.4152935, 0.3547304, 
    0.05606532, -0.06232667, 0.06988382, -0.04556251, -0.107167, 0.07758236, 
    0.1755314, 0.2639432, 0.4382753, 0.6745386, 0.8013775, 0.625499, 
    0.4136341, 0.4972603, 0.588097, 0.3648384, 0.2871853, 0.4935815, 
    0.569607, 0.4399519, 0.1310329, 0.04200292, -0.09562731, -0.2691302, 
    -0.2909236, -0.3173726, -0.2761943, -0.09307241, 0.2160258, 0.6505151, 
    0.7850368, 0.6818955, 0.8034286, 0.8950471, 0.8275988, 0.7098254, 
    0.5313261, 0.4713001, 0.5426054, 0.5326281, 0.3946723, 0.0377712, 
    -0.2678766, -0.3377171, -0.2676488, -0.01590711, 0.4145131, 0.7591256, 
    1.045844, 1.363715, 1.214008, 1.021186, 0.7158638, 0.5279241, 0.6997008, 
    0.6478784, 0.6600037, 0.2051213, -0.1669813, -0.1552464, -0.1125705, 
    0.1664333, 0.05993915, 0.03609478, 0.2295517, 0.2691839, 0.3867784, 
    0.3513618, 0.2625595, 0.03033304, -0.05806208, -0.1436253, -0.2073947, 
    -0.02585185, 0.1760361, 0.4419383, 0.6836696,
  0.8068955, 0.7734485, 0.6895943, 0.2193789, 0.02647561, 0.1583278, 
    0.1172471, 0.1057236, 0.02432716, 0.0117619, -0.09652305, -0.1073792, 
    -0.07521695, -0.1356989, 0.1420841, 0.2563095, 0.2923608, 0.2222276, 
    0.1039655, 0.03607845, 0.008588314, -0.006336689, -0.1512747, 
    -0.02463055, 0.09931135, 0.1017528, 0.2665315, 0.5350537, 0.7884059, 
    0.7663023, 0.5597112, 0.5050238, 0.5610616, 0.5796492, 0.3407985, 
    0.2457626, 0.4456487, 0.4192162, 0.1716735, -0.08488512, 0.08410978, 
    0.05570841, -0.2083225, -0.3934464, -0.4650283, -0.3651588, -0.09526968, 
    0.2506125, 0.4047139, 0.5211208, 0.6823511, 0.7274853, 0.5718533, 
    0.5463163, 0.492296, 0.4069282, 0.3544053, 0.2929469, 0.1289009, 
    -0.1668024, -0.4188043, -0.3653865, -0.1670954, 0.08353939, 0.4082302, 
    0.7958604, 1.017914, 0.997732, 0.9670519, 0.8037056, 0.6754339, 0.587055, 
    0.6517191, 0.5429471, 0.2471962, 0.2844834, 0.1463327, 0.1258733, 
    0.07299256, -0.08361542, 0.008751005, 0.007302403, -0.0009983703, 
    0.2850368, 0.2788031, 0.1029079, 0.07961631, 0.06181026, -0.0664773, 
    -0.08346963, -0.09937143, 0.03884482, 0.2073019, 0.4130635, 0.5484641, 
    0.6944444,
  0.4666939, 0.4256463, 0.1888137, -0.02770758, 0.09517682, 0.1591254, 
    0.06299902, 0.09524187, 0.02986097, 0.0656358, 0.05341244, -0.2572484, 
    -0.226096, 0.07079506, 0.4121361, 0.1813588, 0.2311959, 0.241775, 
    0.2437444, 0.1848249, 0.05639124, -0.03027868, -0.1546597, -0.104692, 
    -0.1256719, 0.1130643, 0.3960886, 0.5385361, 0.5937276, 0.4179301, 
    0.2278428, 0.276036, 0.1982367, 0.09198713, -0.08013201, -0.002284288, 
    0.0315218, -0.3199763, -0.281158, -0.1441941, -0.04749918, -0.4392304, 
    -0.7419815, -0.7930555, -0.5620337, -0.274143, -0.06983042, 0.3108664, 
    0.4979923, 0.5892034, 0.531863, 0.3341583, 0.1795355, 0.1774033, 
    0.100727, 0.01719832, -0.1497451, -0.2462617, -0.2865451, -0.3461319, 
    -0.2502171, -0.123622, -0.0257867, 0.2258734, 0.4651475, 0.5856065, 
    0.653852, 0.6060493, 0.6021923, 0.6231878, 0.6515403, 0.5268168, 
    0.4039989, 0.1616492, 0.09986448, 0.3610945, 0.4089791, 0.1903916, 
    0.09755313, 0.02732193, 0.008327961, -0.02119693, 0.006228209, 0.1097113, 
    -0.08382726, -0.141721, 0.2607532, 0.08946371, -0.1438694, 0.04727626, 
    0.05917406, 0.1650987, 0.2996526, 0.4239204, 0.4472601, 0.4856224,
  0.06856537, 0.1369905, -0.0536027, -0.01318908, 0.07533626, 0.06295031, 
    0.02004659, -0.08866107, -0.09328341, -0.0654186, -0.2380753, -0.540647, 
    -0.3619847, 0.08449888, 0.323595, 0.217525, 0.1456819, 0.1421332, 
    0.1850696, -0.1188045, -0.1679573, -0.3019414, -0.4631886, -0.5398002, 
    -0.643055, -0.1847382, -0.002235413, 0.004778862, -0.01786089, 
    -0.1506572, -0.2725811, -0.1825252, -0.1804097, -0.4583062, -0.4336643, 
    -0.2390354, -0.1965225, -0.3302789, -0.1028371, 0.01032972, -0.3971567, 
    -0.9085016, -0.9548392, -0.7000709, -0.3057349, -0.1623759, 0.08454776, 
    0.4485135, 0.3416774, 0.09732533, -0.1038954, -0.05698788, -0.1287652, 
    -0.1864151, -0.26218, -0.2627658, -0.3057345, -0.2877009, -0.1913629, 
    -0.08519417, 0.005316973, -0.03210151, 0.06607521, 0.2388618, 0.3253365, 
    0.3905544, 0.4657984, 0.5691187, 0.6716573, 0.5930114, 0.5790143, 
    0.4115348, 0.2228789, 0.1168232, 0.05691099, 0.2271104, 0.1257921, 
    0.04294693, -0.006825149, 0.05783963, 0.1140084, 0.05144304, 0.03682745, 
    -0.06314027, -0.08473897, 0.1183696, 0.3011179, 0.002777576, 0.01825619, 
    0.03446722, -0.1963596, -0.1106987, -0.000705719, 0.01229906, 0.02977943, 
    0.1019964,
  -0.1759329, -0.08648014, -0.2114477, 0.06081796, 0.02457166, -0.06309152, 
    -0.0693574, -0.1770887, -0.1637262, -0.1121475, -0.310667, -0.6346574, 
    -0.2229061, 0.3701439, 0.387413, 0.3549752, 0.3193307, 0.1159616, 
    -0.1708226, -0.4739802, -0.3233128, -0.4853246, -0.7567763, -0.9489639, 
    -0.8819878, -0.4473205, -0.4868388, -0.4024794, -0.4524957, -0.6663955, 
    -0.5415423, -0.5882215, -0.6745176, -0.6635959, -0.61428, -0.6799209, 
    -0.4669979, -0.3722878, -0.08649635, -0.08241129, -1.168511, -1.199517, 
    -0.9099014, -0.6143126, -0.2656636, -0.354954, -0.1539774, 0.07125139, 
    -0.1901259, -0.2361058, -0.2194228, -0.1575087, -0.2862523, -0.2761122, 
    -0.2262588, -0.2416558, -0.1813856, -0.1528375, -0.1674697, -0.121034, 
    -0.1378798, -0.04811752, 0.07665479, 0.09416771, 0.2073019, 0.3111429, 
    0.3951275, 0.4073188, 0.3847275, 0.2987251, 0.1829209, 0.06970501, 
    -0.06050348, -0.1059623, -0.06078053, -0.005946279, -0.02380109, 
    -0.07474512, 0.09630013, 0.1186957, -0.01686746, 0.007253885, 
    -0.06063378, -0.1470596, -0.03333926, 0.08285522, 0.1512313, -0.1915259, 
    -0.1411352, -0.3083713, -0.5131893, -0.4530005, -0.4409885, -0.3114963, 
    -0.2411194, -0.2360568,
  -0.2832901, -0.3113012, -0.3633194, 0.09325624, -0.08009994, -0.355702, 
    -0.1904188, -0.2267962, -0.157004, -0.2564996, -0.228456, -0.1843157, 
    -0.03420067, 0.2511826, 0.4577737, 0.4682565, 0.2820582, 0.04345179, 
    -0.1446509, -0.1284726, -0.2058325, -0.4554255, -0.6701391, -0.8854554, 
    -0.6870337, -0.3536676, -0.4863173, -0.08555293, -0.09316957, -0.5402563, 
    -0.2562723, -0.187115, -0.3319716, -0.5591528, -0.7683814, -0.5478573, 
    -0.1779675, -0.2905328, -0.1070693, -0.1482801, -1.579075, -1.137977, 
    -0.5158265, -0.3699436, -0.1799535, -0.1746962, 0.07683396, 0.2339791, 
    0.1684191, 0.1485787, 0.1406686, 0.2175075, 0.2853136, 0.2989529, 
    0.3012966, 0.267361, 0.2633083, 0.2236598, 0.1697374, 0.1351346, 
    0.08629018, 0.1442654, 0.149604, 0.2060819, 0.2836697, 0.1971943, 
    0.2179625, 0.2085719, 0.09641361, 0.01127338, -0.1332736, -0.2010312, 
    -0.2497125, -0.3388567, -0.1320863, -0.04800358, -0.1540583, -0.1255915, 
    -0.03509665, -0.04938704, 0.03225368, -0.004709303, -0.02010643, 
    -0.0445205, -0.1363823, -0.4655173, -0.329514, -0.2041721, -0.2766168, 
    -0.5344458, -0.7087619, -0.6583714, -0.6287978, -0.4398491, -0.3573787, 
    -0.3946345,
  -0.26913, -0.3660538, -0.4239964, -0.02996957, -0.2160863, -0.3007216, 
    -0.1891494, -0.1133518, -0.1939996, -0.2639215, -0.3382056, 0.2048926, 
    0.3846941, 0.3532658, 0.3552351, 0.3760366, 0.1888132, 0.08165145, 
    -0.112473, -0.1386781, -0.202529, -0.3811095, -0.5242407, -0.4809465, 
    -0.1526754, -0.07551008, -0.1839085, 0.02297624, -0.1425185, -0.3890843, 
    0.07919395, -0.0003473163, -0.03006727, -0.7704647, -0.7665746, 
    -0.1427301, -0.09162338, -0.07393131, -0.2198135, -0.913336, -1.478456, 
    -0.6613499, -0.2328343, -0.1395562, 0.0641709, 0.1346787, 0.1297145, 
    0.03568786, 0.05902767, -0.04746634, -0.1129937, 0.04460728, 0.15421, 
    0.1483183, 0.1388942, 0.1423123, 0.1323024, 0.1520616, 0.1474065, 
    0.1218206, 0.1250758, 0.06601009, 0.03119576, 0.03383243, -0.02699113, 
    0.01443124, -0.03910065, -0.125885, -0.2079325, -0.353163, -0.421962, 
    -0.4449279, -0.4613988, -0.4831274, -0.3853081, -0.2438695, -0.07254779, 
    -0.09479719, -0.1391331, -0.1553115, -0.067958, 0.1239528, 0.1175726, 
    -0.2467015, -0.4253311, -0.9170952, -0.4918842, -0.0376687, -0.1952528, 
    -0.4240614, -0.5009007, -0.4036838, -0.3810112, -0.4015522, -0.3161845, 
    -0.3583226,
  -0.1243713, -0.2162821, -0.1902887, -0.04733626, 0.01231542, 0.04546973, 
    0.09179135, 0.03404395, -0.05085182, 0.04345191, -0.06161094, -0.0217824, 
    0.33992, 0.6436625, 0.4256454, 0.3358178, 0.2617292, 0.07842851, 
    -0.1499898, -0.3070691, -0.2905335, -0.4028542, -0.5289934, -0.3804092, 
    -0.2479386, -0.1643283, 0.09361428, -0.03132063, -0.8848524, -0.5929906, 
    -0.2430068, -0.08713119, -0.1149958, -1.069765, -0.8016655, -0.2569389, 
    -0.1922255, 0.04708105, -0.1828666, -0.8035381, -0.8543836, -0.4319717, 
    -0.351096, -0.3014866, -0.1007377, -0.1217338, -0.316672, -0.5499728, 
    -0.5454317, -0.6672904, -0.7588106, -0.7850965, -0.8113171, -0.7544488, 
    -0.715256, -0.6887587, -0.6493382, -0.6007543, -0.4962946, -0.368251, 
    -0.2608128, -0.1916393, -0.1037489, -0.100917, -0.09312081, -0.05090141, 
    -0.1176331, -0.1124732, -0.2195044, -0.3432999, -0.3335512, -0.2828836, 
    -0.2266335, -0.1385145, -0.08379459, -0.1995986, -0.2905329, -0.1563043, 
    -0.05588118, 0.06630307, 0.1728623, 0.09592546, -0.1884008, -0.3396378, 
    -0.2261934, -0.07730046, 0.2007269, 0.2024523, -0.1947159, -0.1906305, 
    0.01161556, 0.0561794, -0.09245312, -0.1814182, 0.07300901, 0.01076865,
  0.1605413, 0.09511113, 0.1201606, 0.05230567, 0.0581001, 0.09708118, 
    0.09600684, 0.08350682, 0.0272572, -0.02293846, 0.06495225, -0.1018929, 
    0.02112007, 0.6467524, 0.7093191, 0.5781026, 0.3893986, 0.1051695, 
    0.04421651, -0.08381081, -0.1591361, -0.1632712, -0.1208706, -0.1034231, 
    -0.1711149, -0.1391008, -0.06670475, -0.06690006, -0.6357646, -0.6021707, 
    -0.2598849, -0.1320042, -0.3852104, -0.71052, -0.5436258, -0.1971573, 
    0.003998399, -0.0778701, -0.2056371, -0.3353571, -0.364654, -0.2103408, 
    -0.1233942, -0.05832231, 0.02045345, -0.01976466, 0.02930772, 0.07805443, 
    0.04545355, -0.06081295, -0.1828994, -0.2862685, -0.3338434, -0.4248101, 
    -0.5479057, -0.5788465, -0.5676811, -0.5582249, -0.5116429, -0.4765192, 
    -0.512831, -0.5086969, -0.5336644, -0.5231826, -0.3326551, -0.3565979, 
    -0.3907933, -0.3673396, -0.5352757, -0.6072805, -0.5495825, -0.2846733, 
    -0.1872451, -0.2273166, -0.007167101, -0.01115462, -0.2392959, 
    0.05422664, 0.1428005, -0.01652569, -0.2433974, -0.2650936, -0.008566618, 
    0.2022243, 0.2490505, 0.3167746, 0.3180447, 0.2686632, 0.05989027, 
    -0.001665354, 0.1396104, 0.1719835, 0.09004998, -0.1350803, 0.03345811, 
    0.08918738,
  0.05158985, 0.04822052, 0.001801252, 0.1125273, 0.2532662, 0.5395126, 
    0.4888779, 0.2800076, 0.05390072, -0.1057673, -0.00267446, 0.08295298, 
    0.1984, 0.6718683, 0.9427662, 0.8009529, 0.6227975, 0.4320583, 0.1425238, 
    -0.190484, -0.2972549, -0.2896872, -0.3546281, -0.2099028, -0.1434612, 
    -0.2951393, -0.7488501, -0.1313044, 0.1633898, -0.3167052, -0.5973363, 
    -0.695204, -0.8565166, -0.2814183, -0.2299209, -0.3948134, -0.09665257, 
    -0.06738824, -0.02458236, 0.017361, 0.03314885, -0.001307487, 0.06544042, 
    0.1332628, 0.1227973, 0.1165304, 0.1674418, 0.1865988, 0.1400168, 
    0.1393168, 0.1139097, 0.04577851, 0.07216239, 0.1038682, 0.1249454, 
    0.1001573, 0.04223084, 0.02002978, -0.004889011, -0.01473522, 
    -0.06982994, -0.1065322, -0.1687717, -0.2858939, -0.2971408, -0.3624567, 
    -0.5230523, -0.6305717, -0.556109, -0.6964247, -0.7154351, -0.303863, 
    -0.2895401, -0.4808646, -0.1830948, -0.1755262, -0.2635307, -0.3350639, 
    -0.4586644, -0.4628799, -0.4781799, -0.1265848, 0.2090433, 0.293988, 
    0.2105737, 0.1267035, 0.1215603, 0.2011337, 0.1322043, 0.128103, 
    0.1599557, 0.02505958, 0.01132286, 0.1536891, 0.1918727, -0.008208513,
  0.344542, 0.4126898, 0.4409288, 0.3754991, 0.1770291, 0.1858506, 0.2350532, 
    0.433035, 0.4444926, 0.1624451, -0.1177627, -0.1855524, 0.03419042, 
    0.3144317, 1.000578, 1.150465, 0.8617449, 0.5503201, 0.2817328, 
    -0.08049047, -0.2951553, -0.2678115, -0.4811416, -0.2030649, -0.09094048, 
    -0.3073621, -0.5667219, -0.2707574, -0.175103, -0.3038791, -0.5264215, 
    -1.150347, -1.563173, -0.7547582, -0.5197489, -0.5312879, -0.1691298, 
    -0.0775283, 0.02328548, 0.098139, -0.02541247, -0.2687879, -0.04479694, 
    0.1346625, 0.06905377, 0.1199977, 0.2187114, 0.2668884, 0.2391381, 
    0.1608016, 0.1294861, 0.0602808, -0.05737853, -0.1578019, -0.2160375, 
    -0.171669, -0.1421442, -0.1674209, -0.1796443, -0.1296282, -0.04095626, 
    0.07733798, 0.1506941, 0.1328063, 0.01478887, -0.05983639, -0.357476, 
    -0.4189021, -0.04176983, -0.4162165, -0.4280654, -0.07830957, -0.394618, 
    -0.724143, -0.718154, -0.5827368, -0.5600476, -0.7426977, -0.5955949, 
    -0.2227104, -0.09149301, 0.0515244, 0.1158798, 0.1591904, 0.2196722, 
    0.2324975, 0.2037544, 0.1873479, 0.1982856, 0.3020616, 0.439122, 
    0.3901638, 0.3401637, 0.5713811, 0.8173447, 0.5813257,
  0.5967394, 0.3519803, 0.2802191, 0.3082464, 0.1754665, -0.0006239414, 
    -0.2498596, -0.06773019, 0.4138618, 0.4386176, 0.1433206, -0.392714, 
    -0.3813043, -0.1174859, 0.3518169, 0.6358166, 0.9740658, 0.8981881, 
    0.407872, 0.0386014, -0.1045791, 0.1546984, -0.03980023, -0.2034559, 
    -0.07935143, -0.1409564, -0.03122306, -0.07008982, -0.2798883, 0.2612739, 
    0.3611436, -0.8714252, -1.51161, -1.392454, -1.160928, -0.6650933, 
    -0.1715875, -0.07612842, -0.03543842, 0.09240985, -0.1685439, -0.510406, 
    -0.3498102, -0.1866428, -0.07096899, 0.0303005, 0.1140568, 0.1682403, 
    0.1754661, 0.1299093, 0.1148052, 0.08723354, 0.03622437, -0.01803994, 
    -0.1060607, -0.1660049, -0.1942925, -0.2062557, -0.2300024, -0.2340224, 
    -0.2220106, -0.1541562, -0.1446509, -0.0129776, 0.0564723, 0.129096, 
    -0.09333301, -0.2814183, -0.07843977, -0.2402236, -0.240598, 0.1592067, 
    -0.1395563, -0.6485407, -0.775087, -0.640891, -0.5890192, -0.5804417, 
    -0.5379939, -0.3967339, -0.2795792, -0.1264708, -0.023525, 0.04781342, 
    0.04542065, 0.05588627, 0.06140423, 0.03199339, 0.07621479, 0.1000433, 
    0.2954865, 0.4859972, 0.3381455, 0.3589465, 0.9237577, 1.076297,
  0.2949489, -0.01615136, -0.34356, -0.2096896, -0.04281151, -0.0471735, 
    -0.1160862, -0.2101781, -0.003993273, 0.5285263, 1.050824, -0.05178022, 
    -0.397629, 0.1251087, 0.4709256, 0.3612895, 0.5587506, 0.7747016, 
    0.3169374, 0.1474879, 0.1966255, 0.3991645, 0.3202745, -0.04437387, 
    -0.03259087, -0.06012917, -0.1635146, -0.05910373, 0.1693794, 0.8451932, 
    0.8617132, 0.2149677, -0.18648, -0.9346247, -1.285552, -0.7623426, 
    -0.3828017, -0.2871637, -0.1610244, -0.1127658, -0.3326064, -0.4388401, 
    -0.3233128, -0.155572, -0.03467333, 0.006895542, 0.1024685, 0.1640083, 
    0.2285428, 0.2027128, 0.1609483, 0.08943152, 0.03811288, 0.08181429, 
    0.1832139, 0.1388618, 0.03322959, 0.05023789, -0.06232643, -0.1144912, 
    -0.1218805, -0.08625269, -0.05010319, 0.02172375, 0.04094458, 0.02673578, 
    0.06789804, -0.06746972, 0.1302682, 0.08783633, -0.2763402, -0.1832085, 
    0.04639757, -0.5863825, -0.8686903, -0.7402562, -0.6340712, -0.5396703, 
    -0.4944228, -0.3331108, -0.2797905, -0.1668186, -0.04635966, 0.0390563, 
    0.09379315, 0.1464462, 0.1586208, 0.07909632, 0.02512455, -0.06314087, 
    -0.2143946, -0.2430401, -0.3875537, -0.298378, 0.1607692, 0.4214626,
  -0.1203831, 0.05609798, -0.02892807, -0.0452528, -0.2264539, -0.49968, 
    -0.4059138, -0.4239972, -0.5288458, 0.1655705, 0.9384065, 0.09216571, 
    -0.3405653, 0.08964276, 0.7139269, 0.6864855, 0.6398218, 0.9856715, 
    0.6038029, 0.1996851, 0.2744737, 0.3274199, 0.2887967, -0.1326394, 
    -0.2930233, 0.01509863, -0.002316773, -0.002511859, 0.555512, 1.282254, 
    1.142914, 1.046967, 0.6165637, -0.3419979, -0.8611221, -0.2195694, 
    0.1069444, -0.07970929, -0.05677629, -0.1675185, -0.6306045, -0.7439508, 
    -0.4991103, -0.1731175, -0.1170954, -0.0221898, 0.09004998, 0.06361759, 
    0.1565541, 0.1412543, 0.1556098, 0.1142687, 0.03921962, -0.009755135, 
    0.003103256, 0.05256605, -0.02565646, 0.0476501, 0.12851, 0.1821558, 
    0.1549261, 0.1781349, 0.2551694, 0.235167, 0.1356559, -0.1241422, 
    0.1225204, 0.2196071, 0.1849229, 0.1782173, -0.07329625, -0.09289277, 
    -0.09557915, -0.5003474, -0.509657, -0.6190971, -0.6746311, -0.5238174, 
    -0.5034562, -0.4502497, -0.4427464, -0.3110406, -0.1336317, 0.06335723, 
    0.2180934, 0.1790955, 0.1202908, 0.09885502, 0.06163216, -0.04152584, 
    -0.1895404, -0.2409897, -0.2595925, -0.3748264, -0.2978573, -0.2005914,
  -0.08311087, -0.1745985, -0.1970921, -0.2081761, -0.1214411, -0.3837621, 
    -0.5331435, -0.5973201, -0.7695527, -0.1818581, 0.1167264, -0.1999403, 
    -0.2151423, 0.08583403, 0.4416287, 0.5424424, 0.7752387, 1.35421, 
    1.075971, 0.599246, 0.7962509, 0.8307726, 0.6360136, 0.5205998, 
    0.2844186, 0.07602024, -0.01045513, -0.1083558, 0.4185168, 1.365196, 
    1.365848, 1.203803, 1.220112, 0.6479924, 0.1272569, 0.2155707, 0.5164658, 
    0.3212998, 0.2556586, 0.04953861, -0.4763246, -0.7531306, -0.5950087, 
    -0.2660048, -0.1468804, -0.06812075, -0.03571516, -0.06932518, 
    0.07903099, 0.1089788, 0.1722438, 0.06783307, 0.01985133, 0.06368291, 
    -0.07806528, -0.1251517, -0.1994846, -0.2111709, -0.08482051, 0.03401136, 
    0.1237903, 0.2858181, 0.4959912, 0.5665474, 0.3738556, 0.008718014, 
    -0.05498588, 0.105154, -0.1765029, -0.432053, -0.02638912, 0.4973583, 
    0.1721296, -0.2906142, 0.005007625, -0.02380157, -0.542665, -0.7347227, 
    -0.6992079, -0.6969456, -0.7221573, -0.5920953, -0.4085016, -0.1388727, 
    0.1162546, 0.2236437, 0.2005804, 0.07403421, 0.02862406, -0.05413914, 
    -0.2597704, -0.3400602, -0.09587193, -0.01063347, 0.227322, 0.2314886,
  0.5615504, 0.5138943, 0.1940211, -0.1555393, -0.337245, -0.3733623, 
    -0.5509989, -0.6495008, -0.8370993, -0.4504941, -0.3313208, -0.6238339, 
    -0.2264054, 0.1886667, 0.1259711, 0.05749786, 0.03830767, 0.4940052, 
    0.9138126, 1.091075, 0.8273057, -0.01180536, -0.5615615, -0.4779352, 
    -0.440305, -0.5209696, -0.3085668, -0.1767144, 0.1803818, 0.4478787, 
    0.5331162, 0.5358831, 0.5938749, 0.5734164, 0.5569937, 0.3751736, 
    0.578933, 0.5110133, 0.4809027, 0.3817978, -0.06048727, -0.3669164, 
    -0.4677463, -0.3263245, -0.2107804, -0.1895888, -0.230637, -0.2407281, 
    -0.08167845, -0.005734563, 0.04087988, -0.08355045, -0.178277, 
    -0.06392155, -0.1382868, -0.2595108, -0.306695, -0.3022351, -0.3073784, 
    -0.2759984, -0.1322484, 0.008979321, 0.3586698, 0.7294378, 0.7576118, 
    0.4693304, 0.1976182, 0.1649033, 0.2172308, 0.07894945, -0.01014566, 
    0.1024034, 0.07261753, -0.3158095, -0.06896698, 0.3018663, -0.03083277, 
    -0.5519426, -0.7068577, -0.8090224, -0.8721902, -0.8227593, -0.6984756, 
    -0.4124078, -0.1492242, -0.008176103, 0.0552029, 0.009239316, 
    -0.06532073, -0.2630427, -0.4935765, -0.5944552, -0.5084534, -0.1345263, 
    -0.00772047, 0.4318142,
  -0.08892155, -0.08895373, 0.1439398, 0.1804795, -0.0701226, -0.4617081, 
    -0.3929741, -0.2745334, -0.4505913, -0.2150934, -0.1821675, -0.2225153, 
    -0.07314992, -0.03338754, -0.1834202, -0.09751606, -0.132802, -0.2400451, 
    0.139236, 0.7150499, 0.6259548, 0.2218858, 0.163227, 0.1232367, 
    0.03397885, 0.06596126, -0.1035374, -0.06663965, 0.1943304, 0.134223, 
    -0.01751855, -0.05116099, -0.1147839, -0.1162164, 0.005658627, 
    -0.1366916, 0.05097115, 0.1236598, 0.1613224, 0.2799425, 0.2117782, 
    0.1091089, -0.02285719, -0.02274323, -0.05846906, -0.09354448, 
    -0.2269914, -0.3916728, -0.2364156, -0.01628149, 0.0316515, -0.068609, 
    -0.2682184, -0.3742894, -0.3913954, -0.4077688, -0.398557, -0.3894587, 
    -0.4951553, -0.4493707, -0.30357, -0.2897515, 0.04398823, 0.6395125, 
    0.6497667, 0.6327745, 0.2379829, -0.03283429, 0.302387, 0.8630648, 
    0.6008892, -0.01286364, -0.1930068, -0.2890842, -0.3367568, -0.1474502, 
    -0.09705949, -0.2364314, -0.5098364, -0.8494358, -1.004336, -0.9362204, 
    -0.87538, -0.6294978, -0.3224669, -0.1898981, -0.1456923, -0.07853743, 
    -0.09564352, -0.4501357, -0.8220437, -1.103358, -1.156532, -0.7632875, 
    -0.1872449, -0.1866274,
  -0.4778213, -0.7662653, -0.3517306, 0.2047959, 0.1907009, -0.4056205, 
    -0.7143935, -0.4380101, -0.4408094, -0.5676324, -0.509348, -0.4290416, 
    -0.4511123, -0.5209364, -0.2741916, -0.1589572, -0.09100473, -0.2796113, 
    -0.4741268, -0.3953505, -0.08890527, 0.3994086, 0.6822047, 0.5656196, 
    0.5846624, 0.6201279, 0.2114691, -0.03088117, 0.2411242, 0.3594347, 
    0.2110133, 0.03840593, -0.1561252, -0.1279839, -0.1605035, -0.369081, 
    -0.3939832, -0.3530328, -0.3446344, -0.2338438, 0.0730083, 0.4491313, 
    0.5907331, 0.5250263, 0.3451109, 0.1696553, -0.07445216, -0.3646214, 
    -0.3445206, -0.1824112, -0.07866812, -0.01473546, -0.1454647, -0.3602107, 
    -0.485846, -0.5136611, -0.4860244, -0.5222874, -0.6606012, -0.622206, 
    -0.470318, -0.4614964, -0.1710505, 0.182579, 0.2875109, 0.5383409, 
    0.3888617, 0.04812288, 0.08871531, 0.7895291, 1.229161, 0.7966247, 
    0.2413681, 0.05463314, -0.1345592, -0.1957411, -0.07472885, -0.12678, 
    -0.2027075, -0.3543513, -0.5300028, -0.6518614, -0.7258687, -0.6920307, 
    -0.4028864, -0.1284399, -0.1084204, -0.1294489, -0.1125704, -0.3638565, 
    -0.8046767, -1.334771, -1.817486, -1.531418, -0.8810277, -0.3021052,
  -0.3397842, -0.7427463, -0.6338921, -0.2291232, 0.03824329, -0.1117893, 
    -0.52232, -0.486594, -0.3519749, -0.383583, -0.1921442, -0.3363661, 
    -0.6449437, -0.3823135, -0.3631727, -0.1549532, -0.03359926, 0.02728975, 
    -0.2039117, -0.2530166, -0.1510631, -0.0712291, -0.1431533, -0.1846572, 
    -0.03177636, 0.1589788, 0.1572047, 0.1830023, 0.4189562, 0.5256132, 
    0.5498968, 0.5126573, 0.3242623, 0.2538683, 0.246528, 0.1583279, 
    -0.0409559, -0.1276422, -0.2174206, -0.4050673, -0.3311903, 0.115294, 
    0.4741642, 0.6368597, 0.5761011, 0.2864847, 0.02733755, -0.1910539, 
    -0.4534073, -0.5993865, -0.4837296, -0.3027725, -0.236692, -0.1854224, 
    -0.134104, -0.1756241, -0.2943094, -0.4979715, -0.6877658, -0.6368382, 
    -0.475917, -0.3611872, -0.2045956, -0.06050301, 0.1600693, 0.3393011, 
    0.3848091, 0.1765895, -0.09914291, 0.06184343, 0.5613064, 0.7593045, 
    0.7079861, 0.6327908, 0.1714464, -0.01385617, -0.07827693, -0.172027, 
    -0.3082907, -0.3016982, -0.3043838, -0.1734436, -0.005621195, -0.1540589, 
    -0.286139, -0.002984047, 0.2720158, 0.3090601, 0.2132268, -0.1333225, 
    -0.553342, -0.9576715, -1.681515, -1.931809, -1.217893, -0.2848524,
  -0.1587458, -0.06408429, -0.3598035, -0.5719945, -0.3583877, -0.01626521, 
    -0.02365434, -0.06429577, -0.08070219, -0.05327702, 0.2355253, 0.4036729, 
    0.08811295, -0.1703994, -0.03810775, -0.0158584, -0.06025943, -0.1086805, 
    -0.2301649, -0.240598, -0.004693031, 0.147195, 0.1456001, 0.04794371, 
    -0.01813674, -0.02883029, 0.1135525, 0.3262153, 0.4317327, 0.4239854, 
    0.4301378, 0.5093207, 0.5209255, 0.491466, 0.4486762, 0.3689561, 
    0.3596138, 0.4054307, 0.3522242, -0.01416552, -0.09557843, 0.1596463, 
    0.4953235, 0.6973413, 0.7034123, 0.5036895, 0.3090274, 0.2134709, 
    -0.07987213, -0.583746, -0.8575413, -0.9360244, -0.9062557, -0.6139541, 
    -0.1925187, 0.07473397, 0.1034606, -0.1287496, -0.4168355, -0.4644586, 
    -0.3193251, -0.1455295, -0.05010313, -0.06092677, 0.07182065, 0.1769313, 
    0.2819118, 0.2833279, 0.1829373, 0.1230576, 0.2210231, 0.3870876, 
    0.6068793, 0.4384221, 0.4308214, 0.1588976, 0.1210394, 0.05154073, 
    -0.1721084, -0.4188043, -0.4913797, -0.3274307, 0.1418564, 0.2893171, 
    0.1746032, 0.234792, 0.4846454, 0.6475856, 0.6220808, 0.3203394, 
    -0.04541564, -0.4123101, -1.064572, -1.561464, -1.187424, -0.6050186,
  -0.3267143, 0.2941516, 0.3838649, 0.01612403, -0.1189834, 0.02613379, 
    0.1372015, 0.2279893, 0.2233672, 0.2169379, 0.2660264, 0.2944444, 
    0.1929795, 0.08749447, 0.2250107, 0.335346, 0.2647731, 0.07868913, 
    -0.1439183, -0.3977269, -0.5086644, -0.3299696, -0.04497612, 
    -0.0002170801, -0.06716049, -0.07874902, 0.0340765, 0.2201117, 0.3485948, 
    0.3328069, 0.1554797, 0.01547313, 0.1002387, 0.3335882, 0.3702256, 
    0.2535752, 0.2728135, 0.4783474, 0.5337836, 0.3943469, 0.5150988, 
    0.7317654, 0.8731065, 0.988829, 1.164382, 1.19713, 1.058214, 0.8904569, 
    0.6095161, -0.01792538, -0.6944064, -1.121181, -1.272678, -1.082558, 
    -0.5694554, -0.06903219, 0.1282165, -0.01454043, -0.1384828, -0.0130589, 
    0.1478786, 0.1108019, 0.04379326, 0.0187282, 0.2324814, 0.3043402, 
    0.2619573, 0.219005, 0.2916612, 0.5205511, 0.6820421, 0.6390569, 
    0.6802842, 0.7650986, 0.732514, 0.5528591, 0.3667262, 0.2490016, 
    0.1603623, 0.1560329, -0.02528222, -0.06143117, 0.005056381, 0.3025656, 
    0.6483014, 0.8986268, 1.074311, 1.015733, 0.8719509, 0.6651473, 
    0.4054308, 0.08280706, -0.4281467, -0.9116102, -1.083469, -0.7685602,
  -0.5354384, -0.3058811, -0.2234756, 0.05383561, 0.2879339, 0.3203721, 
    0.2214138, 0.2003689, 0.274083, 0.2729274, 0.2199978, 0.1787543, 
    0.09901828, 0.04395616, 0.1624945, 0.3086371, 0.2433864, 0.08052833, 
    -0.0945856, -0.3742406, -0.6579645, -0.6830622, -0.4110407, -0.1420301, 
    -0.07788634, -0.05070531, -0.05780166, 0.00655365, 0.1886663, 0.3485948, 
    0.3277288, 0.1354764, 0.09838307, 0.2279892, 0.2611436, 0.1506618, 
    0.01360118, -0.02349186, 0.1272082, 0.3790472, 0.8236436, 0.9368759, 
    0.9783799, 0.7571886, 1.110672, 1.543484, 1.506293, 1.353592, 1.157514, 
    0.6784124, -0.1207575, -0.9417536, -1.358778, -1.279189, -0.842307, 
    -0.3987198, -0.2224996, -0.2593648, -0.1436255, 0.16907, 0.3504506, 
    0.3749456, 0.2319771, 0.2636663, 0.29407, 0.2597275, 0.1577418, 
    0.1072535, 0.1907334, 0.3865179, 0.5602973, 0.6689236, 0.7899197, 
    0.9256293, 1.01186, 0.5870714, 0.5525661, 0.2321885, 0.08511817, 
    0.112234, 0.1744412, 0.06181091, 0.07206479, 0.2659612, 0.6510526, 
    1.132921, 1.43865, 1.408214, 1.216661, 1.09464, 0.8523061, 0.3533962, 
    -0.2635472, -0.6308649, -0.6620985, -0.5861545,
  -0.5635796, -0.6460178, -0.4440648, -0.04810122, 0.4053981, 0.4947536, 
    0.3987087, 0.2702258, 0.1420681, 0.09937599, 0.05018979, 0.0904243, 
    0.1007921, 0.08306745, 0.1223578, 0.1923121, 0.1558052, 0.05079228, 
    -0.070611, -0.2740616, -0.5647516, -0.7670628, -0.7928604, -0.6653212, 
    -0.5034723, -0.3798068, -0.3030003, -0.2232477, -0.04911035, 0.1592393, 
    0.2710231, 0.2293728, 0.206505, 0.1869249, 0.2058376, 0.1937119, 
    -0.01226139, -0.2275771, -0.1976129, -0.01647693, 0.382807, 0.5746365, 
    0.6279079, 0.5051866, 0.5810328, 0.9279242, 1.086013, 1.15421, 1.103575, 
    0.7241154, 0.053738, -0.6123428, -0.8658258, -0.6526098, -0.5237845, 
    -0.2203505, -0.1844131, -0.1397353, 0.02706158, 0.1831814, 0.3654079, 
    0.4740669, 0.4624621, 0.3692817, 0.2724553, 0.2400986, 0.2555446, 
    0.2147731, 0.1560654, 0.1281195, 0.2713975, 0.5568793, 0.5515896, 
    0.6087511, 0.4462999, 0.3271267, 0.2573187, 0.01963979, -0.219032, 
    -0.2756563, -0.08130425, 0.05725366, 0.316238, 0.5603135, 0.824376, 
    1.101183, 1.353233, 1.407726, 1.267491, 1.240782, 1.160118, 0.7290474, 
    0.07263446, -0.4016819, -0.4628311, -0.5436579,
  -0.7095431, -0.7050346, -0.5626031, -0.2386449, 0.0664821, 0.243891, 
    0.3902777, 0.339936, 0.2117458, 0.06537563, -0.01172405, 0.01714969, 
    0.04682094, 0.08368611, 0.1151801, 0.1554633, 0.1538358, 0.05365682, 
    -0.0910697, -0.221555, -0.4260632, -0.5873588, -0.700396, -0.7185439, 
    -0.6293186, -0.5402724, -0.5008681, -0.5068415, -0.4849828, -0.4009658, 
    -0.2906956, -0.1902725, -0.07173404, 0.001866221, 0.09167741, 0.2029407, 
    0.2431913, 0.1566028, -0.0182671, 0.0147731, 0.184988, 0.3597276, 
    0.3780381, 0.4153103, 0.504324, 0.5894313, 0.8017849, 0.8340602, 
    0.9076278, 0.6375922, 0.09359789, -0.4247939, -0.7259983, -0.5390031, 
    -0.235829, 0.004307747, 0.006537437, -0.06004775, -0.04876816, 
    -0.02524936, 0.08866644, 0.2082466, 0.2302517, 0.231277, 0.2360785, 
    0.2940049, 0.343712, 0.3281032, 0.2931097, 0.3215277, 0.5429307, 
    0.5026801, 0.7490992, 0.6917101, 0.3629991, 0.03015435, -0.3428438, 
    -0.558534, -0.3883845, -0.3729059, -0.1824436, 0.150792, 0.2445745, 
    0.1661566, 0.2157497, 0.5921983, 1.001573, 1.086941, 0.9760525, 
    0.8235622, 0.7571234, 0.6383572, 0.4427028, 0.1745876, -0.1454645, 
    -0.4807509,
  -0.1978083, -0.3469293, -0.350445, -0.3998428, -0.263889, -0.09588772, 
    0.116173, 0.09939224, 0.04708129, -0.0276258, -0.05676007, -0.01947165, 
    0.1096137, 0.3067979, 0.5013129, 0.6070421, 0.5452908, 0.4118598, 
    0.1867298, -0.03883982, -0.2297579, -0.4214409, -0.5284884, -0.6360245, 
    -0.6619846, -0.5772353, -0.559885, -0.6071507, -0.6967666, -0.8100476, 
    -0.8401747, -0.7037815, -0.5228406, -0.3611383, -0.1829156, 0.06508261, 
    0.3025337, 0.4136014, 0.394412, 0.3133411, 0.3576933, 0.4403755, 
    0.4914821, 0.4916936, 0.3968531, 0.2623805, 0.3365016, 0.6207789, 
    0.7873644, 0.9663352, 0.6609316, 0.06990016, -0.2468804, -0.3130589, 
    -0.2036188, -0.08171123, 0.006244481, -0.03193915, -0.1460829, -0.242844, 
    -0.286301, -0.254693, -0.2025283, -0.1186253, -0.04787338, 0.0195744, 
    0.1313422, 0.2437934, 0.3327745, 0.4487576, 0.5664659, 0.7069119, 
    0.7713813, 0.702973, 0.5848252, 0.3163848, -0.03452688, -0.4038463, 
    -0.4735081, -0.298736, 0.1626572, 0.3874619, 0.2765407, -0.04162323, 
    -0.2697484, -0.2294813, 0.113292, 0.7345157, 0.9177189, 0.7403423, 
    0.4501085, 0.4277452, 0.2516872, 0.2883571, 0.1856065, -0.02907446,
  0.1186468, 0.1022081, 0.1053169, 0.1369736, 0.1817002, 0.1951605, 
    0.2712672, 0.3382269, 0.3973903, 0.3826933, 0.3602321, 0.3061305, 
    0.2483833, 0.1822699, 0.433393, 0.5612087, 0.6581652, 0.6945906, 
    0.6706643, 0.5346456, 0.2858016, -0.01408422, -0.2826225, -0.4653538, 
    -0.5166559, -0.3897841, -0.3171767, -0.4169326, -0.642486, -0.8248426, 
    -0.9195203, -0.8892795, -0.7182019, -0.5390028, -0.3856663, -0.2272028, 
    -0.1601618, -0.07692611, -0.09559473, -0.07131087, 0.002256837, 
    0.1553167, 0.296723, 0.3213651, 0.2370227, 0.08311623, -0.02466363, 
    0.01438248, 0.3237087, 0.4815699, 0.583035, 0.479031, 0.3355739, 
    0.1577095, 0.0776962, 0.08523211, 0.16671, 0.2114366, 0.06343865, 
    -0.1169976, -0.3676323, -0.5895073, -0.6370497, -0.57315, -0.3981988, 
    -0.2007055, -0.07718652, 0.02206475, 0.04659277, 0.1185004, -0.08711481, 
    -0.1207249, -0.03553605, 0.2444608, 0.354975, 0.3969345, 0.2403591, 
    0.03275847, -0.01899967, 0.04278418, 0.190766, 0.4327095, 0.4637479, 
    0.2449165, -0.03420115, -0.2162978, -0.1673558, -0.023036, 0.1987739, 
    0.3553981, 0.3020128, 0.2110298, 0.2056587, 0.2622016, 0.2066514, 
    0.1532335,
  0.2079209, 0.2422633, 0.2864692, 0.3743924, 0.4668239, 0.5505477, 
    0.6116317, 0.6382431, 0.7040471, 0.7743272, 0.7745064, 0.6335557, 
    0.4649197, 0.3298285, 0.3131293, 0.3546169, 0.4239855, 0.5071722, 
    0.5739855, 0.4470968, 0.3323996, 0.1853948, 0.002484798, -0.123866, 
    -0.1506563, -0.1387588, -0.1317926, -0.2049372, -0.3494521, -0.4932345, 
    -0.5849012, -0.6297417, -0.5854057, -0.5020237, -0.4192437, -0.2147354, 
    -0.2312067, -0.2099014, -0.3058812, -0.2866755, -0.177626, -0.1653701, 
    -0.1335342, -0.09245345, -0.0697972, -0.04437402, -0.03838444, 
    -0.01849511, 0.03827572, 0.1290146, 0.215766, 0.2381944, 0.2190213, 
    0.1894639, 0.1751899, 0.1961695, 0.2437608, 0.2824978, 0.2795192, 
    0.2032499, 0.07600367, -0.06730682, -0.1968316, -0.3798558, -0.321734, 
    -0.2308974, -0.195318, -0.2126682, -0.2282768, -0.03018129, -0.4224989, 
    -0.467437, -0.213661, -0.3231336, -0.1663629, -0.04325068, 0.02525496, 
    0.05121541, -0.001079738, 0.0509873, 0.1424098, 0.3442816, 0.2830186, 
    0.2383246, 0.08918715, -0.09032118, -0.244081, -0.2603571, -0.1747777, 
    -0.1025119, 0.1137966, 0.2035103, 0.2430121, 0.1854275, 0.1741318, 
    0.188764,
  0.1153916, 0.1520615, 0.1977972, 0.2594183, 0.3279405, 0.3835232, 
    0.4119574, 0.4720322, 0.5763617, 0.6732692, 0.7073349, 0.6925564, 
    0.6518825, 0.6267035, 0.5966579, 0.554975, 0.5311958, 0.5228136, 
    0.5054307, 0.4622343, 0.4595324, 0.4439236, 0.3970163, 0.3171659, 
    0.2110135, 0.04154742, 0.03687626, 0.0573678, -0.02266157, -0.1581596, 
    -0.2923393, -0.2192762, -0.274029, -0.305279, -0.3149958, -0.3213271, 
    -0.3343643, -0.3490289, -0.3774632, -0.4040908, -0.4187393, -0.4451715, 
    -0.4284071, -0.3518609, -0.2249891, -0.08605695, 0.01780033, 0.08158618, 
    0.1167912, 0.1414984, 0.1128363, 0.0618923, 0.01527774, -0.02389866, 
    -0.03268784, -0.01869041, 0.02030697, 0.06120866, 0.09042415, 0.09737396, 
    0.07050234, 0.04353285, 0.0328722, 0.06975365, 0.07483184, -0.3169489, 
    -0.3168348, -0.3310113, -0.3302952, -0.3308973, -0.3021213, -0.2791719, 
    -0.276877, -0.240907, -0.2031953, -0.04741764, -0.06873927, -0.03516179, 
    -0.04186751, -0.006776363, 0.1097926, 0.1633245, 0.1901311, 0.1609482, 
    0.09800875, 0.008360445, -0.0843479, -0.1437718, -0.136236, -0.1063044, 
    -0.0349502, 0.1942328, 0.1020454, 0.1471462, 0.1038681, 0.03052834,
  0.2409124, 0.2394313, 0.2465439, 0.2904893, 0.3364528, 0.3858506, 
    0.4402777, 0.4848578, 0.5163031, 0.5626408, 0.6069769, 0.65421, 
    0.6888453, 0.7030381, 0.7170519, 0.7255643, 0.7361274, 0.7378038, 
    0.7147409, 0.6807891, 0.6363064, 0.570828, 0.4835884, 0.3835722, 
    0.3143501, 0.238048, 0.1757922, 0.1226506, 0.07875422, 0.01981869, 
    -0.02669826, -0.08102767, -0.1107315, -0.1250544, -0.1384495, -0.1507868, 
    -0.1808975, -0.2342829, -0.2931533, -0.3439996, -0.3914443, -0.4248264, 
    -0.435178, -0.4283258, -0.3923069, -0.3327204, -0.2649469, -0.1857803, 
    -0.1066786, -0.05267465, -0.04090708, -0.04707569, -0.06608623, 
    -0.08368063, -0.0920465, -0.08634993, -0.05348861, -0.0159235, 
    0.02901465, 0.05028744, 0.06172949, 0.03869888, 0.001003623, -0.05483943, 
    -0.1192763, -0.156939, -0.1918999, -0.1900283, -0.1713922, -0.1429253, 
    -0.1434135, -0.3470919, -0.3689833, -0.2494196, -0.2335342, -0.1994521, 
    -0.1464411, -0.0908584, -0.04391831, -0.00596261, 0.01885831, 0.04063565, 
    0.06264091, 0.08002377, 0.0922471, 0.09656021, 0.09127051, 0.09732519, 
    0.1189072, 0.1519964, 0.1917262, 0.1917263, 0.1953883, 0.2123968, 
    0.2331813, 0.2374619,
  0.1673447, 0.1598903, 0.1536728, 0.1643011, 0.1907659, 0.2157008, 
    0.2350205, 0.2667914, 0.3083441, 0.3591254, 0.4243761, 0.4893663, 
    0.5506781, 0.6093368, 0.66448, 0.7134383, 0.7584742, 0.7826278, 
    0.7860132, 0.7725692, 0.7464461, 0.706863, 0.6644964, 0.6073513, 
    0.5510688, 0.48546, 0.419135, 0.3616644, 0.2926377, 0.2286891, 0.1713649, 
    0.1214951, 0.07281348, 0.02178809, -0.02202702, -0.05230045, -0.08363181, 
    -0.1134333, -0.1446506, -0.1752497, -0.2079645, -0.2398818, -0.2760471, 
    -0.2912164, -0.2992568, -0.3014703, -0.2958225, -0.2877009, -0.2804417, 
    -0.2761774, -0.2790419, -0.2848362, -0.2929417, -0.2953342, -0.3035048, 
    -0.3063207, -0.2907282, -0.2666885, -0.2407282, -0.2267471, -0.2044001, 
    -0.1871475, -0.1800999, -0.1747614, -0.1775935, -0.1893772, -0.1948298, 
    -0.2174046, -0.2381403, -0.255751, -0.2644912, -0.2652887, -0.2628799, 
    -0.2576553, -0.2491266, -0.2694717, -0.266249, -0.252626, -0.2400283, 
    -0.2225479, -0.1927464, -0.1612034, -0.1227594, -0.08136946, -0.04746646, 
    -0.02554265, 0.0003199875, 0.03021907, 0.05515397, 0.07357845, 
    0.09670671, 0.1093695, 0.1237087, 0.1410264, 0.1580023, 0.1691514,
  0.06060644, 0.07099056, 0.07629654, 0.08329524, 0.09797625, 0.1148871, 
    0.1333766, 0.1571885, 0.1773708, 0.2020615, 0.2388454, 0.2694443, 
    0.3016709, 0.3345973, 0.3678167, 0.394835, 0.4216253, 0.450434, 
    0.4747667, 0.4945583, 0.5019476, 0.5053819, 0.5028428, 0.4964463, 
    0.4864039, 0.4804958, 0.4633083, 0.4495387, 0.4279893, 0.407807, 
    0.3877549, 0.361404, 0.3282985, 0.2904567, 0.2611273, 0.2254502, 
    0.192361, 0.1529567, 0.1111924, 0.07227637, 0.02789161, -0.009022459, 
    -0.0585179, -0.1002659, -0.1418838, -0.1861709, -0.2206924, -0.2475804, 
    -0.2841038, -0.3202529, -0.3482152, -0.3703506, -0.390891, -0.4014867, 
    -0.4033421, -0.4067276, -0.406223, -0.4027725, -0.3921605, -0.3793838, 
    -0.3636123, -0.34107, -0.3172093, -0.3014053, -0.2779189, -0.2551162, 
    -0.2350804, -0.2218805, -0.2128148, -0.205637, -0.1944391, -0.194195, 
    -0.1923232, -0.1904515, -0.1861546, -0.1824763, -0.1748102, -0.1697484, 
    -0.1655492, -0.1608454, -0.1506566, -0.1368057, -0.1205947, -0.1029515, 
    -0.0896377, -0.0686416, -0.0557998, -0.03524316, -0.01981347, 
    -0.0008844398, 0.009792645, 0.01970476, 0.02834734, 0.03669694, 
    0.04607195, 0.05237076,
  0.4243007, 0.4060707, 0.3881021, 0.3700361, 0.3523111, 0.3354001, 
    0.3183103, 0.3016605, 0.2839026, 0.2667317, 0.2498045, 0.2317052, 
    0.2127118, 0.1927571, 0.1714678, 0.1487303, 0.1245277, 0.09850192, 
    0.07011676, 0.0386548, 0.004019737, -0.03489631, -0.07815805, -0.1253749, 
    -0.1755214, -0.2277185, -0.2814621, -0.3363776, -0.392123, -0.4474447, 
    -0.5019042, -0.5548348, -0.6056638, -0.6531415, -0.6959476, -0.7336917, 
    -0.7661304, -0.7930679, -0.8141594, -0.8290367, -0.8371429, -0.8385429, 
    -0.8333025, -0.821681, -0.8039074, -0.7813978, -0.7551765, -0.7122087, 
    -0.6732264, -0.6382809, -0.5986977, -0.5591149, -0.4915204, -0.4351239, 
    -0.3836432, -0.339828, -0.3021808, -0.2253742, -0.1875, -0.1560063, 
    -0.1204586, -0.06710625, -0.0527997, -0.005419731, 0.03567696, 
    0.07944298, 0.1249666, 0.1730299, 0.2135901, 0.2474442, 0.2892418, 
    0.3223147, 0.342432, 0.4062829, 0.3977056, 0.4368172, 0.4487958, 
    0.5183432, 0.526237, 0.5492668, 0.5626297, 0.5731606, 0.5790522, 
    0.5824375, 0.582242, 0.5790849, 0.5735509, 0.5652989, 0.5546546, 
    0.5423661, 0.5285151, 0.5127113, 0.4951818, 0.47806, 0.4605303, 0.4422359,
  0.1647296, 0.1623368, 0.1533203, 0.1433597, 0.1310382, 0.1198244, 
    0.1182942, 0.1246257, 0.1346354, 0.1458654, 0.1546381, 0.1599445, 
    0.1584308, 0.1496902, 0.1331048, 0.1132157, 0.09570241, 0.08404875, 
    0.08247018, 0.08946896, 0.1045893, 0.1229649, 0.1391271, 0.1436193, 
    0.1307449, 0.1043452, 0.06638932, 0.01573849, -0.04576874, -0.1120605, 
    -0.1785965, -0.2457685, -0.3139, -0.3812995, -0.444499, -0.4999332, 
    -0.5425129, -0.5679359, -0.5683088, -0.5487289, -0.529068, -0.4499016, 
    -0.3213873, -0.1808758, -0.09088564, 0.01551056, 0.07128859, 0.1268554, 
    0.1541014, 0.1853518, 0.1048174, 0.1462886, 0.1308916, 0.1184239, 
    0.06109953, 0.07792902, 0.04881108, 0.027978, 0.01643831, -0.0008142889, 
    -0.007096887, -0.002946734, -0.002132893, 0.0003085136, 0.01175046, 
    0.02273679, 0.04142177, 0.07255805, 0.0906896, 0.1112788, 0.1147293, 
    0.1096997, 0.1041336, 0.1055825, 0.1793947, 0.219173, 0.3048339, 
    0.3960614, 0.4411292, 0.4396491, 0.4956701, 0.44554, 0.4869626, 
    0.4547845, 0.4538569, 0.4179194, 0.3824866, 0.3404942, 0.2980795, 
    0.2578609, 0.2210937, 0.1899252, 0.1678548, 0.1553221, 0.1522131, 0.156559,
  0.101253, 0.1012211, 0.08413029, 0.08640933, 0.1059887, 0.1146965, 
    0.1058263, 0.08419544, 0.07431591, 0.08201444, 0.1058751, 0.129003, 
    0.1392736, 0.1312985, 0.1141925, 0.1027832, 0.1093421, 0.1291828, 
    0.158772, 0.1956537, 0.2312658, 0.2636551, 0.2881505, 0.2993321, 
    0.3061193, 0.2955725, 0.2438632, 0.1542472, 0.05201769, -0.03818369, 
    -0.09858441, -0.1248868, -0.1209962, -0.09830737, -0.07285166, 
    -0.06534863, -0.07319403, -0.09833956, -0.124577, -0.1307945, -0.119206, 
    -0.09026718, 0.1853027, 0.3479488, 0.3990228, 0.5170405, 0.5329257, 
    0.5396476, 0.5295401, 0.4798168, 0.3772457, 0.2343583, 0.06541276, 
    -0.09588265, -0.221078, -0.3158208, -0.3696132, -0.4221356, -0.3954756, 
    -0.3726397, -0.3082361, -0.2490726, -0.1949711, -0.1330729, -0.08328485, 
    -0.07088256, -0.07225013, -0.07893932, -0.08043671, -0.06925511, 
    -0.03624725, 0.002018452, 0.02353477, 0.07996416, 0.08806944, 0.08071232, 
    0.07273769, 0.1095371, 0.1560059, 0.1580563, 0.1912754, 0.2314609, 
    0.2128086, 0.2067704, 0.2384109, 0.2358068, 0.2395015, 0.2328444, 
    0.2061844, 0.1670406, 0.139111, 0.1087403, 0.07954121, 0.07888937, 
    0.09327793, 0.1060219,
  -0.1456384, -0.2217941, -0.2723312, -0.302621, -0.3197271, -0.3329595, 
    -0.3298995, -0.3029463, -0.2549162, -0.1893229, -0.1110678, -0.02690458, 
    0.04246426, 0.06609678, 0.04430342, 0.04378223, 0.02091455, 0.02745724, 
    0.08696222, 0.1699702, 0.2752109, 0.4166501, 0.4870276, 0.4524899, 
    0.3497714, 0.3113927, 0.3076981, 0.2555981, 0.1785481, 0.1355138, 
    0.1295726, 0.1509758, 0.1893059, 0.2390944, 0.2774732, 0.2761384, 
    0.2339021, 0.1453769, 0.02206969, -0.09619164, -0.1663737, -0.2017903, 
    -0.01749706, 0.2206054, 0.4476397, 0.6784832, 0.5423174, 0.5519526, 
    0.4524407, 0.2889478, 0.05589128, -0.2339686, -0.477035, -0.6282719, 
    -0.7153163, -0.7275721, -0.730567, -0.6608568, -0.5606127, -0.4296882, 
    -0.3033372, -0.2277674, -0.1882004, -0.16766, -0.155811, -0.1362963, 
    -0.1085782, -0.08029008, -0.04457998, -0.02936172, 0.006933212, 
    0.06370401, 0.12609, 0.1528482, 0.2062168, 0.2506833, 0.2656245, 
    0.2482095, 0.2004876, 0.1867507, 0.2004876, 0.1889803, 0.1928381, 
    0.1818029, 0.1945145, 0.2375646, 0.303629, 0.34082, 0.3755367, 0.347037, 
    0.3525059, 0.3003573, 0.2700675, 0.1822746, 0.06879807, -0.05175841,
  -0.1717448, -0.229671, -0.1814938, -0.1700521, -0.1417813, -0.1272798, 
    -0.1416016, -0.2247868, -0.1371098, -0.2279625, -0.1778979, -0.1226234, 
    -0.1065106, -0.1078944, -0.07892299, -0.03637695, 0.03538322, 0.1670241, 
    0.2551265, 0.2426913, 0.2490067, 0.2978996, 0.321044, 0.3316076, 
    0.3295242, 0.3077471, 0.2712073, 0.2518711, 0.2486162, 0.2514157, 
    0.2671545, 0.2922363, 0.3329103, 0.3537595, 0.3314128, 0.2270026, 
    0.06796837, -0.1093421, -0.3026042, -0.4726567, -0.561882, -0.5074873, 
    -0.3291674, -0.09370184, 0.1928706, 0.3402667, 0.3386064, 0.3517735, 
    0.2743807, 0.1217443, -0.08704472, -0.3295252, -0.5355312, -0.6423508, 
    -0.6419113, -0.5343267, -0.4058436, -0.251563, -0.08766326, 0.002326965, 
    0.02789664, 0.04798138, 0.01723582, 0.01555938, 0.01811469, 0.003254652, 
    -0.04694057, -0.07968783, -0.1093104, -0.09012103, -0.07657921, 
    0.01162052, 0.1845046, 0.3511064, 0.5249507, 0.5994624, 0.6504064, 
    0.5889643, 0.4859533, 0.368668, 0.2954748, 0.2342606, 0.1909499, 
    0.1734695, 0.1895177, 0.2089839, 0.2474279, 0.2607091, 0.2593256, 
    0.2673009, 0.3061194, 0.2094721, 0.1454259, 0.06282502, -0.0312345, 
    -0.1091144,
  0.2980952, 0.2665522, 0.2731601, 0.2833163, 0.3089838, 0.2813311, 
    0.2125649, 0.1661777, 0.1365232, 0.1160319, 0.04941344, -0.06487679, 
    -0.07887411, -0.06974363, -0.07594442, 0.004621983, -0.02543926, 
    0.05708027, 0.2488284, 0.3309245, 0.2498205, 0.1962072, 0.182356, 
    0.2295732, 0.2132154, 0.2024407, 0.1684074, 0.07571602, -0.0182457, 
    -0.0634284, -0.006640911, 0.09658241, 0.2113776, 0.335042, 0.3147941, 
    0.1053867, -0.2430997, -0.6114583, -0.8319826, -0.9764814, -0.9275718, 
    -0.8538899, -0.6332197, -0.4188318, -0.2005374, -0.1191733, -0.05187249, 
    -0.04711986, -0.1290207, -0.2724615, -0.4638352, -0.6739913, -0.8455896, 
    -0.9107915, -0.8369471, -0.6473638, -0.4412928, -0.2599777, -0.1356288, 
    -0.09638721, -0.08115286, -0.04270881, 0.01264596, 0.06339467, 0.1145014, 
    0.1419428, 0.163883, 0.2397944, 0.2932124, 0.3326492, 0.3656082, 
    0.4471024, 0.5664709, 0.6619787, 0.7038895, 0.6414057, 0.499967, 
    0.3378413, 0.2536128, 0.1641759, 0.07877553, 0.0954259, 0.1063797, 
    0.1283361, 0.1183751, 0.08758089, 0.07753855, 0.09729767, 0.1358068, 
    0.1640783, 0.2180659, 0.3060542, 0.3660313, 0.3601556, 0.3287266, 
    0.2871414,
  0.2397944, 0.2436844, 0.239827, 0.2311679, 0.1913244, 0.1510571, 0.1429191, 
    0.1717441, 0.2352369, 0.2889967, 0.3263016, 0.3283849, 0.2789708, 
    0.2516759, 0.2581375, 0.2188797, 0.1939614, 0.1908526, 0.1815913, 
    0.1586256, 0.09573507, 0.07389259, 0.0990715, 0.1728669, 0.1736482, 
    0.08896399, -0.005469561, -0.1270843, -0.2367034, -0.2560556, -0.2231125, 
    -0.1778978, -0.2275562, -0.2780607, -0.3263512, -0.5191245, -0.4565759, 
    -0.3898282, -0.3009605, -0.2864918, -0.3171066, -0.3541183, -0.3194666, 
    -0.2122074, -0.09628958, -0.06460012, -0.1422205, -0.3302251, -0.5089036, 
    -0.7071621, -0.941749, -1.116081, -1.298796, -1.306446, -1.13143, 
    -0.9172207, -0.6923347, -0.3883145, -0.2861498, -0.2473313, -0.1574875, 
    -0.04746142, -0.02037811, 0.07146758, 0.06927033, 0.03315379, 
    -0.04375051, -0.002295434, 0.0324702, 0.06689402, 0.08678335, 0.08264923, 
    0.2153804, 0.3290359, 0.29873, 0.2021642, 0.1746089, 0.1464025, 
    0.1216141, 0.1445145, 0.1750483, 0.155452, 0.1021642, 0.04633737, 
    0.002880394, -0.01014048, -0.01816458, -0.001742035, 0.01264599, 
    0.05478464, 0.09921824, 0.1502762, 0.1665685, 0.1581212, 0.1728836, 
    0.2040848,
  0.4434728, 0.343131, 0.2276362, 0.1847163, 0.1088048, 0.0168452, 
    -0.06126344, -0.03227586, 0.01020455, -0.008740723, -0.1108078, 
    -0.1757492, -0.2279953, -0.2121912, -0.1326991, -0.01806693, 0.0675776, 
    0.09812784, 0.08095652, 0.09197539, 0.09910446, 0.1260086, 0.1352047, 
    0.1050615, 0.05178982, -0.04436886, -0.2090337, -0.385645, -0.4858729, 
    -0.5410486, -0.5858728, -0.5601894, -0.5671555, -0.4766119, -0.3844081, 
    -0.126856, 0.02405548, 0.147851, 0.1540685, -0.049366, -0.3156579, 
    -0.4622233, -0.466032, -0.2861006, -0.1144371, -0.1511395, -0.3926756, 
    -0.7509441, -1.114193, -1.422933, -1.595557, -1.661085, -1.628826, 
    -1.486003, -1.264096, -1.09297, -0.9209969, -0.647543, -0.5243008, 
    -0.3450039, -0.2255863, -0.1852055, -0.1055017, -0.02918339, -0.03862363, 
    -0.1373053, -0.2736659, -0.3655441, -0.3440597, -0.2536463, -0.174919, 
    -0.1643071, -0.2146815, -0.3119797, -0.3837895, -0.4015955, -0.3647141, 
    -0.3057134, -0.2513677, -0.2544764, -0.2839849, -0.2366379, -0.1188482, 
    -0.1156255, -0.2012212, -0.2005213, -0.1448898, -0.08341515, -0.03466848, 
    0.01725209, 0.07438101, 0.1244136, 0.1734207, 0.2180496, 0.371549, 
    0.4682124,
  0.4236974, 0.2053545, 0.1155596, 0.009765029, -0.2179207, -0.4104174, 
    -0.650212, -0.6979656, -0.6638999, -0.739372, -0.8599286, -0.9590008, 
    -0.9532554, -0.8680179, -0.767139, -0.6896818, -0.6302578, -0.6374681, 
    -0.6860358, -0.6679694, -0.6569341, -0.6682785, -0.7804367, -0.8997727, 
    -0.9660811, -0.9882004, -1.020508, -0.9847825, -0.9815434, -1.016195, 
    -1.051726, -0.9575201, -0.6810229, -0.3163581, -0.0243659, 0.1413896, 
    0.1725259, 0.1328936, -0.07114267, -0.3398604, -0.4960618, -0.3984871, 
    -0.1698246, 0.02037764, 0.009586334, -0.2181482, -0.5675292, -1.014812, 
    -1.485807, -1.757324, -1.832292, -1.818002, -1.814567, -1.733236, 
    -1.541293, -1.415381, -1.326287, -1.088266, -0.6412444, -0.244597, 
    -0.03818411, -0.01204491, -0.04252994, -0.01458395, -0.03180403, 
    -0.1052089, -0.1625168, -0.1246587, -0.01676482, 0.06682897, 0.1146317, 
    0.06204391, -0.1464852, -0.4089037, -0.5840503, -0.5805672, -0.5387703, 
    -0.58698, -0.6311531, -0.6315763, -0.584164, -0.5409673, -0.6519701, 
    -0.8755866, -0.9318366, -0.9318202, -0.8371263, -0.7699386, -0.5599126, 
    -0.331104, -0.1572433, 0.03598582, 0.2061681, 0.3867345, 0.5605463, 
    0.6005365,
  0.1867994, 0.05460525, -0.05480218, -0.1967614, -0.4000816, -0.6166179, 
    -0.6393716, -0.4726071, -0.3249669, -0.2487144, -0.1407876, -0.0393548, 
    -0.01752949, -0.05315781, -0.1542809, -0.325212, -0.5257814, -0.7451663, 
    -0.9906745, -1.238249, -1.429965, -1.492107, -1.496225, -1.4653, 
    -1.421355, -1.387647, -1.303695, -1.149496, -1.041179, -1.000115, 
    -0.9286791, -0.772559, -0.5124681, -0.173975, 0.0300777, 0.01948309, 
    -0.06181622, -0.1183438, -0.1527352, -0.1390953, -0.0823245, 
    -0.009261131, -0.03411531, -0.05559969, -0.2072592, -0.5286288, 
    -0.8834145, -1.261637, -1.674577, -1.808512, -1.588819, -1.493246, 
    -1.599463, -1.598161, -1.429363, -1.306023, -1.319451, -1.133041, 
    -0.6397953, -0.1943854, 0.00507763, -0.07291716, -0.1585453, -0.1739099, 
    -0.1933924, -0.2590011, -0.2231125, -0.06959695, -0.01575571, 
    -0.05670619, -0.03281295, -0.04067457, -0.2211596, -0.4868171, 
    -0.5632821, -0.5381677, -0.5493004, -0.6240234, -0.6562827, -0.6978188, 
    -0.7549319, -0.7903161, -0.8317711, -0.9331219, -1.030795, -1.022494, 
    -0.9436859, -0.8602709, -0.7209967, -0.48641, -0.2527837, -0.1026047, 
    0.07060498, 0.286816, 0.4175289, 0.33706,
  -0.04085374, -0.1973147, -0.293571, -0.3628907, -0.3816898, -0.3367834, 
    -0.1265464, 0.1697102, 0.3552408, 0.3664389, 0.3397789, 0.2636881, 
    0.0643878, -0.2364097, -0.5682616, -0.8940914, -1.085075, -1.13029, 
    -1.17487, -1.253695, -1.232846, -1.144988, -1.120655, -1.151905, 
    -1.153305, -1.114161, -0.9918951, -0.8151376, -0.739112, -0.7076503, 
    -0.5982425, -0.4435713, -0.2893229, -0.1008139, 0.05091095, 0.01183271, 
    -0.1187663, -0.2083988, -0.2324553, -0.2095542, -0.1666346, -0.2104983, 
    -0.3137374, -0.3894043, -0.5292969, -0.7944334, -1.049138, -1.241292, 
    -1.375033, -1.285775, -0.9764491, -0.8598641, -1.092839, -1.27697, 
    -1.209327, -1.203093, -1.21058, -1.007374, -0.5868984, -0.167481, 
    0.03959914, -0.03185269, -0.1520839, -0.1151372, -0.03841192, 
    -0.0004236698, 0.1326818, 0.2232742, 0.1326982, 0.01455021, 0.04819286, 
    -0.0007494688, -0.2673998, -0.5154469, -0.5906415, -0.605355, -0.6453938, 
    -0.6690431, -0.6907876, -0.7214198, -0.7702963, -0.7210288, -0.6194012, 
    -0.5841959, -0.6271977, -0.6387215, -0.5910164, -0.5385098, -0.3969569, 
    -0.2027348, -0.03457081, 0.1729813, 0.3928868, 0.4560868, 0.3390456, 
    0.1552564,
  -0.08247137, -0.1406739, -0.05940795, 0.01707315, 0.01933575, 0.1072588, 
    0.3101726, 0.4798989, 0.4141765, 0.2279625, 0.082129, -0.1093102, 
    -0.513525, -0.9402018, -1.200245, -1.266553, -1.199952, -1.158154, 
    -1.161556, -1.146257, -1.057862, -0.9982269, -1.116472, -1.27977, 
    -1.267497, -1.111768, -0.9496267, -0.8290535, -0.7531743, -0.6652992, 
    -0.4623864, -0.2283044, -0.05413342, 0.08077812, 0.1241212, 0.06481075, 
    0.006494045, -0.02091503, -0.0057621, 0.03217697, -0.01954794, 
    -0.1270504, -0.2483401, -0.3872399, -0.5579104, -0.8157222, -1.057585, 
    -1.156707, -1.129835, -0.9313483, -0.6548182, -0.6840174, -0.9782394, 
    -1.148991, -1.131267, -1.139193, -1.066846, -0.766244, -0.3621262, 
    0.06966095, 0.3213699, 0.2698237, 0.1608231, 0.1971674, 0.2385575, 
    0.2642899, 0.3249344, 0.2247066, 0.001952529, -0.04751027, 0.08891535, 
    0.1321442, 0.01533127, -0.1418297, -0.3234046, -0.4756351, -0.5071287, 
    -0.5251465, -0.5134599, -0.378516, -0.2888994, -0.3034835, -0.2585289, 
    -0.2381191, -0.2831552, -0.2986987, -0.2700526, -0.2186854, -0.1253911, 
    -0.0514816, 0.04882753, 0.2302567, 0.3334956, 0.2040848, 0.05916297, 
    0.004931211,
  0.05136681, -0.006835938, -0.01126337, -0.1062012, -0.1750331, 0.02177668, 
    0.2740884, 0.2807775, 0.08878517, -0.1689782, -0.5063801, -1.039063, 
    -1.497234, -1.628125, -1.550439, -1.400488, -1.309961, -1.427165, 
    -1.487468, -1.398699, -1.318653, -1.350375, -1.417741, -1.383855, 
    -1.20586, -0.9442879, -0.7825855, -0.7117031, -0.5045085, -0.1752117, 
    0.1025226, 0.2460608, 0.2552078, 0.1954751, 0.1754556, 0.2654457, 
    0.3463864, 0.229671, 0.1048822, 0.05211592, -0.0874517, -0.1862798, 
    -0.2160974, -0.4312179, -0.7519376, -0.9753264, -0.9759448, -1.015121, 
    -0.9534512, -0.8214848, -0.6012049, -0.5447271, -0.6857589, -0.7606612, 
    -0.745671, -0.7685877, -0.6827804, -0.3180669, 0.1258621, 0.4971838, 
    0.6834143, 0.6813471, 0.67067, 0.6624995, 0.561344, 0.5078609, 0.5082841, 
    0.3607578, 0.2008457, 0.2402985, 0.4036779, 0.4279616, 0.3343585, 
    0.1012852, -0.09990239, 0.009830475, 0.1591468, -0.0538578, -0.09140611, 
    0.2046704, 0.2384269, 0.03850842, 0.03870368, 0.06642175, 0.02306271, 
    -0.0241704, -0.01718795, 0.0609858, 0.09628856, 0.1341629, 0.2125647, 
    0.2852048, 0.3222816, 0.2481115, 0.1505203, 0.1187494,
  -0.1240728, -0.2618814, -0.3590174, -0.256592, -0.01918983, 0.2024574, 
    0.1268227, -0.1412275, -0.4682136, -1.000521, -1.62697, -2.043441, 
    -1.920833, -1.521305, -1.328158, -1.276937, -1.293978, -1.365007, 
    -1.411508, -1.394629, -1.283432, -1.153207, -0.9702317, -0.6892585, 
    -0.4840176, -0.301384, -0.02534258, 0.2770499, 0.6513338, 0.798437, 
    0.6256179, 0.4414706, 0.2801588, 0.1986973, 0.3427896, 0.5127926, 
    0.5046058, 0.3104491, 0.1431479, -0.001578808, -0.1179044, -0.0168463, 
    -0.01855522, -0.4326667, -0.9125983, -1.186426, -1.212077, -1.047185, 
    -1.049268, -0.9010096, -0.467009, -0.07159881, 0.008577108, -0.1030279, 
    -0.1298183, -0.1501796, -0.1762538, 0.07521102, 0.4248204, 0.6566727, 
    0.8643061, 0.9344233, 0.8510575, 0.7178544, 0.6258786, 0.6381993, 
    0.5976396, 0.4365065, 0.2998531, 0.298779, 0.3723786, 0.466975, 
    0.5192866, 0.4893875, 0.497314, 0.8663077, 1.047379, 0.5141926, 
    0.2106273, 0.3935705, 0.3127925, 0.2648268, 0.4198562, 0.2747554, 
    0.006135464, -0.1374029, -0.1814784, -0.08689833, -0.07571661, 
    -0.0461756, 0.06214154, 0.120361, 0.1657547, 0.1879064, 0.04145455, 
    -0.09388089,
  -0.0366056, -0.1099617, -0.04721761, 0.2685541, 0.463297, 0.4731927, 
    0.3138826, 0.2064614, -0.2303548, -1.189176, -1.595606, -1.367806, 
    -1.052328, -0.8408532, -0.7521818, -0.6388355, -0.6807461, -0.7467455, 
    -0.7257167, -0.6722336, -0.3269699, 0.1089676, 0.3246577, 0.4895503, 
    0.6234532, 0.7070795, 0.7977371, 0.8579584, 0.9152176, 0.6999018, 
    0.3424473, 0.3937492, 0.5605464, 0.618196, 0.7787919, 0.7799146, 
    0.5279779, 0.2947102, 0.1840494, -0.02376342, -0.07501674, 0.07058868, 
    -0.2162929, -0.8444178, -1.122315, -1.211491, -1.257178, -1.143099, 
    -0.8879399, -0.3168788, 0.4158361, 0.7763829, 0.8029292, 0.6228674, 
    0.4978673, 0.4770177, 0.4067215, 0.5943191, 0.8399246, 0.8881668, 
    0.9667639, 0.9789058, 0.8159502, 0.5996089, 0.4402177, 0.4176263, 
    0.3293126, 0.07325816, -0.04558969, 0.09840417, 0.4541011, 0.6486971, 
    0.8278148, 1.038524, 1.032812, 1.191129, 1.273177, 0.5952302, 0.1190262, 
    0.184521, 0.3754878, 0.5260575, 0.432047, -0.1717941, -0.6282885, 
    -0.7931812, -0.7953621, -0.5041838, -0.1975428, 0.0007970333, 0.1791662, 
    0.2677892, 0.2022945, 0.08048439, 0.01967716, -0.03295958,
  -0.03476612, 0.09623972, 0.3996577, 0.6919755, 0.781803, 0.5602372, 
    0.3213537, 0.1194007, -0.344239, -1.162419, -1.127556, -0.771436, 
    -0.7455246, -0.4159998, -0.06987357, -0.08346403, -0.1678391, -0.1583338, 
    0.04780224, 0.336409, 0.6336259, 0.9121088, 0.9092767, 0.7237787, 
    0.6565748, 0.7232905, 0.7059727, 0.580403, 0.4788731, 0.3797196, 
    0.3382645, 0.4267571, 0.5210116, 0.4719234, 0.5060863, 0.4666986, 
    0.3118322, 0.2306149, 0.1455724, -0.03769583, -0.1081222, -0.3704273, 
    -0.9978684, -1.403435, -1.343832, -1.164372, -0.9056646, -0.5268885, 
    -0.1291021, 0.4985835, 1.07443, 1.163476, 1.180566, 1.087207, 0.827392, 
    0.7782059, 0.7912593, 0.8803217, 0.9895014, 0.8958979, 0.8726557, 
    0.9117508, 0.8075191, 0.5488278, 0.2747555, 0.1893058, 0.03316975, 
    -0.1337898, 0.04007149, 0.4078603, 0.8138011, 0.9683913, 1.061442, 
    1.228011, 1.154899, 1.295767, 1.393586, 0.6205237, -0.007259607, 
    0.1965164, 0.5630692, 0.387467, -0.06650472, -0.6120777, -1.120801, 
    -1.0507, -0.6024747, -0.102686, 0.2063309, 0.4200353, 0.4363602, 
    0.3789546, 0.2876948, 0.157812, 0.122021, 0.01004181,
  0.3332024, 0.436116, 0.650537, 0.8221188, 0.5907871, 0.3364415, -0.1646979, 
    -0.3783699, -0.4124028, -0.8028651, -0.5871099, -0.2621912, -0.3799646, 
    -0.1537603, 0.143782, -0.08274794, 0.008072495, 0.2719069, 0.419091, 
    0.6561841, 0.7065097, 0.6497227, 0.683821, 0.6387041, 0.5827794, 
    0.5226724, 0.3571937, 0.2339354, 0.1453941, 0.2452142, 0.3592116, 
    0.299674, 0.3610184, 0.4352697, 0.3547195, 0.2359532, 0.1293615, 
    0.1550613, 0.1801753, 0.08139598, -0.198503, -0.7715993, -0.9835939, 
    -0.7802414, -0.6119146, -0.4037603, -0.09534562, 0.1710443, 0.3675287, 
    0.685237, 0.9599441, 1.106835, 1.193017, 1.044905, 0.817008, 0.7526525, 
    0.7566076, 0.8129227, 0.8003576, 0.7407384, 0.702327, 0.6132319, 
    0.4126297, 0.2200842, -0.02604222, -0.170313, -0.2595874, -0.1926765, 
    0.2802728, 0.583235, 0.8088538, 1.008056, 1.069254, 1.254231, 1.277783, 
    1.468701, 1.151123, -0.008968592, -0.416993, 0.05948848, 0.4782872, 
    0.06603134, -0.07560301, -0.2395188, -0.6626635, -0.6897306, -0.07858121, 
    0.4354324, 0.4470047, 0.5432287, 0.5674636, 0.4860671, 0.4365227, 
    0.3376133, 0.2649734, 0.2060542,
  0.3345048, 0.3532877, 0.5721192, 0.5491858, 0.01464792, -0.1752775, 
    -0.3030281, -0.1923833, -0.1310878, -0.2983403, -0.3254077, 0.1611814, 
    0.04160094, -0.3945643, -0.1513839, 0.01048136, 0.2110834, 0.4973955, 
    0.6761553, 0.7290201, 0.6696777, 0.5936685, 0.574007, 0.4906573, 
    0.4275713, 0.3554521, 0.2053218, 0.06152296, -0.01971054, 0.01476216, 
    0.1273108, 0.1702632, 0.2933751, 0.3244457, 0.2268387, 0.2992183, 
    0.3951492, 0.3622394, 0.2924309, 0.01233649, -0.2370777, -0.4703941, 
    -0.2616212, -0.0711267, -0.07338929, -0.03336644, 0.06450129, 0.08938742, 
    0.3098626, 0.7274246, 0.8981277, 0.9688144, 1.042301, 1.077229, 1.063215, 
    0.8965814, 0.8289219, 0.8519037, 0.7409174, 0.5579911, 0.2929194, 
    0.09480743, -0.07729539, -0.1896001, -0.3167811, -0.4274421, -0.3262864, 
    -0.111524, 0.2086258, 0.4573888, 0.7303869, 0.8771317, 0.9053867, 
    1.144629, 1.13278, 1.115121, 0.7179689, -0.1669763, -0.4972175, 
    -0.03193402, 0.3012202, 0.02001905, -0.07949269, 0.05515897, -0.03510791, 
    -0.1907883, 0.01897736, 0.544612, 0.5800774, 0.4724114, 0.4871575, 
    0.4575841, 0.3328443, 0.2721674, 0.2555497, 0.2590489,
  0.3027344, 0.317627, 0.260725, -0.1099119, -0.2148768, -0.234278, 
    -0.1682785, 0.01507111, -0.0002121031, -0.03401768, -0.2799647, 
    -0.2577312, -0.1454595, -0.2188644, -0.009766102, 0.1906247, 0.4361658, 
    0.6070311, 0.817301, 0.7640302, 0.6068361, 0.629102, 0.6249838, 
    0.5791507, 0.4394207, 0.1619787, -0.09109735, -0.2500978, -0.2063966, 
    -0.03794003, 0.1209955, 0.241715, 0.4046223, 0.3419275, 0.2302076, 
    0.3415194, 0.4066892, 0.35848, 0.08067942, -0.03974628, -0.03500986, 
    0.03740215, 0.1485507, -0.07277107, -0.2143722, -0.2358239, -0.04122758, 
    0.3378904, 0.5480301, 0.8363769, 0.9662921, 0.9611326, 1.057552, 
    1.193961, 1.049901, 0.8000317, 0.7543774, 0.6580235, 0.4301102, 
    0.1937495, -0.1162114, -0.3077641, -0.4233892, -0.4625331, -0.3642909, 
    -0.285938, -0.1078944, 0.1236649, 0.3359045, 0.5441563, 0.6725578, 
    0.7640786, 0.9733393, 1.011312, 0.6954746, 0.6481762, 0.4896808, 
    0.006916821, -0.2116379, 0.003336072, 0.1731929, 0.06279242, 
    -0.007943228, 0.08422804, 0.1478348, -0.04178119, 0.1260898, 0.4732416, 
    0.4837565, 0.4394534, 0.4694176, 0.4647946, 0.3759439, 0.3819008, 
    0.4044592, 0.3726072,
  0.01448536, 0.01455069, -0.1563153, -0.2836106, -0.009570837, 0.0569331, 
    0.01777293, 0.1333165, 0.1043777, 0.03442323, -0.186801, -0.6479981, 
    -0.2574548, 0.2488935, 0.3506012, 0.3711748, 0.7517414, 0.7754564, 
    0.8412275, 0.7906575, 0.6400557, 0.4972324, 0.3353348, 0.2067051, 
    -0.02181005, -0.2535806, -0.3459797, -0.2146158, -0.02913427, 0.09305, 
    0.2224448, 0.330631, 0.2294924, 0.2018061, 0.1857905, 0.2725747, 
    0.3151689, 0.12111, -0.03195, 0.05068398, 0.02854824, -0.164176, 
    -0.1532717, -0.4628739, -0.5079265, -0.3391767, -0.02119207, 0.3176754, 
    0.4730303, 0.741683, 0.9197099, 0.9425128, 0.9604975, 0.9275057, 
    0.6857252, 0.6306471, 0.5166008, 0.272737, 0.09589791, -0.06477916, 
    -0.244369, -0.4095546, -0.4579107, -0.363412, -0.207992, -0.09322965, 
    0.03098917, 0.2853998, 0.4539869, 0.6023433, 0.7599125, 0.7768388, 
    0.8007646, 0.5524411, 0.3888836, 0.6524892, 0.5142409, 0.08860627, 
    0.05167592, 0.101855, 0.1334305, -0.01526743, -0.06988983, -0.01316783, 
    -0.07561934, -0.1475103, 0.1513023, 0.2266598, 0.1852536, 0.3414712, 
    0.3571284, 0.2732415, 0.2651522, 0.2960935, 0.2396321, 0.2006502,
  -0.229589, -0.1876626, -0.1451011, -0.02293324, -0.01157276, 0.1167312, 
    0.1021805, 0.05165958, 0.00506115, -0.07980192, -0.3115243, -0.6693692, 
    -0.1906252, 0.3428378, 0.501399, 0.6636062, 0.7735343, 0.695117, 
    0.6997066, 0.3790522, 0.1942377, 0.06230402, 0.03455353, -0.08478212, 
    -0.3296552, -0.3659177, -0.2366371, -0.03961611, 0.05105782, 
    0.0003089905, -0.05880594, 0.09210563, 0.1203122, -0.09646893, 
    -0.1436524, -0.06209326, 0.1416337, 0.04498672, -0.02070379, 0.06785536, 
    -0.2167478, -0.4757485, -0.4764485, -0.6143546, -0.5806804, -0.2342124, 
    0.1526849, 0.3896482, 0.6932943, 0.9570634, 0.9448727, 0.9290197, 
    0.8152174, 0.6732739, 0.4993156, 0.3697909, 0.09646761, -0.1073084, 
    -0.09490621, -0.1625329, -0.2501143, -0.3120446, -0.2343431, -0.04474342, 
    -0.004199743, 0.09488845, 0.2474115, 0.388037, 0.4268715, 0.4982741, 
    0.6152024, 0.4953933, 0.4531574, 0.4335446, 0.3875642, 0.2556469, 
    0.05797476, 0.01039982, 0.007746935, 0.03530216, 0.06321561, -0.01611376, 
    -0.102393, -0.22238, -0.1482263, 0.09173131, 0.3523593, 0.2637529, 
    0.227962, 0.1859703, 0.109261, 0.1477051, 0.2136717, 0.2627115, 
    0.1218586, -0.01534843,
  -0.4178715, -0.1657877, -0.1048665, 0.2152996, 0.08622992, 0.1208162, 
    0.03417897, -0.1196949, -0.2181646, -0.1745285, -0.3490074, -0.7575369, 
    -0.04571962, 0.4779286, 0.4705887, 0.5598793, 0.5428543, 0.508235, 
    0.3689938, 0.1026859, 0.06790304, -0.1101403, -0.2818198, -0.4281411, 
    -0.4983559, -0.4057617, -0.2465007, -0.2043295, -0.2978847, -0.380795, 
    -0.2748868, -0.2715011, -0.3198249, -0.3154302, -0.2214196, -0.3897953, 
    -0.2410975, -0.1985841, -0.1012213, -0.1256189, -0.8534017, -0.7595215, 
    -0.7091632, -0.7598801, -0.6237149, -0.2506838, 0.2403805, 0.4712238, 
    0.5360186, 0.5555661, 0.3939774, 0.3574538, 0.3243318, 0.3014803, 
    0.2146475, 0.04985273, 0.03279543, 0.01997018, -0.04064202, -0.06897831, 
    -0.1732104, -0.155567, -0.1127613, -0.06354189, 0.0566237, 0.1584468, 
    0.20555, 0.2373855, 0.3112302, 0.3186522, 0.2347331, 0.2069821, 
    0.1841145, 0.1524086, 0.1380696, -0.03995818, -0.03992563, 0.01673126, 
    0.07288361, 0.02397418, -0.02999723, -0.03388727, -0.137468, -0.1561692, 
    0.02053976, 0.1128578, 0.1257486, -0.121891, -0.06381798, -0.09096718, 
    -0.1544271, -0.02823925, -0.003613472, -0.1680665, -0.4053221, -0.5133619,
  -0.1450195, 0.01896119, -0.06735039, 0.2881668, 0.1241202, -0.03566146, 
    0.02937746, -0.1119962, -0.2557946, -0.3856612, -0.3341963, -0.3258305, 
    0.156023, 0.3998213, 0.3758135, 0.346777, 0.3892088, 0.3770828, 
    0.08204746, -0.0215826, -0.1612306, -0.2133307, -0.2526364, -0.280046, 
    -0.2312007, -0.2059572, -0.1873217, -0.09956098, -0.1225429, -0.4998701, 
    -0.1743655, -0.1152837, -0.1778328, -0.3514163, -0.4884119, -0.5834641, 
    -0.4141936, -0.3153327, -0.09516652, -0.09798217, -1.065821, -0.9052567, 
    -0.7768395, -0.5637863, -0.08473349, 0.3909829, 0.7744952, 0.8808099, 
    0.7981927, 0.8674308, 0.8677237, 0.845426, 0.8443679, 0.7179031, 
    0.627978, 0.4880529, 0.3687169, 0.189827, -0.03787482, -0.1326501, 
    -0.2264328, -0.1748868, -0.1309741, -0.08790755, 0.05891895, 0.077034, 
    0.1271968, 0.1395993, 0.03133059, 0.007942677, -0.003564358, -0.01544571, 
    -0.07682323, -0.1814456, 0.001855135, 0.08136338, -0.03974658, 
    -0.1248052, -0.1122563, -0.1148117, -0.04825896, -0.08312225, 0.01617789, 
    0.04134071, 0.07538986, -0.09625721, -0.09301805, -0.1087732, 
    -0.07403994, -0.2146163, -0.3022943, -0.1887374, -0.1606607, -0.4643888, 
    -0.4807463, -0.3196459,
  -0.1350427, -0.2021813, -0.3955731, -0.05918014, -0.3260747, -0.2409836, 
    -0.0715012, -0.0606125, -0.1338384, 0.02814078, -0.1735516, 0.1007967, 
    0.3013668, 0.2583504, 0.2834468, 0.2358069, 0.06770802, -0.02633476, 
    -0.1949222, -0.1674318, -0.2013516, -0.1788089, -0.2695639, -0.2568851, 
    -0.3373051, -0.3778329, -0.2786956, -0.09292042, -0.1930995, -0.4244466, 
    -0.03968155, -0.1455734, -0.1366379, -1.080648, -1.158025, -0.2545089, 
    -0.1117844, -0.06445363, -0.2880214, -0.6345873, -1.063509, -0.7409511, 
    -0.3939786, 0.008527875, 0.2654942, 0.3203608, 0.4485998, 0.535579, 
    0.5761877, 0.602034, 0.6046708, 0.6662104, 0.6848953, 0.5737299, 
    0.4795893, 0.4194005, 0.2488113, 0.1154455, 0.04684195, -0.06406301, 
    -0.1122889, -0.1921228, -0.2267257, -0.2042813, -0.2081549, -0.189909, 
    -0.2000172, -0.1743331, -0.2091801, -0.213721, -0.2315757, -0.3292975, 
    -0.3393557, -0.4860027, -0.4600102, -0.2195969, -0.03212941, -0.1011561, 
    -0.1423019, -0.1807948, -0.2421229, -0.1716151, -0.04711965, -0.2698085, 
    -0.2348313, -0.5031095, -0.340755, -0.05738974, -0.352767, -0.7021818, 
    -0.4094083, -0.2175624, -0.3927248, -0.6482265, -0.4726238, -0.2929201,
  -0.2489424, -0.3978841, -0.3901376, -0.1306646, -0.1359705, -0.1966965, 
    -0.103451, -0.08229217, -0.008822083, 0.2576654, 0.20345, 0.1588702, 
    0.3662105, 0.5443525, 0.3277006, 0.2108231, -0.0007491112, -0.3806968, 
    -0.5495934, -0.4491215, -0.3371911, -0.3256679, -0.367774, -0.2149904, 
    -0.4497561, -0.5206549, -0.02654672, -0.1085292, -1.025717, -1.094011, 
    -0.4787603, -0.08128306, -0.1299647, -1.637273, -1.489356, -0.3630377, 
    -0.008105993, -0.0452479, -0.5861177, -1.143051, -1.019711, -0.4728032, 
    -0.1832036, -0.1553553, -0.168246, -0.2211756, -0.2475591, -0.399203, 
    -0.4421392, -0.5751632, -0.7395188, -0.8108404, -0.838591, -0.7518397, 
    -0.6893885, -0.6108729, -0.4974777, -0.427816, -0.2996262, -0.2364591, 
    -0.2095873, -0.2096195, -0.09599662, -0.1440272, -0.2454429, -0.1873863, 
    -0.2387373, -0.2226892, -0.2632976, -0.3418458, -0.4042156, -0.4456871, 
    -0.4142091, -0.4116707, -0.2580897, -0.2187993, -0.3767746, -0.2791021, 
    -0.1547368, -0.06471405, -0.05984751, -0.04104869, -0.2158045, 
    -0.4432297, -0.3587407, -0.1763353, 0.07237864, -0.03642631, -0.4374352, 
    -0.5557461, -0.1624192, -0.2127285, -0.4649744, -0.3989103, -0.08359432, 
    -0.2341473,
  0.004214764, -0.1280117, 0.007714331, 0.01183218, 0.01448512, -0.0222173, 
    -0.04746142, -0.03494519, -0.1691412, -0.08295947, 0.02848232, 
    -0.01217413, 0.1273913, 0.4769526, 0.3326836, 0.07242823, -0.1217775, 
    -0.3719893, -0.3833661, -0.3514168, -0.3060226, -0.1348476, 0.06865215, 
    0.07965469, -0.3132653, -0.6344407, -0.219076, -0.1119797, -0.9720058, 
    -1.352458, -0.8914719, -0.2356776, -0.4039232, -1.069076, -1.225375, 
    -0.6676112, -0.3232428, -0.4976567, -0.8709314, -0.9671228, -0.7125819, 
    -0.3658208, -0.3250982, -0.4716964, -0.3445806, -0.1488124, -0.1052576, 
    -0.193783, -0.2075688, -0.3228358, -0.5170089, -0.6661137, -0.7833338, 
    -0.9212081, -0.9583013, -0.9707037, -0.9338383, -0.8896977, -0.7775884, 
    -0.6179692, -0.6429533, -0.7150562, -0.739063, -0.8359706, -0.9132161, 
    -0.8904135, -0.7257974, -0.7146161, -0.7824223, -0.5599775, -0.5368171, 
    -0.4686532, -0.4535165, -0.3696785, 0.04003835, -0.0003911406, 
    -0.4787929, -0.2858729, 0.01290639, -0.1175135, -0.4390305, -0.3700851, 
    -0.1786302, -0.1238286, -0.1592779, 0.06170195, 0.1813309, 0.01878208, 
    0.03928986, -0.03948618, -0.05208385, -0.1544766, -0.2827642, -0.3236175, 
    0.01964468, 0.05397069,
  0.02724552, -0.02504969, -0.04830778, -0.02517956, -0.03175509, 0.1066239, 
    0.2342442, 0.2905267, 0.02670848, -0.04895878, 0.06863558, 0.210742, 
    0.2939777, 0.5162277, 0.5557451, 0.2423029, 0.05099201, -0.1838212, 
    -0.3994634, -0.572494, -0.3893723, -0.2135751, -0.1891599, -0.1380215, 
    -0.1683273, -0.6384768, -1.019027, -0.1922531, -0.08471727, -0.7155116, 
    -0.9465663, -0.7381842, -1.060353, -0.5557458, -0.6921391, -0.9723312, 
    -0.5458336, -0.544727, -0.5967452, -0.6809087, -0.3969406, -0.1359217, 
    -0.2000005, -0.251856, -0.2410324, -0.2757981, -0.2975429, -0.1586268, 
    -0.05317426, -0.09967494, -0.1029794, -0.1522143, -0.1246264, -0.1926277, 
    -0.1847339, -0.2372078, -0.3430183, -0.3812017, -0.4196945, -0.3994798, 
    -0.4241704, -0.6882329, -0.958643, -1.091732, -1.302214, -1.460336, 
    -1.195036, -1.188314, -1.331999, -1.17142, -0.9168299, -0.2751144, 
    -0.2391118, -0.4202642, -0.194369, -0.2886888, -0.4496425, -0.585043, 
    -0.6902025, -0.5710943, -0.7462893, -0.5765955, -0.2683274, -0.1682625, 
    -0.2185879, -0.1234708, -0.1198736, -0.03253639, 0.02971953, -0.1440272, 
    -0.2368983, -0.3441737, 0.03041935, 0.2420566, 0.3039707, 0.1464026,
  0.2627271, 0.3394361, 0.1522617, 0.128938, 0.07810819, -0.01106846, 
    -0.1863611, 0.1030433, 0.1884604, -0.08608437, -0.2358729, -0.2448899, 
    0.08826447, 0.3148432, 0.586587, 0.3776026, 0.08453751, -0.1239753, 
    -0.4678712, -0.8160653, -0.7046716, -0.5391443, -0.3894699, 0.1190586, 
    -0.03055, -0.6847973, -0.9204259, -0.3166835, -0.1151372, -0.2379889, 
    -0.5713377, -0.9752603, -1.707064, -1.036898, -0.8917003, -1.149155, 
    -0.7837244, -0.7456548, -0.529981, -0.6178065, -0.3876958, -0.1237635, 
    -0.1734055, -0.05519256, -0.09765673, -0.1962082, -0.2138841, -0.1804368, 
    -0.1515307, -0.2484384, -0.1834319, -0.2038579, -0.2631514, -0.2356775, 
    -0.1965988, -0.1491706, -0.1062994, -0.159164, -0.1792648, -0.2430503, 
    -0.1752121, -0.2141604, -0.4099617, -0.5931485, -0.9746913, -1.288054, 
    -1.071241, -0.7473801, -0.570492, -0.5183599, -0.2058111, 0.3788569, 
    -0.1118823, -0.6096842, -0.5577636, -0.5953617, -0.6123381, -0.9898443, 
    -0.8522139, -0.3260099, -0.2081876, -0.1961272, -0.15695, -0.02607465, 
    0.001611233, 0.001333952, 0.02268839, 0.1133788, 0.1162105, 0.09728146, 
    0.08863878, -0.3002771, -0.0740242, 0.3878899, 0.7213207, 0.5043774,
  0.3061841, 0.2989252, 0.3383459, 0.5275059, 0.4839676, 0.5418451, 
    0.3170567, 0.2792802, 0.429215, 0.1805499, -0.1090174, -0.2383959, 
    -0.1337085, -0.1368499, 0.5222001, 0.3776846, 0.1862783, -0.001741409, 
    -0.3782392, -0.6730797, -0.6545578, -0.4121424, -0.2606939, 0.258121, 
    0.1642914, -0.4789543, -0.2239754, -0.1189299, -0.08138084, 0.5969394, 
    0.735791, -0.1272459, -1.307015, -1.53239, -1.385239, -1.133073, 
    -0.8064946, -0.7716801, -0.5558435, -0.4982916, -0.3463546, -0.2526534, 
    -0.3047531, -0.07325898, -0.06235403, -0.2469732, -0.2514329, -0.3080735, 
    -0.3002449, -0.3904141, -0.4166512, -0.3290534, -0.325098, -0.2675946, 
    -0.2306321, -0.1895511, -0.08876967, -0.04544353, 0.06606436, 0.08403254, 
    0.1606278, 0.252295, 0.1128905, -0.1334801, -0.3466797, -0.6918623, 
    -0.956788, -0.8976892, -0.6942062, -0.2180669, 0.1008784, 0.2720372, 
    -0.226742, -0.4666184, -0.4088385, -0.4461593, -0.448552, -0.4720708, 
    -0.4331549, -0.3512865, -0.3416023, -0.2620118, -0.1914721, -0.07670903, 
    -0.02335644, -0.03222704, -0.03235674, 0.01625967, 0.1194172, 0.1814451, 
    0.3283849, 0.1619949, -0.07407284, 0.004133224, 0.6970046, 0.839371,
  0.2233393, -0.09895888, -0.4372241, -0.3039069, -0.1791675, 0.1052895, 
    0.3494465, 0.3840656, 0.4017901, 0.6372066, 0.7331209, 0.2931147, 
    0.03691387, 0.2897291, 0.5935868, 0.2496743, -0.04178143, 0.1918283, 
    -0.2058272, -0.3119147, -0.3320482, -0.297787, -0.1814783, 0.3006505, 
    0.4447589, -0.1595218, -0.2994959, -0.08011138, 0.1865067, 0.9452302, 
    1.042237, 0.6381667, -0.00727582, -0.7676604, -1.135564, -0.985222, 
    -0.8343428, -0.8355474, -0.7807785, -0.6776373, -0.4376796, -0.3038091, 
    -0.3291835, -0.1236659, 0.04400992, -0.05074918, -0.1336594, -0.3145677, 
    -0.4113775, -0.3761561, -0.3658048, -0.3078132, -0.2344732, -0.1286466, 
    -0.01665115, -0.02928114, -0.01515341, 0.09503555, 0.1782548, 0.302897, 
    0.4225745, 0.4775882, 0.5838218, 0.4065752, 0.139811, -0.2593589, 
    -0.3877774, 0.01739858, -0.02843475, -0.2843267, -0.4061204, -0.407276, 
    0.08164012, -0.1398118, -0.2738774, -0.2459803, -0.3191899, -0.3517908, 
    -0.3677741, -0.282097, -0.2158208, -0.2097337, -0.1906583, -0.1753912, 
    -0.1090009, -0.0302577, -0.005973339, -0.02125645, -0.01001024, 
    -0.02356815, 0.06626034, 0.2308912, -0.0469892, -0.03299204, 0.4769364, 
    0.6152501,
  0.1634598, -0.007943034, -0.7417649, -0.9798671, -0.8138355, -0.702214, 
    -0.338249, 0.02771783, 0.1489744, 0.3711259, 0.438525, 0.1110833, 
    0.2264645, 0.8670888, 1.161425, 0.6746411, 0.4799962, 0.5083165, 
    -0.4532871, -0.7411139, -0.4888186, -0.3027349, 0.01031852, 0.216617, 
    0.4709468, 0.4823563, 0.1760086, 0.03227484, 0.6794751, 1.628141, 
    1.425326, 0.9834309, 0.5630852, 0.006949663, -0.6315763, -0.596794, 
    -0.4117193, -0.5771978, -0.6544276, -0.589779, -0.4135584, -0.2310876, 
    -0.1798996, -0.1411301, -0.02727915, 0.06181589, -0.03658903, -0.2505539, 
    -0.3878424, -0.4298671, -0.3582852, -0.2859708, -0.1831713, -0.1001472, 
    -0.04231858, 0.02910089, 0.05743766, 0.1494787, 0.1987953, 0.3795733, 
    0.5589843, 0.5772457, 0.8042483, 0.6221685, -0.01127958, -0.6385584, 
    -0.4550298, 0.3987949, 0.4929683, -0.05102587, -0.6680182, -0.5145513, 
    -0.05105877, -0.119727, -0.2795741, -0.2581059, -0.2354334, -0.1585291, 
    -0.1889654, -0.2765142, -0.3604172, -0.3881679, -0.2695808, -0.1453621, 
    -0.08611703, -0.08471704, -0.04855204, -0.07530928, -0.1409669, 
    -0.1320152, -0.1860352, -0.1620102, -0.1955404, -0.1376302, 0.08771086, 
    0.09425402,
  0.3205236, 0.2465164, -0.2143234, -0.68252, -0.6868006, -0.6047692, 
    -0.3411627, 0.005191565, 0.143815, 0.5078602, 0.3604321, 0.1873528, 
    0.312223, 0.4523106, 0.7539382, 1.074528, 1.363606, 1.350471, 0.3476396, 
    -0.6279631, -0.5829757, -0.1872892, -0.0211432, -0.1639979, -0.3740401, 
    0.02939415, -0.1092126, -0.2491868, 0.4594882, 1.687907, 2.08164, 
    1.689551, 1.470199, 1.250993, 0.2841146, -0.3013842, -0.06282604, 
    -0.1638514, -0.2918137, -0.3624517, -0.3061529, -0.02822304, 0.09524685, 
    0.05820262, 0.05133414, 0.2144364, 0.1717443, -0.09545949, -0.2597824, 
    -0.3458014, -0.2592291, -0.1568853, 0.02635038, 0.1756017, 0.1103671, 
    0.1582512, 0.1845858, 0.2387688, 0.293473, 0.3691239, 0.5693851, 
    0.6871905, 0.9384279, 0.7628093, 0.07281876, -0.2058923, -0.4436691, 
    -0.2672206, -0.2028325, -0.3903488, -0.2695806, -0.0267415, 0.158463, 
    0.2738765, 0.1628901, 0.0799799, -0.1868496, -0.4554044, -0.4600265, 
    -0.5406744, -0.7048671, -0.6902186, -0.6450688, -0.5151861, -0.3154629, 
    -0.1775885, -0.1017585, -0.1147137, -0.1512537, -0.1710296, -0.2319016, 
    -0.211833, -0.06739902, -0.1324711, 0.2326982, 0.3822749,
  0.7769852, 0.7831699, 0.4962234, 0.103157, -0.5470387, -0.6916182, 
    -0.5048985, -0.09441757, 0.2404132, 0.3980305, 0.2201171, 0.207845, 
    0.4670405, 0.2004715, 0.2438797, 0.4341786, 0.5231609, 0.8109531, 
    0.7475906, 0.7370763, 0.4728671, 0.1514318, 0.08775985, 0.03771108, 
    -0.2595708, -0.4541997, -0.5195317, -0.1236498, 0.595914, 0.9338372, 
    1.325927, 1.243131, 1.524951, 1.525, 0.9193847, -0.02309632, -0.07861376, 
    -0.07854915, 0.04887652, -0.0522306, -0.1681323, 0.1789055, 0.3779781, 
    0.3279943, 0.2434239, 0.1959142, 0.2211258, 0.07005173, -0.1557948, 
    -0.3324224, -0.3633957, -0.2783534, -0.02338916, 0.2013178, 0.1753088, 
    0.1917313, 0.2342604, 0.2627759, 0.2368484, 0.190527, 0.3097167, 
    0.4420567, 0.7915196, 0.9929681, 0.4905431, 0.2811844, 0.314241, 
    0.2610509, -0.1035001, -0.662077, -0.4791996, -0.167676, -0.003662348, 
    0.1929845, 0.2849439, 0.6466794, 0.6861649, 0.1285968, -0.2557454, 
    -0.6545904, -0.9121754, -1.011833, -1.067513, -0.9344079, -0.7704432, 
    -0.6425462, -0.4477059, -0.3257813, -0.2359214, -0.2112474, -0.2380538, 
    -0.1475925, -0.04397869, 0.1514311, 0.1362627, 0.5574865,
  0.1703931, 0.1912918, 0.2978836, 0.4369136, -0.3190435, -0.9481771, 
    -0.416537, -0.1425292, 0.01634097, 0.3905917, 0.2947097, 0.3354974, 
    0.4710933, -0.1071784, -0.332618, -0.0249846, 0.1665037, -0.01647139, 
    -0.01598358, 0.3263831, 0.2075516, -0.07112694, -0.007129669, 0.08759689, 
    0.2372553, 0.4110835, 0.1009109, -0.1138677, 0.1542475, 0.160644, 
    0.3049149, 0.4683426, 0.7821937, 1.070377, 1.226937, 0.6661787, 
    0.4475257, 0.01974201, -0.07529259, -0.01437187, -0.3383307, -0.2144208, 
    0.1252439, 0.3735836, 0.3772945, 0.2301099, 0.2148755, 0.1636221, 
    0.1057608, -0.01962948, -0.3322597, -0.489356, -0.3074549, 0.008088678, 
    0.2075516, 0.2529943, 0.2331212, 0.2593256, 0.1818352, 0.05608702, 
    -0.01041698, -0.06638956, 0.3685379, 1.013689, 0.6784989, 0.3264478, 
    0.00579375, 0.1351232, 0.4751625, -0.04925203, -0.6131511, -0.8030767, 
    -0.6418625, -0.3827316, -0.1178228, 0.2959954, 0.7503417, 1.019499, 
    0.807178, 0.1264648, -0.3960614, -0.7751141, -1.048585, -1.063119, 
    -1.121388, -1.098975, -0.8705083, -0.7209967, -0.5717454, -0.4490883, 
    -0.4063811, -0.4249682, -0.247314, 0.3209305, 0.7250323, 0.264827,
  -0.2037605, -0.3710129, 0.2377923, 0.4064936, -0.274203, -0.7032392, 
    -0.7955898, -0.8991054, -1.131299, -0.7452638, -0.6447921, -0.6365726, 
    -0.4786303, -0.9085941, -1.076351, -0.4458661, 0.408365, 0.3119464, 
    -0.3292158, -0.4041181, -0.4295092, -0.1934575, 0.1352859, 0.08518803, 
    -0.06770885, 0.12609, 0.08253527, -0.02972056, 0.2906571, 0.1825842, 
    -0.1144373, -0.09181362, 0.1836092, 0.543571, 0.6583986, 0.8550451, 
    0.8592935, 0.4130852, -0.01801801, -0.01402998, -0.1715989, -0.3286459, 
    -0.326905, -0.2252283, -0.09016991, 0.07932949, 0.04034781, -0.2001631, 
    -0.1911139, -0.003971815, -0.08380556, -0.3398607, -0.4596198, 
    -0.3702482, -0.0573411, 0.164534, 0.2613764, 0.3125646, 0.1452632, 
    -0.004346609, -0.239779, -0.6666675, -0.3861656, 0.159163, 0.3850093, 
    0.4087723, -0.09666383, -0.4560714, 0.01373649, 0.6747231, 0.525553, 
    -0.09293652, -0.5042484, -0.4607917, -0.2787927, -0.1459478, 0.1133946, 
    0.5862951, 1.081771, 0.9410155, 0.5000658, -0.00161171, -0.4346199, 
    -0.6463537, -0.8111815, -1.007259, -1.032586, -0.8935224, -0.7233891, 
    -0.5820158, -0.4686036, -0.648747, -1.141244, -0.4751306, 0.2880695, 
    0.3537755,
  3.20673e-005, -0.07044315, 0.04376578, -0.2998378, -0.7572597, -0.8686042, 
    -0.5337737, -0.7832201, -1.217302, -0.7791024, -0.2410812, -0.3528655, 
    -0.4787117, -0.4704596, -0.9507819, -0.5211595, 0.1707349, 0.4553382, 
    0.3517416, 0.1815424, -0.08224368, -0.2843429, -0.1091639, -0.05351615, 
    -0.06473033, -0.03502655, -0.0708013, 0.1702794, 0.5690748, 0.482812, 
    0.1176916, 0.005647302, 0.1424797, 0.2408521, 0.09806263, 0.1922524, 
    0.4640946, 0.4760089, 0.2453282, 0.1257479, 0.1101887, 0.03465128, 
    -0.1135914, -0.3284838, -0.5045741, -0.3722825, -0.2105632, -0.3535645, 
    -0.525456, -0.5681646, -0.4070318, -0.3109052, -0.3590665, -0.4311533, 
    -0.3049161, -0.07648182, 0.2314774, 0.3687496, 0.2279617, 0.188818, 
    -0.008317947, -0.6673837, -0.7883143, -0.5616376, -0.1756189, 0.336653, 
    0.4018875, -0.09983775, -0.3532231, 0.03855743, 0.2643224, 0.1714512, 
    0.03715777, -0.0654465, -0.1237961, -0.09817761, -0.02749074, 0.2133946, 
    0.3980789, 0.6983075, 0.6237299, 0.1862469, -0.1012864, -0.2525234, 
    -0.3524094, -0.3901043, -0.5042977, -0.5556645, -0.4697598, -0.4733567, 
    -0.4486171, -0.4838059, -1.158415, -1.531625, -0.7630208, 0.06129515,
  -0.367839, -0.2425461, -0.2853034, -0.4421228, -0.7047206, -0.8098151, 
    -0.4292974, -0.4107426, -0.8333504, -0.7717942, -0.2084315, 0.1953445, 
    -0.0354009, -0.6341313, -0.8176764, -0.7096034, -0.1977056, 0.1192377, 
    0.1652825, 0.1789871, 0.1400385, -0.03600311, -0.2107264, -0.2836593, 
    -0.1626309, -0.2187831, -0.3405441, -0.4824224, -0.431267, -0.2725916, 
    -0.1276861, -0.01560923, 0.02942657, 0.1263826, 0.08331656, -0.06621146, 
    -0.07472396, 0.04483962, 0.07353425, 0.01526618, 0.05589151, 0.1577632, 
    0.1702633, -0.003597736, -0.232048, -0.3638844, -0.3591478, -0.3322268, 
    -0.4391112, -0.7518232, -0.9320152, -0.836931, -0.6989582, -0.5590823, 
    -0.3229825, -0.1325529, 0.1865714, 0.4369296, 0.4098791, 0.3252436, 
    0.1068517, -0.3542812, -0.4134283, -0.4508307, -0.4188156, -0.1454757, 
    0.288834, 0.3564285, 0.2791336, 0.2664545, 0.1591792, 0.0294103, 
    0.06196237, -0.04488987, 0.005500793, 0.02472281, 0.05603796, 0.06111601, 
    0.1843092, 0.4762366, 0.4563639, 0.3243976, -0.0144372, -0.2460289, 
    -0.405664, -0.3622074, -0.3854008, -0.3930669, -0.2083335, -0.1225431, 
    -0.1283045, -0.1120773, -0.3357591, -0.885271, -1.004916, -0.7754726,
  -0.4304855, -0.2877772, -0.05612028, 0.06254832, -0.01663461, -0.201563, 
    -0.2774419, -0.3092616, -0.4546881, -0.6406745, -0.4685715, -0.130632, 
    -0.06834361, -0.3197922, -0.5249029, -0.5372075, -0.3623052, -0.07413788, 
    0.1027176, 0.1653803, 0.1356603, 0.1142085, 0.04824167, -0.1149257, 
    -0.2229334, -0.1344243, 0.002668768, -0.1181156, -0.3266934, -0.3826666, 
    -0.249154, -0.2037278, -0.2764167, -0.2542486, -0.1280602, -0.09474337, 
    -0.1605963, -0.1544113, -0.117481, 0.002066612, 0.183593, 0.1799797, 
    0.139192, 0.2090161, 0.1920077, 0.01515234, -0.102849, -0.2127774, 
    -0.3362963, -0.579639, -0.8576181, -1.03462, -1.084506, -0.9104168, 
    -0.5524421, -0.2225103, 0.1417966, 0.4545728, 0.480826, 0.3662918, 
    0.1144201, -0.1308762, -0.1733241, -0.1175624, -0.1083989, -0.1458013, 
    -0.140479, -0.1185063, -0.02863008, 0.145605, 0.1563146, 0.08844355, 
    0.0952794, 0.149023, 0.1056961, 0.06676382, 0.06425731, 0.05076447, 
    0.09975541, 0.2582514, 0.3284338, 0.4442701, 0.2770994, 0.07317781, 
    -0.2208333, -0.3101726, -0.2076006, -0.1557455, -0.03852534, 0.1702468, 
    0.30039, 0.3346348, 0.4137202, 0.3688471, 0.1017085, -0.2181971,
  0.298616, 0.1327306, -0.03956756, -0.07978567, -0.0142909, 0.01966095, 
    -0.09768927, -0.2975428, -0.3605474, -0.2634608, -0.174089, -0.2162277, 
    -0.276921, -0.3403163, -0.3356287, -0.4181971, -0.4705408, -0.2709152, 
    0.1005204, 0.3120113, 0.2103836, 0.02469025, -0.02360076, -0.1172043, 
    -0.2066903, -0.2480961, -0.2416021, -0.2827154, -0.429688, -0.36613, 
    -0.1595708, 0.07460886, 0.1133296, -0.02612358, -0.1519699, -0.1752934, 
    -0.1884608, -0.1718918, -0.0686366, 0.1473463, 0.3350904, 0.2701651, 
    0.1414216, 0.1351395, 0.3049149, 0.427213, 0.3453119, 0.1913242, 
    -0.0476079, -0.3079758, -0.5112963, -0.6539073, -0.9069998, -1.079868, 
    -0.8156583, -0.416163, -0.02950883, 0.2554518, 0.3280267, 0.2038081, 
    0.006216943, -0.09747767, -0.1021164, -0.0291509, 0.1082515, 0.18706, 
    0.149088, 0.0411616, -0.01681367, 0.04300079, 0.1311681, 0.1609695, 
    0.1456212, 0.1640783, 0.1866856, 0.1662267, 0.2288081, 0.2807449, 
    0.3248042, 0.2968582, 0.1872879, 0.1072749, 0.1971184, 0.1279125, 
    -0.1359379, -0.2968755, -0.1616211, 0.05794239, 0.2503257, 0.510644, 
    0.7399247, 0.7569817, 0.6700191, 0.6343907, 0.6108393, 0.4799637,
  0.64873, 0.6520014, 0.3194494, -0.004167169, -0.05166066, 0.06549428, 
    0.1895991, 0.08338165, -0.1425135, -0.1895025, -0.08929089, 0.01803336, 
    0.07262319, 0.1206538, 0.1616531, 0.1756668, 0.1362625, 0.1945795, 
    0.4038569, 0.6095371, 0.5849604, 0.4263016, 0.296728, 0.2115718, 
    0.1300939, 0.01940054, -0.1501144, -0.3190923, -0.4945155, -0.5258143, 
    -0.3003586, -0.08667043, 0.03771108, -0.04485727, -0.1017746, -0.1382655, 
    -0.1547695, -0.241895, -0.1612147, 0.02563426, 0.2634923, 0.3366531, 
    0.3137528, 0.2693192, 0.2502273, 0.4559728, 0.6423986, 0.5858719, 
    0.3314449, 0.03624624, -0.2092617, -0.3257656, -0.4871424, -0.6066736, 
    -0.6668792, -0.3815925, -0.1604662, 0.1118157, 0.2415845, 0.1067541, 
    0.07036054, 0.03077745, 0.0688796, 0.07120717, 0.08600211, 0.1356603, 
    0.1612788, 0.1273758, 0.1098465, 0.1410639, 0.2082352, 0.2140619, 
    -0.02358449, -0.114584, -0.05006576, 0.1642085, 0.4080073, 0.5150875, 
    0.607454, 0.5730139, 0.3469722, 0.1541499, 0.190299, 0.2337072, 
    0.1800123, 0.1259923, 0.04072189, 0.05439401, 0.09586501, 0.4038568, 
    0.784065, 0.9906569, 0.959537, 0.7221185, 0.54484, 0.63234,
  1.027815, 1.029492, 0.7686844, 0.2398758, -0.1909836, -0.3019862, 
    -0.08592173, 0.1500158, 0.1661128, 0.07618761, 0.02630156, 0.1051753, 
    0.1864904, 0.190185, 0.167838, 0.1590164, 0.1541173, 0.2303218, 
    0.3612462, 0.4857255, 0.5414546, 0.4419106, 0.2802404, 0.1066727, 
    -0.003792822, -0.05862683, -0.183871, -0.3481613, -0.537354, -0.62391, 
    -0.5225266, -0.3554204, -0.2639003, -0.2499842, -0.1908858, -0.1084315, 
    -0.07008505, -0.1744308, -0.2620936, -0.179216, 0.07555288, 0.2753738, 
    0.318782, 0.1759761, 0.1093419, 0.2178706, 0.469726, 0.4528152, 
    0.4268875, 0.2412593, 0.002798975, -0.2125494, -0.3189946, -0.2803879, 
    -0.2134448, -0.1356125, -0.02823925, 0.1528966, 0.2986974, 0.2868644, 
    0.2490878, 0.1759109, 0.09049433, 0.0629715, 0.08539987, 0.09274039, 
    0.09080353, -0.02845104, -0.2462733, -0.3446294, -0.3156418, -0.1870122, 
    -0.2570317, -0.3241053, -0.2052579, 0.01398063, 0.1750808, 0.2464024, 
    0.2035314, 0.3243973, 0.4803055, 0.3975418, 0.2653316, 0.1441401, 
    0.163297, 0.3654454, 0.4937331, 0.3505366, 0.2064122, 0.153759, 
    0.3837558, 0.8356599, 1.186295, 1.251236, 1.107796, 1.002653,
  1.459488, 1.447542, 1.150358, 0.8590326, 0.292301, -0.122738, -0.0836919, 
    -0.06551158, 0.02399039, 0.05908155, 0.04918575, 0.0598464, 0.0867182, 
    0.1055984, 0.1140295, 0.1468908, 0.230338, 0.3373204, 0.533105, 
    0.7302077, 0.873144, 0.8894854, 0.7358232, 0.5151361, 0.3349442, 
    0.1884923, 0.1070145, 0.03754832, -0.06609753, -0.1963384, -0.2068528, 
    -0.253793, -0.3118332, -0.3565109, -0.3511724, -0.2190109, -0.1674484, 
    -0.1485031, -0.2767258, -0.352328, -0.3099778, -0.2589686, -0.2442877, 
    -0.2461756, -0.1759445, -0.1218592, 0.008332834, 0.1232743, 0.1514156, 
    0.09876248, 0.04817657, -0.03867239, -0.06233776, -0.06141007, 
    -0.03043675, -0.01801801, -0.04941458, -0.09104872, -0.0603683, 
    -0.06905967, -0.06337941, -0.07472382, -0.1076503, -0.1474289, -0.131104, 
    -0.1065435, -0.08103895, -0.1101242, -0.2261724, -0.3437667, -0.4267745, 
    -0.5109707, -0.5294115, -0.4653326, -0.1053065, -0.0410974, 0.0951004, 
    0.07625282, 0.06342733, 0.2535151, 0.2090815, 0.2499344, 0.2310541, 
    -0.07981819, -0.2354172, -0.1223149, 0.1684077, 0.3870273, 0.2966628, 
    0.1530594, 0.2584956, 0.617773, 0.8694006, 1.213802, 1.40332, 1.443278,
  1.301009, 1.243505, 1.089355, 0.7943516, 0.4990717, 0.21206, 0.01966095, 
    -0.05572966, -0.0822596, -0.08681691, -0.08294332, 0.05379176, 
    0.002798915, -0.02464247, 0.1172681, 0.2609205, 0.4309561, 0.622704, 
    0.799413, 0.9393055, 1.029426, 1.061116, 1.020442, 0.921663, 0.7901038, 
    0.6362789, 0.5894364, 0.5599116, 0.4988927, 0.3877111, 0.2942704, 
    0.1612138, 0.007502675, -0.1449549, -0.2711105, -0.2724615, -0.1779628, 
    -0.1017583, -0.09007213, -0.148617, -0.2673507, -0.3849777, -0.4304042, 
    -0.4124354, -0.3387538, -0.3258957, -0.3547531, -0.2994797, -0.2158859, 
    -0.04360399, -0.005827308, 0.04801381, 0.1428217, 0.1768712, 0.1473466, 
    0.1263668, 0.1240067, 0.0974767, 0.07539012, 0.002506018, -0.02296603, 
    -0.03942108, -0.0250656, -0.03541714, -0.05001676, -0.05107474, 
    -0.004867047, 0.06362256, 0.1018875, -0.01943409, -0.1377283, -0.4112964, 
    -0.6488128, -0.3925135, -0.5893401, -0.2046229, -0.2002447, -0.09510142, 
    -0.005811065, 0.02216746, 0.1421544, 0.2708492, 0.3316725, 0.09563756, 
    -0.0831548, -0.2185064, -0.2245122, -0.1773607, -0.1074224, -0.05566454, 
    -0.1122237, 0.1081703, 0.4054682, 0.7444982, 1.078678, 1.275895,
  0.9049637, 0.9805821, 0.8864741, 0.6734044, 0.4109045, 0.1597488, 
    -0.02604216, -0.1224126, -0.1297856, -0.1004563, -0.07189178, 
    -0.06640685, -0.06318414, -0.04978895, -0.001416445, 0.242691, 0.2165034, 
    0.3460606, 0.4183915, 0.6636224, 0.7094555, 0.7679031, 0.8124832, 
    0.8635088, 0.871435, 0.8371902, 0.7696122, 0.7096837, 0.6426915, 
    0.5575354, 0.4821285, 0.3976233, 0.2951981, 0.1790848, 0.0768875, 
    0.06341095, 0.1046382, 0.1323888, 0.2334304, 0.250618, 0.0597651, 
    -0.02347058, -0.1326177, -0.2210943, -0.2576177, -0.2657069, -0.2650884, 
    -0.2523117, -0.2217453, -0.1168462, 0.03684845, 0.1785965, 0.2549637, 
    0.2763178, 0.2645828, 0.2375158, 0.2084142, 0.1897619, 0.1350581, 
    0.06741485, -0.002474427, -0.07558644, -0.1328456, -0.2428718, 
    -0.2186693, -0.1465826, -0.03810275, 0.07049102, 0.1340165, 0.02758729, 
    0.001985192, -0.188233, -0.219548, -0.5779303, -0.5593593, -0.5336269, 
    -0.313233, -0.007552624, 0.02781522, 0.08608347, 0.1392248, 0.3447098, 
    0.2072261, 0.1782547, 0.1153316, -0.01069385, -0.149675, -0.2442551, 
    -0.3322922, -0.3926111, -0.411231, -0.3597824, -0.1396001, 0.1350255, 
    0.4131343, 0.7015457,
  0.2166173, 0.3500971, 0.4424637, 0.434049, 0.3162593, 0.1199865, 
    -0.07311243, -0.1097824, -0.1722662, -0.2303391, -0.2396816, -0.1920905, 
    -0.09975648, 0.02579701, 0.09412384, 0.2312657, 0.3060541, 0.389127, 
    0.4019037, 0.4268713, 0.4653314, 0.4383621, 0.506461, 0.591829, 
    0.6260899, 0.8754879, 0.8097001, 0.768131, 0.6929845, 0.6165196, 
    0.5571285, 0.3373042, 0.2492509, 0.1581864, 0.104215, -0.003467306, 
    -0.09619193, -0.1495448, -0.1878586, -0.2092941, -0.2547531, -0.2971685, 
    -0.3260096, -0.3161301, -0.288119, -0.2407557, -0.1673345, -0.1054693, 
    -0.06515349, -0.04279022, -0.03165741, -0.025619, -0.02553764, 
    -0.0254074, -0.01126352, 0.006705225, 0.02807567, 0.04402618, 0.04492137, 
    0.02542268, -0.009717315, -0.0330897, -0.02015024, 0.003889441, 
    0.004052222, -0.1795906, -0.1541673, -0.118311, -0.1214361, -0.171664, 
    -0.222787, -0.1156906, -0.2331873, -0.314535, -0.3860519, -0.1482427, 
    -0.1680506, -0.1204269, -0.110938, -0.02672574, 0.09682566, 0.1578447, 
    0.1826818, 0.1692052, 0.1297521, 0.06839147, -0.004476428, -0.0857427, 
    -0.1580083, -0.217188, -0.2345057, -0.3404302, -0.1166508, -0.1283859, 
    -0.1001633, 0.03154246,
  0.166243, 0.1889155, 0.2479324, 0.2865718, 0.2979813, 0.2850906, 0.2407221, 
    0.3055007, 0.2598139, 0.2053381, 0.1518224, 0.1315425, 0.1436355, 
    0.1799799, 0.234228, 0.3020504, 0.383626, 0.4545569, 0.5156409, 
    0.5605302, 0.5866695, 0.6010413, 0.614648, 0.6363603, 0.639127, 
    0.7093094, 0.6793451, 0.6398432, 0.5807937, 0.5266433, 0.459521, 
    0.3721349, 0.2626622, 0.1277664, -0.02257538, -0.1682948, -0.3000982, 
    -0.4060064, -0.4758469, -0.5055994, -0.5224452, -0.5218755, -0.4986171, 
    -0.4652674, -0.4319178, -0.3863775, -0.3496424, -0.3288417, -0.3209966, 
    -0.317367, -0.313884, -0.3041997, -0.279867, -0.2389002, -0.1755213, 
    -0.1072271, -0.03370819, 0.04218699, 0.09996693, 0.1367996, 0.1451492, 
    0.1216303, 0.08946884, 0.06046498, 0.03320259, 0.00483346, -0.007878065, 
    0.02014923, 0.04477489, 0.0705561, 0.0432775, -0.2767094, -0.3409673, 
    -0.2215825, -0.2538091, -0.2591802, -0.2383957, -0.1778, -0.1308436, 
    -0.06925511, -0.01499081, 0.01783806, 0.03736931, 0.04104769, 0.04174751, 
    0.05672148, 0.07545522, 0.09635366, 0.1134923, 0.1186356, 0.1093419, 
    0.06889598, 0.0537267, 0.03831329, 0.05483348, 0.09383087,
  0.3313309, 0.3290685, 0.3400711, 0.3525874, 0.3550939, 0.3443843, 
    0.3090327, 0.2930008, 0.2805984, 0.2621251, 0.2332026, 0.2144851, 
    0.1932124, 0.1780107, 0.1735021, 0.1775222, 0.2124181, 0.2612137, 
    0.3121414, 0.3649409, 0.41276, 0.4600744, 0.4986648, 0.5377274, 0.56442, 
    0.5646479, 0.5413406, 0.5112136, 0.4890131, 0.4449702, 0.3882482, 
    0.3173009, 0.2398921, 0.1575028, 0.06645457, -0.016716, -0.09734753, 
    -0.1715825, -0.2490565, -0.3173507, -0.3710943, -0.4126958, -0.4494308, 
    -0.4697922, -0.4889653, -0.4948898, -0.4938319, -0.4850591, -0.4731613, 
    -0.4559738, -0.4348312, -0.4139165, -0.4006353, -0.3811203, -0.3499842, 
    -0.3234055, -0.2916183, -0.2675949, -0.2391281, -0.2235357, -0.2197922, 
    -0.2227544, -0.2365239, -0.2564946, -0.2647303, -0.2706385, -0.265772, 
    -0.2594244, -0.2486984, -0.2518722, -0.24655, -0.2547206, -0.2480799, 
    -0.2354009, -0.2484217, -0.2429042, -0.2262213, -0.2049484, -0.1479823, 
    -0.1045904, -0.05802459, -0.01865286, 0.02387643, 0.06583607, 0.09959257, 
    0.1308426, 0.1498042, 0.1682938, 0.2032384, 0.2542638, 0.2700678, 
    0.2689448, 0.289713, 0.3041336, 0.3185705, 0.3288244,
  0.491064, 0.4920405, 0.5004553, 0.5023595, 0.5087072, 0.5039546, 0.493782, 
    0.4810216, 0.4666336, 0.4553218, 0.4389806, 0.4229324, 0.4033686, 
    0.3838048, 0.3688797, 0.3521968, 0.3376948, 0.3183263, 0.3052404, 
    0.2988602, 0.2916987, 0.2829585, 0.2688797, 0.249381, 0.2326004, 
    0.2133947, 0.1943517, 0.1800776, 0.1589188, 0.1314123, 0.104866, 
    0.07613882, 0.0402827, -0.003890481, -0.0404302, -0.08029023, -0.1181646, 
    -0.1574549, -0.1945969, -0.229802, -0.2578456, -0.2877935, -0.3095708, 
    -0.3375005, -0.3540533, -0.3662603, -0.3738286, -0.3848312, -0.3976242, 
    -0.407813, -0.4146164, -0.4133469, -0.4072759, -0.4051926, -0.4014491, 
    -0.4093755, -0.4117517, -0.4022466, -0.3948573, -0.3875656, -0.3874842, 
    -0.3835779, -0.3820317, -0.3798507, -0.3747075, -0.3687017, -0.3611333, 
    -0.3491053, -0.3370611, -0.3277186, -0.3167486, -0.3029302, -0.278923, 
    -0.2504725, -0.2293137, -0.2035324, -0.174854, -0.1465174, -0.1120122, 
    -0.07916716, -0.04095101, -0.001188666, 0.02986601, 0.07311144, 
    0.1172358, 0.1598628, 0.200618, 0.2438146, 0.2798335, 0.3230138, 
    0.3595698, 0.3829911, 0.4051753, 0.4378576, 0.4590002, 0.4785151,
  -0.07391024, -0.0886569, -0.09814548, -0.1020031, -0.1008959, -0.09589958, 
    -0.08798933, -0.07858181, -0.06857204, -0.05805731, -0.0485034, 
    -0.04117918, -0.0360198, -0.03336573, -0.03382206, -0.03719163, 
    -0.04386473, -0.05372787, -0.06634212, -0.08131659, -0.09869921, 
    -0.1185069, -0.1410004, -0.1656586, -0.1924164, -0.2208508, -0.2506685, 
    -0.2806652, -0.3100758, -0.3375983, -0.3620772, -0.3827806, -0.3989921, 
    -0.410841, -0.4170742, -0.4195647, -0.4167976, -0.4087081, -0.3957682, 
    -0.3794613, -0.3592625, -0.3367214, -0.3122091, -0.2865582, -0.2603197, 
    -0.233058, -0.2159042, -0.1841326, -0.1576509, -0.1264324, -0.09516716, 
    -0.0441246, -0.05760145, -0.06224012, 0.002619267, -0.01101971, 
    0.01824474, 0.03834534, 0.06961203, 0.1237459, 0.1184726, 0.1624184, 
    0.2004714, 0.2284017, 0.2515297, 0.2743158, 0.2968092, 0.3188796, 
    0.3413892, 0.3543611, 0.3694005, 0.3821774, 0.3935704, 0.4003086, 
    0.3656731, 0.3810539, 0.3701653, 0.4214184, 0.3989902, 0.3947747, 
    0.3876784, 0.3780262, 0.3639469, 0.3460599, 0.3237782, 0.2965485, 
    0.2651682, 0.2299303, 0.1920397, 0.1524563, 0.1124992, 0.07273674, 
    0.03474855, 0.0009269714, -0.02867842, -0.05367947,
  -0.05869246, -0.0291028, 0.001219749, 0.03142786, 0.05869007, 0.08019114, 
    0.09415627, 0.1000485, 0.1004553, 0.09789944, 0.09013581, 0.07670808, 
    0.06046486, 0.04339123, 0.02638197, 0.01087093, -0.00237751, -0.01292455, 
    -0.02168095, -0.03175569, -0.04324645, -0.05683696, -0.07752381, 
    -0.1067393, -0.1398125, -0.1742363, -0.2076514, -0.2407234, -0.2750986, 
    -0.3109543, -0.3466153, -0.381186, -0.4153004, -0.4485688, -0.4758472, 
    -0.4931641, -0.4978371, -0.4881849, -0.4653015, -0.4395208, -0.3781748, 
    -0.3361664, -0.2740736, -0.2442074, -0.22404, -0.1744146, -0.2272472, 
    -0.2386889, -0.2457037, -0.217546, -0.203728, -0.2389007, -0.2251637, 
    -0.2396328, -0.1352718, -0.1983252, -0.1402682, -0.06368935, 
    -0.002491236, 0.09365132, 0.1977202, 0.2929024, 0.3705879, 0.413475, 
    0.428563, 0.425959, 0.3944974, 0.3478014, 0.3252593, 0.3084625, 
    0.3345041, 0.3487616, 0.3563957, 0.3810701, 0.3485346, 0.33745, 
    0.3556466, 0.3446279, 0.3553548, 0.2528801, 0.2767081, 0.2366526, 
    0.1528633, 0.1278635, 0.08258361, 0.0392732, 0.004946709, -0.02823973, 
    -0.05958748, -0.08909559, -0.1137705, -0.1302581, -0.1300139, -0.1251149, 
    -0.1089525, -0.08608484,
  -0.04983807, -0.006348133, 0.01598215, 0.03217697, 0.03053308, 0.02179217, 
    0.002668023, -0.01468211, -0.008773804, 0.01157117, 0.04010296, 
    0.06362247, 0.07374597, 0.07265615, 0.07137012, 0.07705021, 0.09438515, 
    0.1162264, 0.1298494, 0.1264473, 0.09814364, 0.04461161, -0.01219176, 
    -0.05325621, -0.07159933, -0.0691905, -0.07282031, -0.07405758, 
    -0.06552815, -0.06655335, -0.08854246, -0.1309252, -0.1976082, 
    -0.2673998, -0.3220222, -0.3581548, -0.3686857, -0.3551283, -0.3244476, 
    -0.2790208, -0.239666, -0.1642914, -0.05571318, -0.01079178, 0.04522943, 
    0.05222857, 0.0372709, 9.632111e-005, -0.05535603, -0.1137871, 
    -0.1706231, -0.1972995, -0.1804049, -0.1461112, -0.09837341, -0.03759867, 
    0.006997347, 0.09981966, 0.2090487, 0.3499181, 0.5058751, 0.6430979, 
    0.7453113, 0.8079259, 0.8237786, 0.7734526, 0.6729317, 0.5575836, 
    0.4678211, 0.4284332, 0.4372063, 0.4468098, 0.4347157, 0.4356761, 
    0.4087877, 0.3419747, 0.2938466, 0.3289375, 0.2314606, 0.1689119, 
    0.1371248, 0.09933162, 0.02148306, -0.04117942, -0.09679462, -0.1509289, 
    -0.2128594, -0.2502944, -0.2853198, -0.2822762, -0.2939625, -0.2731442, 
    -0.2280936, -0.1801929, -0.1342297, -0.08756638,
  -0.1330253, -0.1810395, -0.2098155, -0.2240082, -0.217335, -0.195802, 
    -0.1651864, -0.1227546, -0.06105137, -0.005795479, 0.03437376, 
    0.08048439, 0.130012, 0.1754384, 0.1967435, 0.2309723, 0.2324867, 
    0.1701491, 0.1045885, 0.06717002, 0.04080284, 0.004149675, -0.03307343, 
    -0.04638743, -0.02700317, 0.02324116, 0.06228721, 0.1109033, 0.1604159, 
    0.1942213, 0.1966131, 0.161799, 0.08714056, -0.01085734, -0.08567834, 
    -0.1088555, -0.0871594, -0.04498863, -0.02373123, -0.03689861, 
    -0.06736708, -0.1082525, -0.0565114, 0.01510429, 0.111181, 0.2265618, 
    0.08121681, 0.08024025, 0.03847504, -0.0131197, -0.03089321, 
    -0.004558563, 0.02809119, 0.05925977, 0.104133, 0.2151031, 0.2865875, 
    0.2775052, 0.2879219, 0.2809231, 0.3107249, 0.3286285, 0.3401356, 
    0.3936512, 0.4134264, 0.3945467, 0.3493807, 0.3194499, 0.2842927, 
    0.2803698, 0.3149405, 0.3647285, 0.4347649, 0.4861975, 0.4854002, 
    0.4860506, 0.3994946, 0.2338045, 0.06067634, 0.0856111, -0.05686998, 
    -0.09085417, -0.1178724, -0.1428233, -0.1628265, -0.1909353, -0.2321625, 
    -0.278338, -0.3200696, -0.3081553, -0.2498546, -0.150131, -0.09376693, 
    -0.05774808, -0.05628419, -0.09782028,
  -0.1063156, -0.1130047, -0.1160822, -0.07119274, -0.04795027, 0.005093575, 
    0.009977341, -0.06437397, -0.1063004, -0.162632, -0.1985846, -0.1853361, 
    -0.1354985, -0.06334734, 0.05196857, 0.2160959, 0.2569981, 0.2103677, 
    0.05929279, -0.1103041, -0.1287119, -0.1145684, -0.07692122, 
    -0.004688859, 0.06913954, 0.1943679, 0.3045721, 0.3686028, 0.4172683, 
    0.4390297, 0.4485834, 0.4186351, 0.3145335, 0.1798007, 0.02654552, 
    -0.09238338, -0.1566086, -0.1884279, -0.1994629, -0.2153983, -0.24157, 
    -0.2396326, -0.1716647, 0.0131011, 0.1738758, 0.3219719, 0.2378573, 
    0.1915519, 0.08974457, -0.003614545, -0.09070766, -0.09489048, 
    -0.03532004, 0.04718325, 0.1059072, 0.1217438, 0.05094299, -0.05377707, 
    -0.1331553, -0.1325044, -0.05294704, 0.0761708, 0.1675445, 0.2613758, 
    0.2856596, 0.2818835, 0.3202462, 0.3536121, 0.4091295, 0.4164699, 
    0.362808, 0.2482084, 0.2865386, 0.360497, 0.3543447, 0.2822417, 
    0.2470855, 0.07006735, -0.1228039, -0.288787, -0.3217298, -0.3743827, 
    -0.3828952, -0.4024912, -0.4342458, -0.4348317, -0.4365083, -0.4025564, 
    -0.3283866, -0.2227876, -0.1218764, -0.08942175, -0.05600688, -0.0357759, 
    -0.02853322, -0.07573318,
  0.2900867, 0.2242175, 0.08845913, 0.0363431, 0.06140828, 0.07937765, 
    0.1519527, 0.09005451, 0.2859864, 0.3495922, 0.290396, 0.1773751, 
    0.1540352, 0.189013, 0.2360191, 0.3618808, 0.3098783, 0.109601, 
    0.1409497, 0.08513927, 0.04662991, 0.03286004, 0.03852415, 0.08662033, 
    0.1184235, 0.1091471, 0.09506798, 0.09975433, 0.1180983, 0.1186676, 
    0.1236167, 0.1456857, 0.1212554, 0.07268906, -0.05499792, -0.1846204, 
    -0.3121104, -0.4031587, -0.4432468, -0.4012542, -0.2597828, -0.03769636, 
    0.2130523, 0.3258457, 0.1669588, 0.06516838, -0.07254291, -0.1936538, 
    -0.2882663, -0.3539236, -0.3569183, -0.2993988, -0.2257171, -0.1433115, 
    -0.0964691, -0.1038259, -0.1758637, -0.2580252, -0.2845227, -0.2013845, 
    -0.01294047, 0.2050771, 0.4031402, 0.5417633, 0.6231598, 0.7342275, 
    0.8679188, 0.9857085, 1.054166, 1.051041, 0.9514963, 0.7982574, 
    0.7179026, 0.6317535, 0.5165355, 0.3013662, -0.005307008, -0.2862803, 
    -0.4608409, -0.609376, -0.6024424, -0.6326834, -0.6240733, -0.644337, 
    -0.6532562, -0.6471853, -0.6217784, -0.553598, -0.4620453, -0.3434255, 
    -0.2425791, -0.125945, 0.02415264, 0.2049794, 0.3136707, 0.3313303,
  0.3068024, 0.09505107, -0.05079854, -0.08535272, -0.07960737, -0.02900517, 
    0.05981326, 0.1898425, 0.2714018, 0.2905589, 0.2602691, 0.1494782, 
    0.07828674, 0.1164051, 0.2404447, 0.282665, 0.2701325, 0.2604647, 
    0.252636, 0.2009592, 0.09939647, 0.01684439, -0.02492023, -0.03499484, 
    -0.0596205, -0.08180475, -0.03951979, -0.02747536, -0.02511525, 
    -0.002963424, 0.00774622, -0.006755829, -0.08797359, -0.1984386, 
    -0.3260748, -0.3061693, -0.2806976, -0.2077644, -0.2012222, -0.1755383, 
    -0.1285983, -0.1092461, -0.2008151, -0.390089, -0.6509613, -0.8719087, 
    -0.9769216, -1.037159, -1.007732, -0.9659675, -0.9093107, -0.8287932, 
    -0.8215828, -0.8406099, -0.7759778, -0.661134, -0.5360202, -0.406642, 
    -0.3141123, -0.195395, -0.01375428, 0.1677236, 0.3970368, 0.5194325, 
    0.6548005, 0.7329416, 0.8402821, 1.000943, 0.9943675, 0.9255198, 
    0.7221344, 0.5156565, 0.3729156, 0.292512, 0.1691233, -0.01098737, 
    -0.2456228, -0.4821787, -0.674822, -0.7021819, -0.7185557, -0.8346365, 
    -0.8525727, -0.8350108, -0.8080578, -0.758481, -0.6590993, -0.5551443, 
    -0.4722993, -0.3945487, -0.2546072, -0.04070741, 0.2256989, 0.4393056, 
    0.5460765, 0.488557,
  0.309667, 0.2752919, 0.2237783, 0.2387034, 0.265868, 0.3452139, 0.3565582, 
    0.2935862, 0.1812978, 0.05535376, -0.07080168, -0.1037933, -0.02952582, 
    0.1509267, 0.243749, 0.1982737, 0.121288, -0.003467828, -0.1373057, 
    -0.2923349, -0.4505219, -0.5310395, -0.4693043, -0.2808115, -0.06442159, 
    0.04150277, 0.02955616, 0.01422393, 0.07656121, 0.1714019, 0.1993642, 
    0.1584461, -0.06502396, -0.374822, -0.5165211, -0.6545583, -0.6618662, 
    -0.8162446, -1.033823, -1.283709, -1.454086, -1.722201, -1.937712, 
    -2.347868, -2.630161, -2.45713, -2.139877, -1.890332, -1.621713, 
    -1.322071, -1.096778, -0.9365079, -0.8558278, -0.853354, -0.7987641, 
    -0.6408379, -0.5501314, -0.4411144, -0.3631033, -0.4384777, -0.3335297, 
    -0.2105642, -0.0411143, 0.07464093, 0.2052072, 0.2897938, 0.2798165, 
    0.1502918, 0.003172696, -0.08255321, -0.2250499, -0.5236501, -0.7782236, 
    -0.9516287, -1.104656, -1.28423, -1.46198, -1.550473, -1.526889, 
    -1.518556, -1.452556, -1.300343, -1.129461, -1.033579, -0.9533867, 
    -0.8453299, -0.685418, -0.5179212, -0.3948091, -0.2882499, -0.1283541, 
    0.1050442, 0.3407052, 0.4319485, 0.4131173, 0.3679025,
  0.4492826, 0.4136707, 0.2166328, 0.1329904, 0.1182605, 0.04625523, 
    -0.07526171, -0.3376154, -0.5486344, -0.6721691, -0.658286, -0.5777357, 
    -0.5895194, -0.7110201, -0.9040542, -1.158742, -1.350473, -1.384262, 
    -1.332488, -1.145818, -0.8177419, -0.6811208, -0.5812185, -0.5031911, 
    -0.4530121, -0.4364756, -0.480242, -0.4793142, -0.354542, -0.09095154, 
    -0.05898539, -0.2424815, -0.582716, -0.8268567, -0.9033861, -0.8223803, 
    -0.8152678, -0.9873536, -1.304151, -1.591049, -1.715577, -1.756544, 
    -1.887403, -2.037078, -2.05669, -1.881544, -1.743034, -1.675977, 
    -1.543197, -1.283041, -1.002784, -0.8922861, -0.8898447, -0.8213224, 
    -0.5461924, -0.240724, -0.03465295, -0.03198361, -0.2394867, -0.5046397, 
    -0.6111013, -0.4709483, -0.2912282, -0.2310882, -0.2204763, -0.1479991, 
    -0.1147308, -0.1556325, -0.2259125, -0.2972667, -0.4852713, -0.7142263, 
    -0.9460948, -1.157211, -1.364194, -1.565707, -1.693702, -1.768669, 
    -1.864633, -1.945655, -1.902312, -1.708562, -1.524285, -1.430291, 
    -1.236394, -1.003435, -0.7523451, -0.5092947, -0.2878106, -0.1233249, 
    0.03844273, 0.1362128, 0.2889148, 0.3915353, 0.4548327, 0.4502265,
  0.2987943, 0.2222806, 0.09578323, 0.0235343, -0.05939198, -0.1425953, 
    -0.3260748, -0.462045, -0.4911792, -0.502003, -0.5277028, -0.6188812, 
    -0.8405931, -1.125147, -1.380144, -1.543262, -1.548455, -1.469955, 
    -1.442498, -1.436589, -1.425619, -1.349969, -1.302931, -1.340822, 
    -1.377817, -1.362371, -1.269256, -1.079461, -0.8659191, -0.706365, 
    -0.6862154, -0.8048679, -0.9392748, -0.962338, -0.8694344, -0.7815764, 
    -0.8350749, -1.089046, -1.364307, -1.487158, -1.450147, -1.409864, 
    -1.524821, -1.706381, -1.718246, -1.553972, -1.490577, -1.52116, 
    -1.417009, -1.139405, -0.9049814, -0.8899262, -0.8227549, -0.4420099, 
    0.05403519, 0.3306791, 0.3125966, 0.09680891, -0.2990734, -0.6887218, 
    -0.7755544, -0.53296, -0.2271332, -0.1293142, -0.1654795, -0.1256195, 
    0.000438435, 0.02317606, -0.1192557, -0.312094, -0.5207693, -0.702247, 
    -0.840138, -1.058367, -1.363331, -1.51548, -1.404492, -1.221289, 
    -1.151433, -1.222396, -1.186248, -1.016489, -0.8678231, -0.7557139, 
    -0.7040699, -0.6169441, -0.5323577, -0.5354664, -0.3719902, -0.1846855, 
    -0.02695429, 0.1398263, 0.1986966, 0.3210274, 0.3341296, 0.3247871,
  0.3305976, 0.3052728, 0.2430329, 0.1114414, -0.01269603, -0.1615243, 
    -0.2662282, -0.2638679, -0.2743659, -0.3976564, -0.5642581, -0.7599282, 
    -0.9764004, -1.124903, -1.182389, -1.214323, -1.240821, -1.250033, 
    -1.323341, -1.394744, -1.383367, -1.299171, -1.257162, -1.248992, 
    -1.181658, -1.040887, -0.8747734, -0.7543958, -0.6970227, -0.6873542, 
    -0.6701181, -0.6407723, -0.6140308, -0.5580249, -0.5558596, -0.7040205, 
    -0.9511886, -1.17396, -1.282943, -1.292969, -1.204867, -1.123145, 
    -1.265577, -1.50573, -1.515967, -1.309799, -1.180062, -1.128712, 
    -1.005144, -0.8208344, -0.7657398, -0.6828626, -0.426645, -0.01005971, 
    0.3029611, 0.4526519, 0.4658356, 0.2351552, -0.1648448, -0.4910329, 
    -0.5155447, -0.2947927, 0.01438701, 0.1534007, 0.105484, 0.1710765, 
    0.3363759, 0.3193187, 0.1129383, -0.1209648, -0.3960785, -0.6814303, 
    -0.9112637, -1.068181, -1.181821, -1.194824, -1.041456, -0.8748379, 
    -0.8089201, -0.8035817, -0.7561369, -0.5920248, -0.4060879, -0.2827973, 
    -0.2635911, -0.2734382, -0.2620451, -0.2411633, -0.2500339, -0.229461, 
    -0.1263033, -0.02946091, 0.05833197, 0.1885892, 0.3110664, 0.3350738,
  0.3972318, 0.3104973, 0.1725578, 0.02158117, -0.1090336, -0.1680999, 
    -0.2096195, -0.2259121, -0.3677416, -0.6170092, -0.749691, -0.7970872, 
    -0.8729331, -0.9627283, -1.048113, -1.138396, -1.225749, -1.289112, 
    -1.277312, -1.207797, -1.158627, -1.150863, -1.204167, -1.24699, 
    -1.230633, -1.141245, -1.043604, -0.992579, -0.9261076, -0.7878428, 
    -0.6136889, -0.4701993, -0.3905931, -0.3843756, -0.5215492, -0.7089524, 
    -0.7887859, -0.7818689, -0.7429695, -0.7497888, -0.7275233, -0.6785159, 
    -0.8379405, -1.136883, -1.067872, -0.7350268, -0.5059581, -0.345818, 
    -0.2366059, -0.2861014, -0.4144378, -0.3830089, -0.117986, 0.2188955, 
    0.50607, 0.7109201, 0.7312816, 0.4582021, 0.00416565, -0.3130707, 
    -0.3971853, -0.2253428, 0.0726064, 0.2109039, 0.1598623, 0.3148752, 
    0.5058259, 0.4156889, 0.2297027, 0.09002173, -0.1550794, -0.4910977, 
    -0.6958342, -0.7080903, -0.6391122, -0.6211915, -0.5755053, -0.4603353, 
    -0.3046558, -0.1710947, -0.1100104, -1.66893e-005, 0.1283364, 0.1358066, 
    -0.005599737, -0.1442389, -0.2117198, -0.1877291, -0.237664, -0.2958021, 
    -0.2306979, -0.09311652, 0.01070833, 0.191584, 0.3852201, 0.4512032,
  0.4518542, 0.2637689, 0.1171217, 0.04106355, -0.02451229, -0.07923245, 
    -0.1470222, -0.2244148, -0.3783212, -0.6015146, -0.7717292, -0.9634447, 
    -1.18099, -1.352947, -1.435157, -1.412729, -1.351873, -1.284929, 
    -1.250375, -1.204916, -1.185645, -1.274577, -1.368865, -1.357504, 
    -1.276059, -1.076156, -0.8294768, -0.6680347, -0.4773932, -0.2181649, 
    -0.01531649, 0.09365153, 0.1081374, 0.01106691, -0.1760259, -0.2646484, 
    -0.1972985, -0.2112956, -0.269743, -0.3017747, -0.3591967, -0.3291674, 
    -0.4558766, -0.7473152, -0.574806, -0.08294404, 0.2370428, 0.3676095, 
    0.0843904, -0.4029632, -0.5492035, -0.2931162, 0.05478412, 0.3539865, 
    0.5437001, 0.6204742, 0.6032216, 0.5084299, 0.3256337, 0.1657867, 
    0.1051097, 0.144872, 0.241275, 0.1878733, 0.1369781, 0.3966787, 
    0.5767402, 0.4851061, 0.54689, 0.5346665, 0.2058415, -0.1116872, 
    -0.288233, -0.3067229, -0.2661629, -0.1669114, 0.02449512, 0.1467772, 
    0.2005203, 0.2697258, 0.2759433, 0.3049309, 0.3374667, 0.2607903, 
    0.132942, -0.02366686, -0.2101738, -0.3029311, -0.3669283, -0.4006848, 
    -0.2937022, -0.1212575, 0.1012034, 0.3102365, 0.4337227, 0.5041654,
  0.6523913, 0.3644843, 0.1796541, 0.1367016, 0.03754735, -0.05439615, 
    -0.3089535, -0.6017749, -0.846225, -1.210027, -1.576791, -1.787615, 
    -1.712436, -1.463006, -1.280193, -1.121925, -1.000489, -0.9495125, 
    -1.022104, -1.172803, -1.153891, -1.11561, -1.072966, -0.8299979, 
    -0.5822278, -0.375457, -0.120509, 0.136278, 0.4900862, 0.7088201, 
    0.6523097, 0.5503728, 0.4073226, 0.307209, 0.3153801, 0.3555007, 
    0.3307934, 0.1896801, 0.1607909, 0.1310215, -0.04379988, 0.05335164, 
    0.1301097, -0.1462899, -0.1586924, 0.1887522, 0.426529, 0.3167306, 
    -0.1707204, -0.677947, -0.6051605, -0.06128031, 0.3179841, 0.4014313, 
    0.436555, 0.5981272, 0.8982575, 1.090998, 0.921809, 0.6565908, 0.5571605, 
    0.4225576, 0.3259104, 0.3730458, 0.3943509, 0.4882312, 0.517935, 
    0.5336901, 0.7661281, 0.746304, 0.4348626, 0.1610506, -0.0009284019, 
    -0.02786517, 0.04643464, 0.3451002, 0.7504878, 0.6417801, 0.2450509, 
    0.2700508, 0.2864897, 0.3467107, 0.4338689, 0.3129705, -0.02793121, 
    -0.4000176, -0.6124035, -0.6197276, -0.57129, -0.3739593, -0.06416118, 
    0.1731598, 0.3833646, 0.5827949, 0.6420722, 0.7005681,
  0.6496243, 0.5072578, 0.3592275, 0.1871083, 0.05673727, 0.04065657, 
    -0.06855571, -0.105942, -0.2918957, -0.8976246, -1.24463, -1.148536, 
    -0.8628752, -0.5517914, -0.4540048, -0.3943043, -0.3966811, -0.4899426, 
    -0.5864758, -0.6953787, -0.5545746, -0.3106129, -0.1075044, 0.2082184, 
    0.4693513, 0.6048818, 0.7325998, 0.9386547, 1.086002, 0.924885, 
    0.6638173, 0.6625638, 0.6756986, 0.6972804, 0.7855294, 0.7171381, 
    0.5417962, 0.3229322, 0.3216138, 0.310823, 0.232502, 0.3457509, 
    0.2687327, -0.08522238, -0.06417745, 0.2062978, 0.2444651, -0.03048605, 
    -0.3827159, -0.5087249, -0.2597992, 0.291291, 0.6591133, 0.6687976, 
    0.7819974, 1.114468, 1.394725, 1.363166, 1.025227, 0.7117663, 0.5583972, 
    0.3544422, 0.3446115, 0.4985827, 0.3715644, 0.3703923, 0.532111, 
    0.6928048, 0.9598296, 0.8784335, 0.5806797, 0.3339837, 0.1615064, 
    0.2488754, 0.2500476, 0.5547679, 1.07368, 0.5949857, 0.07747287, 
    0.09137267, 0.1917632, 0.2592112, 0.2282214, -0.1679703, -0.6454113, 
    -0.9317229, -0.84948, -0.5544446, -0.2615734, 0.05235875, 0.3463691, 
    0.4956696, 0.5224922, 0.6093412, 0.7939278, 0.79064,
  0.5876291, 0.553726, 0.3828764, 0.3039539, 0.3834134, 0.4469228, 0.3414047, 
    0.1886542, -0.155291, -0.8800142, -1.026157, -0.6615245, -0.4742035, 
    -0.184539, -0.08374155, -0.03549898, 0.1280262, 0.045995, -0.1254892, 
    -0.03509218, 0.1820465, 0.4061188, 0.6757802, 0.7995757, 0.6762522, 
    0.5744129, 0.6557767, 0.819172, 0.8134922, 0.6720369, 0.6779612, 
    0.7031726, 0.6534981, 0.6435534, 0.5788722, 0.4513333, 0.4320951, 
    0.360855, 0.308723, 0.2618804, 0.2254222, 0.2176419, -0.1520683, 
    -0.34227, -0.1566904, -0.034962, -0.03007922, -0.1008799, 0.01432189, 
    0.2288075, 0.5480458, 0.9444652, 1.052636, 1.003482, 1.146125, 1.320848, 
    1.336994, 1.092414, 0.7436026, 0.3833487, 0.08445549, 0.03836161, 
    0.1578763, 0.1777656, 0.1301744, 0.4749333, 0.7558252, 0.7919583, 
    1.019969, 0.9067371, 0.6234205, 0.4590154, 0.3332995, 0.3337066, 
    0.2286611, 0.7289214, 1.074934, 0.3778473, -0.1629567, -0.05986428, 
    0.2719554, 0.2599598, 0.1034981, -0.2755225, -0.6538582, -0.602361, 
    -0.2083507, 0.1541002, 0.3618152, 0.5095205, 0.4487783, 0.4298981, 
    0.470816, 0.5406728, 0.7408519, 0.6660471,
  0.6482415, 0.5934727, 0.4814117, 0.5484538, 0.545279, 0.503482, 0.2058256, 
    -0.3065767, -0.4362642, -0.7601085, -0.6459483, -0.1362804, -0.1946625, 
    -0.1626638, 0.1183746, 0.2305654, 0.3741688, 0.1899729, -0.09409308, 
    0.003465533, 0.1804187, 0.2887357, 0.5031726, 0.4659982, 0.226285, 
    0.1818676, 0.3117507, 0.5217929, 0.6335604, 0.7796869, 0.9695795, 
    0.7155264, 0.4744781, 0.4742665, 0.3358551, 0.2691233, 0.3138987, 
    0.2986642, 0.3380523, 0.2663726, 0.2494293, 0.1531563, -0.05672336, 
    0.1216135, 0.1387683, 0.0372386, 0.1816233, 0.3165517, 0.5370921, 
    0.6223622, 0.6224599, 0.7878896, 0.768342, 0.8204743, 0.9944813, 
    1.029914, 1.067789, 0.8430654, 0.5175771, 0.3119619, 0.1578114, 
    0.2053863, 0.2200835, 0.1864246, 0.3522773, 0.6517888, 0.7317694, 
    0.6229478, 0.7089015, 0.5492826, 0.4838529, 0.510676, 0.30454, 0.1957181, 
    0.3081369, 0.8530588, 0.6603513, -0.09170023, -0.3660494, -0.0974133, 
    0.4965809, 0.3791166, 0.1062813, -0.007357955, -0.3283372, -0.3466969, 
    0.1235335, 0.4318509, 0.3543935, 0.3896148, 0.353417, 0.2810534, 
    0.3599108, 0.4129544, 0.487808, 0.518472,
  0.6613765, 0.5170889, 0.5963044, 0.5856762, 0.2393545, 0.2760893, 
    0.02576381, -0.3441091, -0.1965505, -0.4130707, -0.6241877, -0.02265692, 
    -0.08455527, -0.4371755, 0.00138247, 0.2749988, 0.1423326, -0.1525407, 
    -0.2286963, -0.1209161, 0.09329319, 0.2505851, 0.186897, 0.09160066, 
    0.05040622, 0.2269037, 0.4740067, 0.6675291, 0.8159337, 0.8527169, 
    0.7030759, 0.285269, 0.1935208, 0.3189765, 0.2302396, 0.318065, 
    0.4756987, 0.5939119, 0.4748522, 0.35078, 0.3527168, 0.3302727, 
    0.2613273, 0.2428052, 0.03572512, 0.05844617, 0.278075, 0.2818021, 
    0.2910957, 0.2566068, 0.2476387, 0.5511707, 0.7012848, 0.8410308, 
    0.9733224, 0.9213856, 0.8605621, 0.5546702, 0.283137, 0.2560374, 
    0.1538076, 0.1143545, 0.1154124, 0.1755035, 0.2514474, 0.3101875, 
    0.3537096, 0.3980293, 0.4009268, 0.3525869, 0.4650055, 0.3715159, 
    0.1415024, 0.2526848, 0.403532, 0.5470858, 0.3373852, 0.08679911, 
    -0.1335139, -0.03230906, 0.5667795, 0.2135895, -0.05984819, 0.2668118, 
    0.1206043, 0.07748902, 0.2079743, 0.3610178, 0.2080554, 0.1436019, 
    0.1908519, 0.1417634, 0.1653147, 0.3180006, 0.465445, 0.5952792,
  0.5187488, 0.3905749, 0.4175615, 0.2923818, 0.1504872, -0.01811635, 
    -0.1797048, -0.2281423, -0.2314626, -0.354347, -0.605698, -0.2333503, 
    -0.06176871, 0.02659392, 0.4508131, 0.3073885, 0.0006504059, -0.1886563, 
    -0.1347175, -0.03811932, 0.1182771, 0.1887851, 0.09827423, 0.2551427, 
    0.417448, 0.4945474, 0.5168934, 0.5499992, 0.5606275, 0.4844394, 
    0.2612944, -0.05878997, 0.2060213, 0.3014965, 0.2618151, 0.4714342, 
    0.6989739, 0.7033358, 0.2895329, 0.211164, 0.3454258, 0.3026032, 
    0.1372876, -0.196013, -0.3120451, -0.1537607, 0.06375265, 0.1234369, 
    0.03024006, 0.04996586, 0.1711414, 0.3894519, 0.5424954, 0.6397611, 
    0.660676, 0.5049955, 0.3526193, 0.1926909, 0.119514, 0.04638571, 
    -0.04082143, -0.03219515, 0.07537335, 0.07740784, 0.1237783, 0.2698883, 
    0.3505849, 0.366633, 0.42412, 0.476073, 0.4643704, 0.3312819, 0.2940912, 
    0.3565269, 0.1383944, 0.09016705, 0.08609939, 0.07812397, -0.0594902, 
    0.08103716, 0.3641591, 0.08831269, 0.05525607, 0.3472481, 0.2310049, 
    0.02731019, 0.1314114, 0.3085113, 0.2378411, 0.2052727, 0.2112622, 
    0.3096998, 0.4010735, 0.5309076, 0.6049473, 0.6134601,
  0.304491, 0.2775707, 0.2986159, 0.2826982, 0.2558909, -0.06207788, 
    -0.2291677, -0.1272798, -0.2644704, -0.2999523, -0.3914241, -0.5133798, 
    -0.2721852, 0.08971286, 0.4669099, 0.08974552, -0.01017237, 0.01241827, 
    0.04858303, 0.1853347, 0.2303224, 0.1208167, 0.2185698, 0.3265128, 
    0.3523588, 0.3856759, 0.3692045, 0.4515615, 0.3940582, 0.291894, 
    0.1374183, 0.006737709, 0.03538322, 0.1535146, 0.1915681, 0.3800609, 
    0.5928383, 0.3795733, -0.05555141, 0.008690596, 0.1363435, -0.1456056, 
    -0.3215828, -0.5348153, -0.3970871, -0.1408858, -0.06041765, 0.04181242, 
    0.03435802, 0.1817214, 0.3817377, 0.5214021, 0.6277173, 0.7187655, 
    0.5004869, 0.256086, 0.09459507, -0.02089965, 0.03406441, -0.07754028, 
    -0.1035658, -0.1400239, -0.03121859, 0.06272674, 0.1182281, 0.233788, 
    0.3165514, 0.3822416, 0.3892081, 0.4045076, 0.3419914, 0.2975259, 
    0.2033191, 0.04200745, -0.143816, 0.1440263, 0.3267241, 0.0122874, 
    0.2309558, 0.2027334, 0.2420238, 0.08287674, 0.05240785, 0.08268127, 
    -0.1517754, -0.06233883, 0.4584465, 0.412288, 0.1604972, 0.294091, 
    0.3318028, 0.3855789, 0.4360507, 0.4294267, 0.3766117, 0.3615222,
  0.1680169, 0.2017078, 0.2424469, 0.261735, -0.01831156, -0.1906261, 
    -0.2221203, -0.1291025, -0.1343112, -0.2021332, -0.4378756, -0.7300463, 
    -0.4047863, 0.08800364, 0.4492507, 0.28509, 0.1475739, 0.1482258, 
    0.1575184, 0.1001458, 0.03911018, -0.01855612, 0.1338534, 0.1302891, 
    0.2136383, 0.2732897, 0.2231436, 0.2320304, 0.2007475, 0.1494946, 
    -0.07081747, -0.1765795, -0.1687346, -0.2328138, -0.1593268, -0.08239007, 
    -0.07421947, -0.274447, -0.2599461, -0.03836346, -0.163054, -0.53794, 
    -0.6181974, -0.5196133, -0.4542975, -0.2479339, -0.08396864, 0.04313064, 
    0.1534336, 0.3107901, 0.4378734, 0.5624504, 0.4822578, 0.3121732, 
    0.06004107, -0.03606904, -0.07047653, -0.1546563, -0.06824672, 
    -0.1820977, -0.2053398, -0.1668143, -0.03732228, 0.09044468, 0.09680843, 
    0.120409, 0.261539, 0.3275383, 0.2759922, 0.2959638, 0.2070789, 
    0.1453929, -0.06009197, -0.1624355, -0.4096031, -0.03011131, -0.04956156, 
    0.1472317, 0.158609, 0.2618477, 0.1014638, 0.0818674, 0.08082569, 
    0.002619267, -0.1415706, 0.1651361, 0.4625487, 0.2707028, 0.2362795, 
    0.2695313, 0.2734537, 0.271956, 0.2560058, 0.2425284, 0.2070794, 0.2158518,
  0.01238537, 0.1684885, 0.0533042, 0.1449871, -0.180486, -0.4805026, 
    -0.347739, -0.3518733, -0.3020031, -0.267791, -0.4642913, -0.7773938, 
    -0.2532401, 0.3049798, 0.3952141, 0.2377272, 0.08139515, 0.03056574, 
    -0.1556325, -0.3675461, -0.3227224, -0.2152672, -0.148243, -0.08001375, 
    0.1709628, 0.150959, 0.1523113, 0.1723795, 0.04270744, -0.2034838, 
    -0.3439298, -0.4374356, -0.4913745, -0.3644376, -0.3028655, -0.4919611, 
    -0.4325366, -0.5549164, -0.220737, -0.1536303, -0.8874846, -0.9575362, 
    -0.9634118, -0.778419, -0.7499037, -0.4338222, -0.1382332, -0.05200291, 
    0.04835534, 0.2247224, 0.3042147, 0.3455882, 0.3021469, 0.2301421, 
    0.142349, 0.008283377, -0.0822444, -0.1786634, -0.2758317, -0.3277683, 
    -0.2426772, -0.09624171, -0.01025462, -0.05813885, 0.03950119, 0.1610832, 
    0.1685214, 0.1312652, 0.0927248, -0.01365614, -0.1849937, -0.174171, 
    -0.3300142, -0.370379, -0.372396, -0.04277445, 0.03998911, 0.05123596, 
    0.162271, 0.03377151, 0.1316396, 0.1082344, 0.08100474, 0.05034053, 
    -0.00579524, 0.1814771, 0.2457347, 0.1196933, 0.1937814, 0.02311087, 
    0.09029865, 0.04566956, -0.02495193, -0.05341911, -0.05105925, -0.01167107,
  0.1348796, 0.2150545, -0.0224781, 0.1319165, -0.146746, -0.537322, 
    -0.4438489, -0.4226738, -0.3368014, -0.3694837, -0.4708664, -0.3004723, 
    0.1087885, 0.325748, 0.3403802, 0.2204089, 0.06121349, -0.1016769, 
    -0.3531256, -0.4051924, -0.399219, -0.2764654, -0.09920311, 0.008772373, 
    0.07900429, 0.01360607, -0.08442497, -0.1549325, -0.1198747, -0.5823083, 
    -0.3445315, -0.2974615, -0.328614, -0.4505379, -0.4969082, -0.6031415, 
    -0.4143236, -0.2341973, -0.0645518, -0.08971477, -1.131755, -0.9336267, 
    -0.6711104, -0.4052904, -0.1876147, 0.2541003, 0.4694815, 0.5455879, 
    0.6034167, 0.6954253, 0.7039865, 0.6053211, 0.5092925, 0.3221505, 
    0.1500151, -0.01899529, -0.1781749, -0.258725, -0.3177259, -0.2235689, 
    -0.1462903, -0.09248161, -0.04449964, 0.0145824, 0.08627868, 0.07021403, 
    0.004817009, -0.03328538, -0.1572926, -0.2294278, -0.2188482, -0.2937665, 
    -0.334343, -0.3449388, -0.2895515, 0.1230947, 0.02208558, -0.1254405, 
    -0.08898219, 0.01082256, 0.1421538, 0.1222157, 0.08268142, 0.0670886, 
    0.01790237, -0.1091316, -0.07918358, 0.001886845, -0.02335739, 
    -0.01583767, 0.08753157, -0.07542324, -0.09129286, -0.06642246, 
    0.0442543, 0.1227055,
  0.07737541, 0.0205884, -0.1565599, -0.01388466, -0.272641, -0.3359873, 
    -0.1736013, -0.1653656, -0.1612806, -0.05520892, -0.1381192, 0.0527668, 
    0.108983, 0.2242002, 0.2400546, 0.133625, -0.09651709, -0.1870122, 
    -0.2626636, -0.2534351, -0.2186041, -0.08759832, -0.03881931, 
    -0.02822351, -0.1486659, -0.2538908, -0.2576671, -0.07057399, -0.2117689, 
    -0.728435, -0.1468762, -0.1869314, -0.1388196, -1.280665, -1.225148, 
    -0.2509451, -0.06886496, -0.05716246, -0.1904632, -0.6217289, -0.9908376, 
    -0.5338876, -0.05841565, 0.210269, 0.3631986, 0.7178376, 0.8774241, 
    0.9632965, 0.9855946, 0.887206, 0.7709461, 0.6422842, 0.4442698, 
    0.2258128, 0.02633362, -0.1334971, -0.2748383, -0.3209157, -0.2931001, 
    -0.2805188, -0.2841973, -0.1869805, -0.1371269, -0.02579904, -0.07115984, 
    -0.009717464, -0.04864979, -0.140414, -0.1704435, -0.1857755, -0.2627125, 
    -0.3853197, -0.3702645, -0.5084643, -0.5142754, -0.2070811, -0.09542744, 
    -0.09482523, -0.1269704, -0.199529, -0.1424001, 0.01082253, 0.007713825, 
    -0.3767427, -0.2866547, -0.6577969, -0.4167328, 0.04983616, -0.1330733, 
    -0.2409019, -0.329021, -0.3627775, -0.3716803, -0.3250327, -0.1342616, 
    0.02949142,
  -0.1827478, -0.2271166, -0.1655288, -0.1060069, -0.1275075, -0.07810974, 
    0.03652242, -0.01403096, -0.09326261, -0.04235125, 0.1214343, 0.395751, 
    0.3769522, 0.4740372, 0.3120928, 0.1451001, -0.03405046, -0.2158046, 
    -0.1507494, -0.1630054, -0.191993, -0.2039559, -0.2792487, -0.1835127, 
    -0.3683758, -0.5817065, -0.1798352, -0.1112641, -0.8694506, -1.100587, 
    -0.2710134, -0.08522237, -0.07436626, -1.540137, -1.568182, -0.2839694, 
    0.01835835, -0.1213389, -0.4135587, -0.8903327, -0.8304858, -0.3778821, 
    -0.1169121, -0.009961963, 0.05182177, 0.1018056, -0.03029072, -0.2526378, 
    -0.4602874, -0.5750823, -0.6652682, -0.6577161, -0.6110688, -0.4313815, 
    -0.3601413, -0.3448092, -0.3275243, -0.3531427, -0.4130542, -0.3619964, 
    -0.3254726, -0.3134937, -0.2588875, -0.1325366, -0.1573088, -0.1169605, 
    -0.201726, -0.1273117, -0.09571981, -0.1253264, -0.2241218, -0.2730477, 
    -0.2365406, -0.1349943, 0.08632696, -0.1096039, -0.3940765, -0.3413911, 
    -0.1640798, -0.1238454, -0.205128, -0.2440277, -0.3026867, -0.3637871, 
    -0.2796565, -0.07954121, 0.2286127, 0.02910089, -0.4935553, -0.6948249, 
    -0.8116868, -0.8590825, -0.9963875, -0.8192713, -0.4030604, -0.3013678,
  -0.09323072, -0.1935718, -0.004737496, 0.06611225, 0.02078348, -0.08094177, 
    -0.01534933, 0.1177886, 0.1004219, -0.01920688, -0.07120895, 0.1588531, 
    0.3355947, 0.4105616, 0.223176, -0.1171398, -0.2481289, -0.2952318, 
    -0.1074231, 0.05633008, 0.06697464, 0.06315041, 0.07407236, -0.1818857, 
    -0.549561, -0.6542485, -0.1170746, -0.06097107, -0.7532885, -0.8693204, 
    -0.3423841, -0.05703226, 0.07156456, -0.7959805, -1.18755, -0.4262379, 
    -0.1529146, -0.4421887, -0.5817072, -0.634946, -0.3157889, -0.1038095, 
    -0.00296326, 0.001707971, -0.140919, -0.2230479, -0.4056325, -0.5843923, 
    -0.8066416, -0.9760753, -1.160825, -1.224106, -1.22077, -1.239389, 
    -1.261036, -1.209376, -1.234848, -1.190789, -1.260711, -1.190349, 
    -1.069434, -0.9398279, -0.7219405, -0.7573256, -0.7207856, -0.7545738, 
    -0.7690434, -0.588119, -0.7704437, -0.7227058, -0.7635586, -0.6846688, 
    -0.5398123, -0.1756525, 0.3721018, -0.01285909, -0.7914398, -0.6534678, 
    -0.1500824, -0.2208344, -0.6983899, -0.6039401, -0.3382009, -0.1237803, 
    0.003498197, 0.3255035, 0.3341135, -0.09736443, -0.3727551, -0.4021171, 
    -0.6511408, -0.6641126, -0.7907889, -0.6216805, -0.03354609, 0.01209188,
  0.08857298, -0.07615709, -0.1517916, -0.1484874, -0.1110199, -0.2507336, 
    -0.2478691, -0.03100699, -0.08527148, 0.03543174, 0.09399301, 0.08209538, 
    0.4666491, 0.5232401, 0.4059544, 0.01853657, -0.2235193, -0.2808924, 
    -0.226808, -0.1625988, 0.02495015, 0.05514169, 0.1620598, -0.1451836, 
    -0.5986657, -0.8698411, -0.7464361, -0.06001079, 0.1381823, -0.1615403, 
    -0.3597012, -0.2073412, -0.2519376, -0.2470064, -0.3877122, -0.664438, 
    -0.4658216, -0.4212415, -0.4627942, -0.5202324, -0.1388519, -0.06640726, 
    -0.03781026, -0.1214691, -0.3936045, -0.3030447, -0.25949, -0.2446789, 
    -0.3322277, -0.3962739, -0.4135265, -0.3960786, -0.4747894, -0.5847667, 
    -0.6508312, -0.5985852, -0.6124035, -0.5544608, -0.6890799, -0.8371918, 
    -1.022918, -1.024822, -0.9408867, -1.180991, -1.186248, -1.083676, 
    -1.078908, -1.011313, -0.898048, -0.9274753, -1.182749, -0.6156423, 
    -0.3246755, -0.6240573, -0.2708344, -0.3244478, -0.4115734, -0.6205903, 
    -0.7473153, -0.6424487, -0.7967947, -0.6102551, -0.3342296, -0.1538585, 
    -0.09069133, 0.0504384, 0.01830941, -0.1389334, -0.09868266, -0.04550882, 
    -0.1849947, -0.2013521, -0.1526054, -0.03955209, 0.1315579, 0.2343903,
  0.1528958, 0.08002806, 0.07029486, 0.2605782, 0.407258, 0.2432604, 
    -0.09117949, 0.1788721, 0.4159498, 0.2918122, -0.06232198, -0.338673, 
    -0.01233816, 0.2989082, 0.3358545, 0.008039474, -0.2879562, -0.3329763, 
    -0.2850592, -0.3841321, -0.39463, -0.3628755, 0.01565695, 0.007258415, 
    -0.5386076, -0.9475913, -0.8107102, -0.1544609, -0.01907682, 0.09369946, 
    0.1812329, -0.1935067, -0.9322433, -0.5815279, -0.1373544, -0.5335619, 
    -0.5545261, -0.386476, -0.3651381, -0.5573744, -0.3726575, -0.2984225, 
    -0.2217785, -0.2858247, -0.3634288, -0.3566742, -0.4603362, -0.435255, 
    -0.4104503, -0.3992362, -0.3683932, -0.2965833, -0.3278822, -0.2767105, 
    -0.2288101, -0.1232758, -0.07793069, -0.1276546, -0.1706884, -0.07905388, 
    -0.2283869, -0.5536145, -0.6582043, -0.8459158, -0.8821136, -0.6516775, 
    -0.8537119, -0.8500662, -0.1914073, -0.2755869, -0.493751, 0.1214019, 
    -0.05649513, -0.8354661, -0.7608893, -0.5949551, -0.468979, -0.8412936, 
    -0.923715, -0.5810884, -0.5522797, -0.4826998, -0.380177, -0.2469411, 
    -0.1999848, -0.03344893, 0.04051018, -0.08499432, -0.03574347, 
    0.04296744, 0.07011604, -0.125587, 0.07696819, 0.2618968, 0.1286447, 
    0.1955067,
  0.3777008, 0.3622385, 0.4485666, 0.7429351, 0.8736155, 1.020572, 0.675487, 
    0.4649727, 0.5959624, 0.2811027, -0.4016612, -0.5629569, -0.1389495, 
    0.1691231, 0.6252432, 0.1719694, -0.05478668, -0.0927577, -0.2082853, 
    -0.2640474, -0.3041026, -0.02861464, 0.5340483, 0.2361484, -0.7148447, 
    -1.002474, -0.4184585, -0.2308606, -0.4747734, 0.1955068, 0.7444, 
    0.2901359, -0.4254398, -0.6825039, -0.5634284, -0.5906258, -0.5302095, 
    -0.2588882, -0.02462685, -0.09474409, -0.147332, -0.2790215, -0.3388519, 
    -0.4399262, -0.2824392, -0.337501, -0.4935232, -0.4967297, -0.5435233, 
    -0.4809906, -0.5141288, -0.45158, -0.4182956, -0.3289237, -0.2221038, 
    -0.1266119, -0.1431649, -0.2306974, -0.2815926, -0.1660652, -0.06494212, 
    -0.149138, -0.2388518, -0.4438159, -0.5001636, -0.4109876, -0.6702648, 
    -0.7757823, -0.4207204, -0.237143, 0.0687978, 0.2969553, -0.3157237, 
    -0.5793144, -0.4985363, -0.5495616, -0.7120615, -0.6799815, -0.6512056, 
    -0.5570651, -0.529461, -0.379591, -0.2689135, -0.1672373, -0.110157, 
    -0.07368255, -0.01837635, -0.03616595, -0.006592274, -0.02184319, 
    0.2356925, 0.1415515, 0.3317533, 0.5245919, 0.479377, 0.5085437,
  0.3130521, 0.2514964, 0.03520358, -0.01614642, -0.0358572, 0.2098625, 
    0.3178701, 0.3874507, 0.5326326, 0.4998034, 0.4971342, 0.190022, 
    0.2621078, 0.6083157, 0.8548165, 0.5575347, 0.05146503, 0.01790237, 
    -0.2840664, -0.3015151, -0.3275729, -0.1534027, 0.4197091, 0.5139312, 
    0.08967996, -0.1888199, -0.2295748, -0.2421399, -0.4383962, 0.009683073, 
    0.5200671, 0.5639317, 0.6543282, 0.2833002, -0.2326667, -0.4499037, 
    -0.5726738, -0.1517754, 0.2438302, 0.3230621, 0.2586414, -0.04212368, 
    -0.1715667, -0.3501313, -0.3541026, -0.2868174, -0.2791026, -0.3689952, 
    -0.5242199, -0.4339041, -0.4342135, -0.4229505, -0.2480971, -0.04782021, 
    0.09448123, 0.1880038, 0.1631665, 0.152571, 0.1374829, 0.1785965, 
    0.2116694, 0.1950355, 0.1674314, -0.007064342, -0.08050203, -0.2280445, 
    -0.5327162, -0.3425303, -0.1849619, -0.2778819, -0.2349784, -0.2457044, 
    0.2246409, 0.03790581, -0.4360036, -0.4290375, -0.5122569, -0.5831717, 
    -0.6123872, -0.509132, -0.4951997, -0.3850925, -0.2676769, -0.2157233, 
    -0.08418036, -0.05976629, -0.02945995, -0.04926777, -0.08253717, 
    -0.2323737, -0.1989751, -0.09422302, -0.05576301, 0.3200021, 0.6197416, 
    0.5471669,
  0.008087993, -0.08393651, -0.2957855, -0.2846041, -0.2792493, -0.2758472, 
    -0.1201506, 0.3027501, 0.6317706, 0.595377, 0.5870594, 0.1520169, 
    0.4944161, 0.8777168, 0.903189, 0.8186679, 0.6417797, 0.5376129, 
    -0.1692879, -0.6322608, -0.5976415, -0.4154633, -0.006527722, 0.09461141, 
    0.006671667, 0.05244039, -0.006934613, -0.1126801, -0.2507172, 
    -0.06925553, 0.2110504, 0.3542632, 0.5449209, 0.3823719, -0.03873825, 
    0.003856182, -0.07900506, 0.05146372, 0.4228668, 0.7354318, 0.6909168, 
    0.3040028, 0.2430491, 0.04378153, -0.1110524, 0.01726787, 0.0408681, 
    -0.09381616, -0.232667, -0.3018239, -0.3363456, -0.3989106, -0.2957532, 
    -0.03492975, 0.1388659, 0.2437484, 0.2384107, 0.1923008, 0.1510899, 
    0.2577634, 0.2795243, 0.2396798, 0.3937497, 0.2816243, 0.01834297, 
    -0.2701831, -0.3165375, 0.3850575, 0.509846, 0.01103413, -0.2284515, 
    0.01204325, 0.3621244, 0.09544164, -0.1703786, -0.2153168, -0.3940765, 
    -0.3380544, -0.3953787, -0.4591481, -0.5620453, -0.5377289, -0.358237, 
    -0.2381523, -0.1272471, -0.1109059, -0.06116581, -0.1185708, -0.155014, 
    -0.2528653, -0.4994631, -0.6538916, -0.6795421, -0.4151049, 0.07880735, 
    0.1910144,
  0.1967109, 0.07809138, -0.07379659, -0.203305, -0.2983246, -0.3359706, 
    -0.3606617, 0.08790612, 0.4444332, 0.5730627, 0.4861642, 0.4203763, 
    0.5784009, 0.486588, 0.6027982, 1.204442, 1.409129, 1.119319, 0.4449375, 
    -0.1944022, -0.2157563, -0.168263, -0.1456883, -0.2169929, -0.4360361, 
    -0.07970428, -0.07946038, -0.4782722, -0.4712253, 0.09483933, 0.2512685, 
    0.1902496, 0.5650706, 0.5833486, 0.02239472, -0.02016699, 0.2589669, 
    0.2652659, 0.4765778, 1.037662, 1.15716, 0.8338044, 0.5131987, 0.2799143, 
    0.2570628, 0.3900543, 0.3801911, 0.2067047, -0.04324648, -0.1682954, 
    -0.1542979, -0.1890311, -0.08103955, 0.1698557, 0.3781236, 0.5316391, 
    0.5199533, 0.5428867, 0.4724765, 0.3798332, 0.4200516, 0.4873362, 
    0.7055168, 0.4429679, -0.0289402, -0.009115696, -0.1241709, 0.1605784, 
    0.2619292, -0.04528111, 0.05104089, 0.5701003, 0.4884431, 0.1916004, 
    0.3685049, 0.4269352, -0.151922, -0.3567884, -0.381235, -0.5885754, 
    -0.8229178, -0.7915213, -0.6441091, -0.4936535, -0.3161145, -0.1668472, 
    -0.00195384, -0.06733489, -0.1988769, -0.2725759, -0.377296, -0.3404636, 
    -0.4507008, -0.6391449, -0.3512868, 0.07664287,
  0.4481272, 0.4978668, 0.3066396, 0.06459859, -0.4402031, -0.5105639, 
    -0.5725422, 0.07914972, 0.7447424, 0.4184239, 0.1760571, 0.3012199, 
    0.2070788, -0.1677745, 0.004653931, 0.530972, 0.7951818, 0.6487787, 
    0.5259756, 0.7029288, 0.442121, -0.05981576, -0.2262383, -0.3097503, 
    -0.7498713, -0.7243991, -0.4998063, -0.9552746, -0.9021497, -0.1661306, 
    0.1031077, -0.08146274, 0.1311188, 0.4895986, 0.4269359, 0.1485177, 
    0.2402657, 0.3149401, 0.4868317, 0.9142727, 1.181445, 1.073518, 
    0.5832183, 0.1689117, 0.1021962, 0.2277985, 0.4483551, 0.3945791, 
    0.03725483, -0.05852967, -0.1031423, -0.182667, -0.02016703, 0.1850739, 
    0.3698556, 0.602782, 0.6712875, 0.6668606, 0.5262849, 0.3165197, 
    0.3081703, 0.4705882, 0.8194656, 0.6316724, 0.2063468, 0.1688465, 
    -0.04528093, -0.2976899, -0.04760814, 0.1578119, 0.2092116, 0.1341951, 
    0.1572256, 0.1551094, 0.4581205, 0.9432769, 0.7166984, 0.1275547, 
    -0.08753347, -0.4197278, -0.737534, -0.8445978, -0.8769546, -0.7387708, 
    -0.5575532, -0.3697765, -0.1310396, -0.1006522, -0.1331227, -0.2443037, 
    -0.4199557, -0.395802, -0.2698917, -0.07408905, -0.2382822, 0.02763572,
  -0.04860151, 0.04164922, 0.2514476, 0.3996409, -0.2883965, -0.8577313, 
    -0.6833827, -0.2475104, 0.4473138, 0.5016098, 0.1374667, 0.221565, 
    0.2738268, -0.1438327, -0.4347018, -0.1107926, 0.3441074, 0.2413735, 
    0.1845696, 0.3492991, 0.1803375, 0.106851, 0.2903308, 0.3587549, 
    0.1222157, 0.09376526, 0.2370106, -0.1237315, -0.6365081, -0.6196463, 
    -0.3611989, -0.2271496, -0.2314952, -0.07228303, 0.4076487, 0.5895334, 
    0.3165516, 0.174657, 0.3084464, 0.7170401, 0.8854811, 0.8504059, 
    0.5865057, 0.2494453, -0.07031381, -0.1840506, 0.1280912, 0.189859, 
    -0.08699667, -0.188722, -0.1144544, -0.13436, -0.06167114, 0.07970268, 
    0.3098459, 0.5310374, 0.6748688, 0.7337878, 0.581037, 0.2784986, 
    0.06782246, 0.1059885, 0.7283192, 0.9446931, 0.4248685, 0.2952461, 
    -0.02094847, -0.2566256, -0.04475975, 0.3457832, 0.4778643, 0.1117344, 
    -0.1048191, -0.1312511, 0.004849076, 0.4603828, 0.7202952, 0.6985505, 
    0.5109041, 0.04129171, -0.3473477, -0.6003101, -0.7687345, -0.7211108, 
    -0.6903007, -0.5289401, -0.2898285, -0.2333508, -0.2115088, -0.2805672, 
    -0.4083982, -0.4547696, -0.4266281, 0.1312819, 0.492789, 0.01521683,
  -0.3055838, -0.3121264, 0.3413562, 0.3410797, -0.3512542, -0.5350919, 
    -0.7158862, -1.032162, -0.9509447, -0.4003587, -0.2823577, -0.2875824, 
    -0.1761568, -0.5764172, -1.016358, -0.5547047, 0.2042303, 0.2372062, 
    -0.1559091, -0.2527678, -0.2001151, 0.09702042, 0.2643542, 0.2025052, 
    0.2872546, 0.3883942, 0.5159657, 0.5575023, 0.4072092, -0.0677419, 
    -0.3820159, -0.424822, -0.5632823, -0.5728851, -0.1686696, 0.2820138, 
    0.1880849, 0.04934782, 0.06347537, 0.4311841, 0.6100416, 0.6440098, 
    0.6193514, 0.5346019, 0.2101384, -0.1112484, -0.142319, -0.09397936, 
    -0.2867692, -0.4747411, -0.310353, -0.1264501, -0.1480811, -0.09907365, 
    0.2344875, 0.4709136, 0.6337066, 0.7152008, 0.5520495, 0.2866361, 
    -0.06814861, -0.4322929, 0.1262684, 0.4692864, 0.3301908, 0.2004547, 
    -0.07505012, -0.3240898, -0.389552, -0.09296942, 0.05595636, -0.06946707, 
    -0.2106616, -0.1445651, -0.0002616644, 0.1505848, 0.3074368, 0.5195137, 
    0.6017244, 0.3783193, 0.02661061, -0.3647957, -0.6693525, -0.6717782, 
    -0.5533695, -0.4113126, -0.3988452, -0.3704928, -0.2834646, -0.3604178, 
    -0.4974618, -0.6526532, -1.143181, -0.6788096, 0.1386874, 0.1734527,
  -0.01324981, 0.1729318, 0.3310372, -0.2500661, -0.8776702, -0.7181003, 
    -0.4517591, -0.9147799, -1.391131, -1.022836, -0.4216973, -0.4018241, 
    -0.2737968, -0.2896007, -0.7389661, -0.6049979, -0.07736158, 0.2762852, 
    0.2678704, 0.09962416, 0.00447464, 0.07726109, 0.1899404, 0.1551584, 
    0.04968974, -0.03429464, 0.07766825, 0.2983224, 0.439501, 0.2615712, 
    -0.008041382, -0.2280771, -0.4022148, -0.4206231, -0.2527842, 
    -0.02340627, 0.05147994, 0.002472758, 0.05987835, 0.01443553, 0.1363599, 
    0.2379551, 0.2991204, 0.2346184, 0.1620595, 0.03411317, -0.1740251, 
    -0.3070652, -0.4311373, -0.6036305, -0.4505379, -0.07726312, -0.09430408, 
    -0.147413, 0.04435134, 0.3003409, 0.5537423, 0.6988109, 0.6639964, 
    0.546711, 0.179328, -0.5197115, -0.4783216, -0.2608895, 0.00572753, 
    0.06767464, 0.03543192, -0.1291189, -0.1363942, 0.01264547, 0.04674378, 
    0.02703333, 0.05025923, 0.0430814, 0.06144094, 0.2213042, 0.3115224, 
    0.3934395, 0.3803536, 0.4353992, 0.1818514, -0.2291024, -0.5019538, 
    -0.641309, -0.6259446, -0.3500819, -0.2066412, -0.2021492, -0.1494968, 
    -0.2859384, -0.4298676, -0.4864107, -1.162289, -1.596404, -0.765414, 
    -0.02882588,
  -0.4373872, -0.1401216, 0.005158305, -0.1576672, -0.4356945, -0.5560559, 
    -0.3067232, -0.2618665, -0.5698255, -0.6518402, -0.5059419, -0.328419, 
    -0.3300303, -0.4662445, -0.578891, -0.5470877, -0.2603363, 0.06456542, 
    0.1485667, -0.0352391, -0.2826184, -0.2471529, -0.05745554, 0.1479805, 
    0.1484038, -0.04078889, -0.06603295, -0.1305023, -0.300294, -0.4196137, 
    -0.4073252, -0.3959808, -0.3991873, -0.2876966, -0.07933068, 0.04208851, 
    0.1223295, 0.1543932, 0.2277331, 0.1604159, -0.02755618, -0.1580248, 
    -0.1213713, -0.1361666, -0.1214368, -0.1412776, -0.3421075, -0.5316908, 
    -0.6160984, -0.658448, -0.6124356, -0.3904469, -0.1599617, -0.01943421, 
    0.1251781, 0.2241201, 0.3685863, 0.438508, 0.479654, 0.5403147, 
    0.2283516, -0.3249192, -0.4191253, -0.3878268, -0.1900401, -0.04266065, 
    0.0767892, 0.0001943111, -0.05083109, 0.0544586, 0.05885315, 0.07885635, 
    0.1460274, 0.05393779, 0.1161122, 0.2081532, 0.3086578, 0.3177399, 
    0.338036, 0.4006171, 0.221874, 0.1590812, 0.06109953, -0.1092129, 
    -0.2793622, -0.2095547, -0.1205077, -0.03334999, 0.03998947, -0.1400399, 
    -0.3282728, -0.3461762, -0.5597178, -0.8998222, -0.8468598, -0.6743011,
  -0.3220228, -0.3646171, -0.1991709, 0.04392802, 0.09190978, -0.04319763, 
    -0.1336762, -0.1408539, -0.2022636, -0.2812186, -0.2108085, -0.1874522, 
    -0.2175954, -0.2501313, -0.1942557, -0.1861663, -0.153647, 0.05737203, 
    0.2467437, 0.2702951, 0.09825745, -0.1870942, -0.286964, -0.171111, 
    -0.07316184, -0.05193786, -0.09280701, 0.01718652, 0.01992059, 
    -0.1514823, -0.4410493, -0.5617036, -0.5754731, -0.4582204, -0.2535821, 
    -0.0503267, 0.004295588, 0.226838, 0.4555, 0.7810538, 0.472981, 
    -0.01189899, -0.1754732, -0.106056, -0.05892062, -0.1048354, -0.263299, 
    -0.5028825, -0.6972669, -0.7851088, -0.7680182, -0.6762214, -0.4352386, 
    -0.09122801, 0.2405753, 0.4593418, 0.5839672, 0.4438632, 0.3450997, 
    0.393521, 0.2491201, -0.04355571, -0.2003754, -0.1787608, -0.1880381, 
    -0.1663422, -0.1569021, -0.2500661, -0.3095388, -0.2033213, -0.1039398, 
    -0.05146587, -0.01655364, 0.05240774, 0.1421864, 0.2580069, 0.3138498, 
    0.3340809, 0.3761871, 0.3806956, 0.3456207, 0.2980131, 0.2268221, 
    0.2212722, 0.192512, 0.1287594, 0.06638956, 0.1146965, 0.2624831, 
    0.2231762, 0.01635671, -0.1512057, -0.159718, -0.08248818, -0.007797301, 
    -0.07827252,
  0.4485178, 0.2028635, 0.02016491, -0.01951611, 0.02571505, 0.08004455, 
    0.08022361, -0.03110453, -0.1104177, -0.09352309, -0.01980895, 
    -0.09532979, -0.1787608, -0.1579113, -0.04752719, -0.07107849, 
    -0.08247173, 0.0369944, 0.2775706, 0.4350088, 0.4932119, 0.4397287, 
    0.3507639, 0.2771471, 0.2927558, 0.1841785, 0.02568269, 0.08004445, 
    0.2454254, 0.1292796, -0.1939301, -0.3706065, -0.4336599, -0.3341808, 
    -0.1126963, 0.1473134, 0.2725901, 0.4450673, 0.6083648, 0.8391753, 
    0.7001127, 0.2897449, 0.05911326, -0.1190443, -0.01269633, 0.07900292, 
    0.04282111, -0.1757988, -0.4449557, -0.575555, -0.6223807, -0.6478205, 
    -0.5540047, -0.2879076, 0.05060148, 0.3443351, 0.5330396, 0.5122547, 
    0.3129058, 0.1553372, -0.01062953, -0.09513474, -0.09923637, 
    -0.009880543, 0.06622618, 0.1055491, 0.07068583, -0.08587343, -0.2248057, 
    -0.2032399, -0.06780702, 0.01992086, 0.0103831, -0.03603618, 0.01228739, 
    0.1250641, 0.2524241, 0.3706208, 0.4529937, 0.5652496, 0.5764475, 
    0.3678864, 0.2555816, 0.1866521, 0.3513827, 0.5562491, 0.6404452, 
    0.5495272, 0.4472485, 0.3776686, 0.3078117, 0.1925285, 0.1510406, 
    0.2409493, 0.4167469, 0.5408679,
  0.5557607, 0.4980458, 0.3075673, 0.1720366, 0.03061414, 0.001968384, 
    0.06352437, 0.06564024, -0.02114359, -0.0597992, -0.02806091, 0.01290589, 
    0.08245341, 0.1595693, 0.2344879, 0.1979319, 0.140982, 0.1621084, 
    0.2492991, 0.3892893, 0.5202301, 0.6083485, 0.6319814, 0.6655588, 
    0.6680163, 0.5131987, 0.2738758, 0.1433257, 0.1518219, 0.0994456, 
    -0.1181325, -0.3159516, -0.4660168, -0.4532075, -0.2210786, 0.08058167, 
    0.286441, 0.3846833, 0.4393219, 0.5851389, 0.5956208, 0.4453765, 
    0.3332672, 0.1078278, -0.06297302, 0.04523009, 0.1568837, 0.1356272, 
    -0.04801533, -0.2329274, -0.3393404, -0.3499365, -0.2487645, -0.09459782, 
    -0.05680418, 0.1576807, 0.3609364, 0.4705396, 0.4069979, 0.1394522, 
    -0.04415846, -0.137583, -0.1013359, -0.04617631, 0.008299589, 0.0585112, 
    0.1038889, 0.06129456, -0.03084411, -0.01149191, 0.0671702, 0.05253805, 
    -0.06461692, -0.1708996, -0.2037445, -0.01906026, 0.0657379, 0.1066722, 
    0.2131173, 0.3965157, 0.5252429, 0.4576163, 0.2864573, 0.2471344, 
    0.4257312, 0.8137847, 1.159715, 1.256038, 1.071321, 0.7914219, 0.4991038, 
    0.2871408, 0.2407701, 0.3116198, 0.4363106, 0.5773911,
  0.58885, 0.5998361, 0.4535307, 0.116975, -0.1820648, -0.3151052, 
    -0.1476084, -0.08250427, -0.1761241, -0.2734385, -0.283611, -0.1767263, 
    -0.03986105, 0.04643453, 0.09586487, 0.1311351, 0.1153147, 0.09646708, 
    0.1770007, 0.3192698, 0.4310373, 0.4587067, 0.3936839, 0.3740387, 
    0.4000477, 0.4952951, 0.552717, 0.5531565, 0.5374989, 0.4182444, 
    0.2382477, 0.06254774, -0.06526792, -0.1083019, -0.06805116, 0.01817932, 
    0.07394105, 0.1213369, 0.2130849, 0.4202952, 0.6054677, 0.6556305, 
    0.5542958, 0.3132314, 0.08369046, 0.02994674, 0.1136869, 0.1231922, 
    0.07774955, -0.02321076, -0.1141612, -0.1647635, -0.1414237, -0.126564, 
    -0.03099108, 0.07675648, 0.1185211, 0.1656889, 0.1558093, 0.115168, 
    0.1217275, 0.2144194, 0.2280586, 0.174885, 0.1188304, 0.09187724, 
    0.07823792, 0.01850484, -0.05861104, -0.08688253, -0.06700948, 
    -0.1345714, -0.2622407, -0.3265309, -0.3267102, -0.2648122, -0.3049654, 
    -0.2481293, -0.077003, 0.1946277, 0.3950834, 0.4081208, 0.3472483, 
    0.2590322, 0.1607412, 0.4017079, 0.7728828, 1.216877, 1.42259, 1.300666, 
    0.956184, 0.5667793, 0.3525703, 0.3390777, 0.4394846, 0.5217112,
  0.7925282, 0.7871572, 0.5825347, 0.3382965, 0.01500549, -0.1582855, 
    -0.1925304, -0.1575043, -0.2021821, -0.2920259, -0.3637544, -0.3625337, 
    -0.3299001, -0.2980804, -0.1928885, -0.02418739, 0.06578678, 0.09272349, 
    0.1478339, 0.2991526, 0.5004544, 0.6518544, 0.648697, 0.535611, 
    0.4384104, 0.4463043, 0.5319651, 0.6595694, 0.7309397, 0.6844066, 
    0.4462227, 0.2076809, 0.04872918, 0.01082265, 0.01536357, 0.04256082, 
    0.01158753, 0.01827699, -0.01565856, 0.0143219, 0.09749247, 0.1284007, 
    0.09957594, 0.02195536, -0.06401469, -0.1211436, -0.06484479, 0.03886592, 
    0.09436727, 0.1766915, 0.1780261, -0.08917749, -0.0403657, -0.07791471, 
    -0.02467573, 0.09978724, 0.2041981, 0.1881662, 0.2410635, 0.223827, 
    0.2079579, 0.205663, 0.1869293, 0.1209951, 0.03393453, -0.02478939, 
    -0.08932406, -0.1563486, -0.1997733, -0.1665213, -0.1287283, -0.1688976, 
    -0.3213878, -0.5101736, -0.5637543, -0.5053397, -0.4015636, -0.5051118, 
    -0.3185395, -0.1104504, 0.1204905, 0.1988271, 0.222769, 0.08056533, 
    -0.07931417, -0.1760917, -0.04464674, 0.3018384, 0.6213207, 0.8493474, 
    0.8514963, 0.8302073, 0.5566396, 0.5424469, 0.607551, 0.6936675,
  0.7301422, 0.6672353, 0.5452138, 0.3454742, 0.126122, 0.03264871, 
    -0.1439626, -0.2645192, -0.3228689, -0.3632823, -0.3814465, -0.3000988, 
    -0.2760265, -0.2498547, -0.2909354, -0.1273776, -0.002849579, 0.06101763, 
    0.08884966, 0.2132312, 0.4780749, 0.7424141, 0.8963529, 0.8746408, 
    0.6828765, 0.5391265, 0.5181955, 0.589273, 0.6906891, 0.7409008, 
    0.6357084, 0.4295886, 0.2573067, 0.1099924, 0.05180562, 0.08253479, 
    0.1127431, 0.05642802, -0.01858824, -0.09087008, -0.1491222, -0.168507, 
    -0.1603689, -0.1113292, -0.106544, -0.1600108, -0.180779, -0.1349132, 
    -0.03027451, -0.217856, -0.07918429, -0.0500499, -0.1079437, 0.09135641, 
    0.06780481, 0.09584853, 0.1558909, 0.1963043, 0.1934072, 0.1854807, 
    0.1692209, 0.1277333, 0.0552724, -0.05473736, -0.1658539, -0.2467622, 
    -0.2852387, -0.2846854, -0.2174003, -0.1092297, -0.1450207, -0.2413099, 
    -0.3998872, -0.3993011, -0.6978037, -0.4900076, -0.5803071, -0.4282236, 
    -0.274171, -0.008204147, 0.03989142, 0.1292468, 0.3342432, 0.3147123, 
    0.4265125, 0.3387848, 0.2133288, 0.1068027, 0.03577399, 0.1532218, 
    0.4112785, 0.5850081, 0.6862454, 0.71551, 0.7343088, 0.7489736,
  0.6461741, 0.5012197, 0.3408518, 0.1770823, 0.002017211, -0.1201019, 
    -0.2006683, -0.2533377, -0.2851899, -0.3189139, -0.3539398, -0.3998545, 
    -0.4105643, -0.3749036, -0.2891451, -0.3209811, -0.2528985, -0.2833184, 
    -0.2958997, -0.184653, 0.006802082, 0.2788236, 0.5602038, 0.7410472, 
    0.8055655, 0.775764, 0.6908519, 0.6080556, 0.5329092, 0.5098296, 
    0.4836416, 0.4433258, 0.3723622, 0.3315257, 0.3658844, 0.3209951, 
    0.4330068, 0.4786774, 0.5359365, 0.4147938, 0.2306792, 0.09776914, 
    0.002456665, -0.02928162, -0.01787212, -0.02021586, -0.002979532, 
    0.006737264, 0.02630107, 0.04601133, 0.0726715, 0.1125315, 0.1605621, 
    0.1800608, 0.1541494, 0.1106272, 0.08017477, 0.02703351, -0.02265728, 
    -0.05457467, -0.05232859, -0.04646927, -0.05385858, -0.05986434, 
    -0.09121209, -0.1571137, -0.1993501, -0.2113618, -0.2288749, -0.2084158, 
    -0.3177258, -0.3738292, -0.3397309, -0.3977388, -0.35394, -0.316326, 
    -0.3013847, -0.2772961, -0.2327973, -0.1813324, -0.108725, -0.04560673, 
    0.1230619, 0.3201159, 0.4618965, 0.4711904, 0.4046051, 0.3752917, 
    0.315282, 0.3207181, 0.5747061, 0.5435696, 0.7777816, 0.8509589, 
    0.8229645, 0.7478668,
  0.5924306, 0.4259756, 0.2794423, 0.1240712, -0.03317158, -0.1367686, 
    -0.2171723, -0.2804536, -0.3231456, -0.3435233, -0.3804211, -0.4304537, 
    -0.4282887, -0.4624359, -0.4920908, -0.4736013, -0.4723644, -0.4153496, 
    -0.3015639, -0.1906263, -0.03966594, 0.1273099, 0.3069974, 0.4286445, 
    0.5375479, 0.7682933, 0.7443837, 0.7006826, 0.6260407, 0.5450023, 
    0.5420401, 0.4510733, 0.4068348, 0.3823232, 0.4476064, 0.489094, 
    0.518277, 0.5235993, 0.506135, 0.4333649, 0.3018707, 0.1722158, 
    0.05027568, -0.03004659, -0.05890401, -0.03431091, 0.03670146, 0.14204, 
    0.2402984, 0.3298492, 0.3530751, 0.363736, 0.3493642, 0.3386383, 
    0.3221344, 0.2869293, 0.2505035, 0.2162587, 0.1721181, 0.112678, 
    0.04667866, 0.002782106, -0.03909618, -0.07415473, -0.1249523, -0.131007, 
    -0.1579764, -0.1565117, -0.1550957, -0.1418958, -0.1387707, -0.1031424, 
    -0.09964305, -0.04451597, -0.05537206, -0.03514099, -0.06816506, 
    -0.07073669, -0.133546, -0.1137054, -0.05338669, -0.007732391, 
    0.04576707, 0.101724, 0.126838, 0.159553, 0.2058909, 0.2530751, 
    0.3124011, 0.4051741, 0.4967922, 0.7588204, 0.5446274, 0.6180488, 
    0.7361155, 0.7243153,
  0.38815, 0.4179189, 0.3277171, 0.2450836, 0.1011546, 0.04846904, 
    -0.004183959, 0.04469299, -0.03046978, -0.08987734, -0.1515147, 
    -0.1628917, -0.2049163, -0.1854666, -0.1408865, -0.1111827, -0.03857523, 
    0.01962775, 0.05856019, 0.1116201, 0.166926, 0.2279124, 0.2934884, 
    0.3298817, 0.3579416, 0.322525, 0.3266266, 0.3488759, 0.3730296, 
    0.3833323, 0.3963043, 0.3705556, 0.3508453, 0.3534495, 0.3536611, 
    0.3542958, 0.3221995, 0.285318, 0.2502106, 0.2033356, 0.1496409, 
    0.0936025, 0.04090068, -0.004476931, -0.03354594, -0.04176534, 
    -0.03079529, -0.006137085, 0.02005107, 0.03940328, 0.06274313, 
    0.09220275, 0.1218252, 0.1624339, 0.1909007, 0.2108388, 0.2163401, 
    0.2071604, 0.1698883, 0.1260569, 0.073062, 0.02029508, -0.03296018, 
    -0.06082475, -0.08382279, -0.1198579, -0.1266124, -0.1156098, -0.1314628, 
    -0.1100109, -0.07760531, -0.2247407, -0.1601247, -0.1142751, -0.09477633, 
    -0.07775164, -0.06645632, -0.06227338, -0.08077931, -0.08110476, 
    -0.08121872, -0.0829277, -0.06611454, -0.05752075, -0.02166456, 
    0.03310445, 0.09457907, 0.1565092, 0.2255523, 0.2976875, 0.3772286, 
    0.4427395, 0.5000315, 0.505126, 0.4753571, 0.4313141,
  0.2281402, 0.2221506, 0.2063791, 0.1987294, 0.1740387, 0.1569814, 
    0.1505849, 0.1510406, 0.1470856, 0.1285309, 0.1123851, 0.1033844, 
    0.09168193, 0.09506734, 0.1117503, 0.1400218, 0.1535634, 0.1731109, 
    0.2052561, 0.2416657, 0.2679515, 0.2887034, 0.3054515, 0.3112783, 
    0.304719, 0.2813629, 0.2594065, 0.2418447, 0.23343, 0.2219228, 0.2131012, 
    0.1871735, 0.1536774, 0.1233714, 0.1032542, 0.08328348, 0.06458232, 
    0.04509989, 0.01887919, -0.01575623, -0.05559997, -0.09067485, 
    -0.1262054, -0.1511241, -0.1721527, -0.1817881, -0.1823415, -0.1769867, 
    -0.1739268, -0.1742523, -0.1706879, -0.167628, -0.1538422, -0.1266449, 
    -0.1061859, -0.09202576, -0.08515728, -0.09246522, -0.09290463, 
    -0.1004243, -0.09795028, -0.1032237, -0.1259289, -0.1546561, -0.1823579, 
    -0.2055025, -0.2175792, -0.2236176, -0.2443533, -0.2810883, -0.3118989, 
    -0.3548187, -0.3628754, -0.3850759, -0.3745615, -0.4446789, -0.4814954, 
    -0.4795098, -0.4238132, -0.4349948, -0.3789401, -0.334946, -0.2780936, 
    -0.2305675, -0.1828299, -0.1364593, -0.09638774, -0.05022888, 
    0.001707964, 0.08126526, 0.1472646, 0.1744293, 0.2118968, 0.2194814, 
    0.2225901, 0.2270335,
  -0.0306651, -0.006836951, 0.02063698, 0.03981018, 0.05226135, 0.06485897, 
    0.07332253, 0.07477111, 0.07451069, 0.08006084, 0.08147684, 0.09104717, 
    0.1037913, 0.107665, 0.1191722, 0.1213531, 0.1282216, 0.1362457, 
    0.1404287, 0.1418447, 0.1503408, 0.1553375, 0.1552073, 0.1619944, 
    0.1647776, 0.1664215, 0.1741526, 0.1768707, 0.1746409, 0.1689768, 
    0.160497, 0.1464671, 0.1346669, 0.1198395, 0.103775, 0.08803609, 
    0.06979065, 0.04946186, 0.02529195, 0.004279584, -0.02078553, 
    -0.04056092, -0.0605479, -0.07882589, -0.09741312, -0.1136078, 
    -0.1269867, -0.1416351, -0.1498058, -0.1555187, -0.1684581, -0.172462, 
    -0.1778005, -0.1792165, -0.1731618, -0.1645029, -0.1580088, -0.146225, 
    -0.1482759, -0.1436046, -0.1386241, -0.1325532, -0.1386079, -0.1374522, 
    -0.1480643, -0.1641124, -0.1761892, -0.1903006, -0.2024261, -0.2209157, 
    -0.2392263, -0.2591156, -0.2797862, -0.3049001, -0.3288422, -0.3462738, 
    -0.3588063, -0.3635915, -0.3649262, -0.358432, -0.3471853, -0.3371267, 
    -0.3251964, -0.3062673, -0.2845225, -0.2634288, -0.2385427, -0.21268, 
    -0.1922536, -0.1655284, -0.1386729, -0.1167979, -0.09451601, -0.0870941, 
    -0.0748708, -0.04921979,
  -0.1220279, -0.1429915, -0.1629786, -0.1816959, -0.1982164, -0.2127347, 
    -0.2253971, -0.2360096, -0.2446842, -0.2518787, -0.2576566, -0.2609925, 
    -0.2614164, -0.2583723, -0.2520738, -0.2430887, -0.2318096, -0.2188375, 
    -0.2034895, -0.1867256, -0.16739, -0.1467842, -0.125479, -0.1039132, 
    -0.08140343, -0.05806351, -0.03332353, -0.007591248, 0.0191021, 
    0.04621792, 0.0740819, 0.1022553, 0.1308203, 0.1595802, 0.1864524, 
    0.2137141, 0.2412534, 0.2689543, 0.2960691, 0.322648, 0.3481035, 
    0.3713303, 0.3925858, 0.4112377, 0.4272203, 0.4398022, 0.4540291, 
    0.4449463, 0.4420815, 0.4365311, 0.4261637, 0.3986082, 0.3803482, 
    0.397161, 0.3381772, 0.3555436, 0.3538508, 0.3414645, 0.2702737, 
    0.1851168, 0.2055759, 0.2449479, 0.2137465, 0.2014422, 0.1882906, 
    0.1768003, 0.1714938, 0.1720474, 0.1790459, 0.1722426, 0.1762791, 
    0.1841407, 0.1930437, 0.1928976, 0.1917086, 0.2011328, 0.1967545, 
    0.2161231, 0.2211685, 0.2155538, 0.2122009, 0.2050068, 0.1960706, 
    0.1820894, 0.1647554, 0.1454845, 0.1238862, 0.1000419, 0.0747329, 
    0.04898405, 0.02263379, -0.003359079, -0.0283916, -0.05344057, 
    -0.07739925, -0.1003485,
  -0.2659898, -0.3182354, -0.3600168, -0.391901, -0.4142323, -0.4239645, 
    -0.4219956, -0.4125066, -0.398737, -0.3848209, -0.3717508, -0.3567281, 
    -0.335911, -0.3068259, -0.2710025, -0.2305408, -0.187816, -0.1457748, 
    -0.1052312, -0.06491578, -0.02136111, 0.02544874, 0.07699496, 0.1271577, 
    0.1672622, 0.1918226, 0.2037532, 0.2070739, 0.2028749, 0.192718, 
    0.1764264, 0.1547461, 0.1316667, 0.1081152, 0.08680916, 0.07108593, 
    0.06322289, 0.06224728, 0.067276, 0.08011723, 0.1017323, 0.1397047, 
    0.1304932, 0.1837482, 0.2125583, 0.201117, 0.247992, 0.2534928, 
    0.2374606, 0.2164483, 0.1471777, 0.1846776, 0.1699321, 0.1605897, 
    0.1052506, 0.1232197, 0.09006453, 0.05966091, 0.0428803, 0.02627882, 
    0.02868772, 0.03090131, 0.0390234, 0.04052067, 0.04325509, 0.03397775, 
    0.01329064, -0.01138389, -0.03680724, -0.05174854, -0.05482477, 
    -0.04815137, -0.04855847, -0.0370667, -0.06016278, -0.04808617, 
    -0.03037691, -0.01929379, -0.02113295, 0.009189606, 0.02597046, 
    0.01246095, 0.082057, 0.103004, 0.1827241, 0.2288341, 0.2581149, 
    0.270843, 0.2653911, 0.2363868, 0.1851501, 0.1167254, 0.03890944, 
    -0.04759741, -0.1306705, -0.203197,
  -0.1162014, -0.1876693, -0.230963, -0.2606182, -0.2846088, -0.301488, 
    -0.3154855, -0.3276274, -0.3419666, -0.3591052, -0.3714421, -0.3808987, 
    -0.3676331, -0.3252666, -0.2531314, -0.1568265, -0.0458889, 0.07268286, 
    0.1875422, 0.2894791, 0.3685803, 0.4194429, 0.4289643, 0.4094006, 
    0.3824149, 0.3635997, 0.357285, 0.3493748, 0.3242128, 0.2832947, 
    0.2308209, 0.1782815, 0.1315041, 0.09104156, 0.0501399, 0.01057291, 
    -0.01805687, -0.04660511, -0.07678032, -0.1003642, -0.1331277, 
    -0.1040597, -0.05376625, -0.03639936, 0.03064132, 0.03078771, 0.06366491, 
    0.1113375, 0.1551691, 0.1863215, 0.1898695, 0.1583265, 0.1008561, 
    0.03335881, -0.02502334, -0.05171597, -0.06922919, -0.07733428, 
    -0.05558896, -0.02699184, 0.004078388, 0.008684635, -0.02534819, 
    -0.0722394, -0.1015692, -0.1138244, -0.1106837, -0.109089, -0.1088937, 
    -0.1073308, -0.1098535, -0.1051493, -0.1171937, -0.1596746, -0.1672268, 
    -0.1658268, -0.1373277, -0.1488023, -0.09533453, -0.04312181, 
    -0.00479126, 0.02292585, 0.07483029, 0.1349377, 0.2062593, 0.272405, 
    0.3391856, 0.3978121, 0.4186454, 0.453656, 0.3914814, 0.3199801, 
    0.2171321, 0.1270118, 0.04136705, -0.03693628,
  0.06716424, 0.0256115, -0.03042692, -0.09873754, -0.1704662, -0.2534084, 
    -0.3435774, -0.4389873, -0.5089746, -0.4945054, -0.3888574, -0.225316, 
    -0.05677748, 0.0662365, 0.1429296, 0.2298927, 0.3008237, 0.3573833, 
    0.3539158, 0.3159761, 0.352337, 0.4615009, 0.5237074, 0.5212667, 
    0.4459893, 0.3612723, 0.329062, 0.3158624, 0.2981708, 0.2656512, 
    0.2369401, 0.200156, 0.1427341, 0.07141244, 0.01875925, 0.001018524, 
    0.01006842, 0.01672578, 0.02015996, 0.02416372, 0.02279663, 
    -0.0006251335, 0.02849293, 0.05567408, 0.06192398, 0.09569716, 
    0.06150103, 0.08526397, 0.1256285, 0.1393168, 0.1343522, 0.07357717, 
    -0.04292679, -0.1587145, -0.2245349, -0.2591216, -0.3167225, -0.2673736, 
    -0.2159408, -0.2252839, -0.182429, -0.1709217, -0.1447987, -0.139395, 
    -0.1971097, -0.2421618, -0.2807517, -0.3140686, -0.3040752, -0.2893295, 
    -0.2703028, -0.2558007, -0.2404037, -0.2019601, -0.1608629, -0.1051004, 
    -0.08960557, -0.04873657, -0.01584363, -0.00562191, -0.04336643, 
    0.02985942, 0.08275676, 0.1239026, 0.1840262, 0.2639904, 0.3321381, 
    0.3662202, 0.4033134, 0.4759699, 0.4469335, 0.3962171, 0.4143488, 
    0.3167574, 0.207952, 0.1268649,
  0.02273107, -0.08633471, -0.1707911, -0.3084049, -0.4431705, -0.4934635, 
    -0.5096421, -0.5368242, -0.5466881, -0.4979906, -0.3298078, -0.1608953, 
    -0.003896236, 0.09276724, 0.1403418, 0.07509136, -0.09157562, -0.1811914, 
    -0.1618395, -0.1177638, -0.03264046, 0.1201432, 0.3279886, 0.5024996, 
    0.623284, 0.7214947, 0.6837339, 0.548317, 0.4217377, 0.3372169, 
    0.2661557, 0.2123637, 0.1543722, 0.06786489, -0.02285814, -0.1069889, 
    -0.1690173, -0.1860094, -0.1722722, -0.1555076, -0.1428123, -0.1515689, 
    -0.2279525, -0.2665267, -0.3201561, -0.2753482, -0.2683492, -0.09937143, 
    0.03588223, 0.09878874, 0.08669591, -0.0148344, -0.1774809, -0.3213448, 
    -0.4097075, -0.4776437, -0.5289459, -0.5420643, -0.513858, -0.4248769, 
    -0.3672596, -0.3549548, -0.3842679, -0.4216868, -0.4609935, -0.456029, 
    -0.4057686, -0.3444568, -0.3002021, -0.2720119, -0.197598, -0.1654854, 
    -0.1743072, -0.2209543, -0.2093493, -0.2397693, -0.220466, -0.2063058, 
    -0.2419015, -0.2869373, -0.2567942, -0.2542223, -0.1607329, -0.02676487, 
    0.1183687, 0.2531994, 0.3757743, 0.4354258, 0.4375256, 0.4173595, 
    0.452711, 0.3578707, 0.2594331, 0.2134206, 0.152809, 0.08868194,
  0.1028414, 0.0476979, 0.02452099, -0.0349189, 0.004908562, -0.05609322, 
    -0.03805947, 0.09800816, 0.0152936, -0.04041958, -0.05529642, -0.1239166, 
    -0.1251533, -0.08124053, -0.03076839, 0.008472919, -0.1494379, 
    -0.1918526, -0.1148992, -0.0798893, 0.04411769, 0.07234013, 0.132692, 
    0.1969986, 0.248805, 0.2011647, 0.06810856, -0.08391047, -0.166266, 
    -0.1959538, -0.1769924, -0.1726627, -0.1854072, -0.2747946, -0.3057032, 
    -0.3082252, -0.2470112, -0.2004457, -0.09885073, -0.1075263, -0.1295476, 
    -0.1629949, -0.2225652, -0.2473207, -0.1829975, -0.1307514, -0.01664019, 
    0.0814712, 0.06840134, -0.04308963, -0.2429106, -0.4423572, -0.6076242, 
    -0.6642973, -0.6543527, -0.6490467, -0.6649972, -0.7326894, -0.7936757, 
    -0.8174711, -0.8205799, -0.8252186, -0.8073963, -0.7735096, -0.6924061, 
    -0.5422596, -0.3404692, -0.1304757, 0.04185499, 0.1455008, 0.2115164, 
    0.1890067, 0.1320568, 0.02575797, -0.07678115, -0.1986884, -0.3024647, 
    -0.3217355, -0.4188871, -0.4472075, -0.3686268, -0.236449, -0.01167691, 
    0.2407319, 0.4205496, 0.4884532, 0.510377, 0.512379, 0.4758882, 0.426116, 
    0.3587658, 0.302646, 0.235019, 0.186956, 0.1369884, 0.1137789,
  -0.2443592, -0.2764882, -0.3029041, -0.2419664, -0.1416247, -0.07899451, 
    -0.05018568, -0.06066751, -0.1010973, -0.1209376, -0.1046132, 
    -0.08708382, -0.04940478, -0.01486695, -0.02735031, -0.06528974, 
    -0.1420796, -0.2100973, -0.233144, -0.2529199, -0.2643461, -0.2323312, 
    -0.1503323, -0.03094757, -0.01815462, -0.016397, -0.1061428, -0.2223048, 
    -0.328213, -0.3808987, -0.391771, -0.379743, -0.3103098, -0.286123, 
    -0.3650615, -0.2912498, -0.3091369, -0.3448961, -0.4096583, -0.4515207, 
    -0.4240956, -0.3733958, -0.3326732, -0.2809801, -0.226602, -0.2411854, 
    -0.3571847, -0.5878486, -0.8858793, -1.157152, -1.314688, -1.359463, 
    -1.335114, -1.262474, -1.113809, -1.026618, -1.006257, -1.022354, 
    -1.02766, -0.9705148, -0.8795317, -0.8076567, -0.7133533, -0.5946034, 
    -0.4107004, -0.1915597, 0.002499517, 0.1251883, 0.2744884, 0.3367769, 
    0.3440685, 0.256308, 0.2449148, 0.191562, 0.06542265, -0.03589565, 
    -0.0451405, -0.06784552, -0.08085012, -0.04190159, -0.04719132, 
    0.06123966, 0.200286, 0.3065034, 0.3477794, 0.3395112, 0.3564057, 
    0.3605399, 0.321103, 0.2406831, 0.1109956, -0.005199045, -0.1044341, 
    -0.1499907, -0.1716541, -0.2072173,
  -0.5408762, -0.4825103, -0.3727283, -0.2188058, -0.08311245, -0.02349332, 
    -0.04160857, -0.1066639, -0.1415109, -0.1830799, -0.2426502, -0.2768136, 
    -0.3284413, -0.359561, -0.4562082, -0.5802479, -0.6400948, -0.6672271, 
    -0.6475818, -0.6070707, -0.6131418, -0.6001698, -0.5653228, -0.5472889, 
    -0.6025949, -0.6754953, -0.7503812, -0.8519602, -0.9805735, -1.05458, 
    -1.013972, -0.8740793, -0.7160715, -0.776423, -0.9829333, -1.079613, 
    -1.011889, -1.074632, -1.192422, -1.318529, -1.332689, -1.251374, 
    -1.221605, -1.388824, -1.524469, -1.744602, -1.960765, -2.159804, 
    -2.270367, -2.034804, -1.712279, -1.462637, -1.183942, -1.096426, 
    -0.9197003, -0.8983949, -0.9216539, -0.9255275, -0.9293689, -0.9085032, 
    -1.00974, -0.9669504, -0.8345935, -0.6116932, -0.4722075, -0.3694569, 
    -0.3683989, -0.1974191, 0.01553661, 0.06584597, 0.156487, 0.07043588, 
    -0.1387436, -0.3779364, -0.5217678, -0.6482326, -0.6717841, -0.6379299, 
    -0.6422106, -0.5421293, -0.552497, -0.4731839, -0.296084, -0.2176499, 
    -0.184642, -0.1406153, -0.1119369, -0.109789, -0.1421946, -0.2234932, 
    -0.3204335, -0.3775624, -0.4080799, -0.4189848, -0.4560779, -0.5193104,
  -0.4772529, -0.352904, -0.2172432, -0.08345419, -0.1159412, -0.1181222, 
    -0.2779039, -0.3968005, -0.5384995, -0.7009994, -0.8481512, -1.033291, 
    -1.130817, -1.233503, -1.315355, -1.478604, -1.544424, -1.40821, 
    -1.228473, -1.069115, -0.9163318, -0.9050688, -1.017113, -1.268236, 
    -1.502807, -1.632185, -1.561563, -1.556127, -1.499844, -1.643757, 
    -1.533747, -1.262784, -1.123981, -1.12761, -1.279222, -1.391055, 
    -1.428701, -1.422386, -1.496947, -1.656549, -1.839346, -1.995954, 
    -2.067129, -2.09514, -2.089443, -2.167992, -2.210325, -2.166282, 
    -1.955052, -1.660977, -1.410896, -1.28002, -1.270775, -1.286448, 
    -1.270319, -1.251455, -1.221263, -1.170092, -1.077741, -1.042503, 
    -1.083047, -1.11083, -0.9987211, -0.8305897, -0.7324777, -0.6426828, 
    -0.486742, -0.27294, -0.09217811, -0.01935911, -0.05611038, -0.1558988, 
    -0.3459215, -0.6159248, -0.8853742, -1.029059, -1.040354, -1.017731, 
    -0.9935122, -0.9107318, -0.7617581, -0.6246324, -0.5887432, -0.6635478, 
    -0.6018946, -0.5466865, -0.5065657, -0.4554266, -0.3923246, -0.3185779, 
    -0.3264232, -0.3587796, -0.421459, -0.4857654, -0.5590726, -0.55349,
  -0.7786691, -0.7575263, -0.7312731, -0.6179757, -0.5955956, -0.6508198, 
    -0.800853, -0.8659732, -0.900202, -0.9854558, -1.104108, -1.186302, 
    -1.247728, -1.3482, -1.481582, -1.593431, -1.631143, -1.623932, 
    -1.641364, -1.754629, -1.980556, -2.099193, -2.154043, -2.151374, 
    -2.164411, -2.080117, -1.885977, -1.739183, -1.703864, -1.591104, 
    -1.305931, -1.041331, -0.9612365, -1.009414, -1.155052, -1.383096, 
    -1.586563, -1.660684, -1.721833, -1.825755, -1.906484, -1.976553, 
    -2.002953, -1.928555, -1.821654, -1.742503, -1.657379, -1.611302, 
    -1.568089, -1.466429, -1.273363, -1.079255, -0.9933167, -0.9349673, 
    -0.8393781, -0.778522, -0.7331771, -0.6177316, -0.4996161, -0.4787181, 
    -0.5923898, -0.7108303, -0.7312733, -0.6945382, -0.5772043, -0.3717518, 
    -0.1388251, -0.003441095, -0.003864288, -0.01058638, -0.04352915, 
    -0.2058496, -0.5095763, -0.8036194, -0.9476628, -0.9652247, -0.9325094, 
    -0.898623, -0.7867255, -0.6973212, -0.6622784, -0.5704975, -0.60235, 
    -0.7075427, -0.8067608, -0.8811748, -0.8954487, -0.8333077, -0.7373765, 
    -0.6199615, -0.6895742, -0.7425361, -0.7664782, -0.7942289, -0.9129466, 
    -0.8746979,
  -0.7709213, -0.6857815, -0.6765363, -0.6120176, -0.5393453, -0.5534897, 
    -0.6082909, -0.6102278, -0.6431706, -0.7154851, -0.7601953, -0.807982, 
    -0.8918033, -1.014281, -1.117308, -1.176146, -1.221133, -1.306143, 
    -1.418577, -1.493675, -1.498736, -1.473639, -1.500332, -1.551243, 
    -1.552122, -1.546035, -1.507363, -1.363678, -1.172809, -0.9541892, 
    -0.7582417, -0.7287333, -0.8565335, -0.9591699, -1.053132, -1.272646, 
    -1.409414, -1.377448, -1.400381, -1.455459, -1.402253, -1.307786, 
    -1.345954, -1.404076, -1.279857, -1.076585, -0.9711657, -0.9514554, 
    -0.9920313, -0.9013412, -0.7422426, -0.6092184, -0.3946187, -0.1367257, 
    -0.0298897, -0.006875157, 0.06203747, 0.1153903, 0.01376283, -0.2023344, 
    -0.4009185, -0.4227446, -0.274421, -0.108438, 0.02149373, 0.2017672, 
    0.3365327, 0.2398206, 0.02600229, -0.1381742, -0.2703844, -0.4980366, 
    -0.7408264, -0.8069072, -0.7379949, -0.7934637, -0.873558, -0.7391667, 
    -0.4639547, -0.5346253, -0.644635, -0.5298405, -0.4743717, -0.6046288, 
    -0.699827, -0.6720603, -0.6268134, -0.6196847, -0.6620184, -0.7732491, 
    -0.8744373, -0.9858958, -1.081387, -1.092878, -1.063256, -0.9479235,
  -0.3626698, -0.1914773, -0.1481993, -0.180784, -0.2099187, -0.1635482, 
    -0.06346703, 0.007643223, 0.007642984, -0.05847025, -0.1700912, 
    -0.3679917, -0.6125555, -0.767715, -0.8343003, -0.9225004, -1.074046, 
    -1.190387, -1.204678, -1.185325, -1.16345, -1.158811, -1.229661, 
    -1.311839, -1.34514, -1.346019, -1.289508, -1.116575, -0.8996646, 
    -0.8043029, -0.8037658, -0.805752, -0.7796776, -0.7169824, -0.6978908, 
    -0.6891017, -0.583714, -0.5190172, -0.6339583, -0.7455144, -0.7140203, 
    -0.6452212, -0.7011461, -0.6824121, -0.453099, -0.2163153, -0.2443907, 
    -0.3393614, -0.2724023, -0.125088, -0.0739001, 0.06480432, 0.4511322, 
    0.7376071, 0.6630467, 0.4523534, 0.44262, 0.541025, 0.496575, 0.3084241, 
    0.1371675, 0.1741792, 0.3117118, 0.4263276, 0.4232027, 0.4200613, 
    0.4332124, 0.3351169, 0.1215426, -0.09935582, -0.2675197, -0.3063862, 
    -0.2235413, -0.1477926, -0.1643457, -0.2364163, -0.2677474, -0.206924, 
    -0.01040649, -0.08923149, -0.224534, -0.2142808, -0.2659729, -0.3789449, 
    -0.2963932, -0.1555569, -0.1249743, -0.1839261, -0.3686918, -0.6376694, 
    -0.8535874, -1.013646, -1.082559, -1.012523, -0.855329, -0.6335353,
  0.2243259, 0.1934021, 0.06923199, 0.02263403, 0.1390564, 0.3898051, 
    0.5214615, 0.4665949, 0.3271255, 0.0829854, -0.2685933, -0.6425352, 
    -0.8398335, -0.8667541, -0.8578186, -0.9609761, -1.132151, -1.206923, 
    -1.158323, -1.151618, -1.181647, -1.189883, -1.17984, -1.185553, 
    -1.218105, -1.159544, -1.006175, -0.8923078, -0.688271, -0.3722718, 
    -0.1031148, 0.06693721, 0.126296, 0.1012959, 0.08869791, 0.1949315, 
    0.3736098, 0.3120542, 0.1332946, 0.1016378, 0.05785537, 0.003932714, 
    -0.06434536, -0.09190059, 0.1238546, 0.3512137, 0.3325782, 0.4200944, 
    0.4613699, 0.320273, 0.2194918, 0.4830661, 0.8341563, 0.8896742, 
    0.7248627, 0.5922946, 0.6542412, 0.8330008, 0.9101819, 0.7065196, 
    0.4416596, 0.4179617, 0.5333753, 0.59428, 0.6215101, 0.7152437, 
    0.7306408, 0.5856537, 0.3377862, 0.04498029, -0.09841108, 0.0173924, 
    0.1634867, 0.1734478, 0.2328389, 0.5333436, 0.7963643, 0.6312931, 
    0.3172626, 0.1443291, 0.02624631, -0.04185271, -0.01618505, 0.1939383, 
    0.4548597, 0.4568616, 0.1684501, -0.1871003, -0.5749091, -0.9123765, 
    -1.055996, -1.044717, -0.8288642, -0.5787177, -0.3805895, -0.02541375,
  0.4170182, 0.3370864, 0.4018977, 0.5212498, 0.6153905, 0.647926, 0.4399183, 
    0.1953707, -0.03102899, -0.4297268, -0.8193259, -0.9734273, -0.8891175, 
    -0.8044331, -0.9153218, -1.180849, -1.342406, -1.230215, -1.107493, 
    -1.073297, -0.9463605, -0.7844143, -0.7098211, -0.623835, -0.5498605, 
    -0.4468006, -0.25668, 0.006096601, 0.5247818, 0.9634374, 1.019736, 
    0.902321, 0.7632258, 0.7887468, 0.9351335, 1.050629, 1.104161, 0.9454694, 
    0.8069437, 0.6540956, 0.3031185, 0.1647556, 0.3293062, 0.4450778, 
    0.5826589, 0.7965752, 0.8697032, 0.9059989, 0.8297781, 0.4667086, 
    0.3782157, 0.585361, 0.6570244, 0.6608653, 0.7102793, 0.8361911, 
    1.046705, 1.245696, 1.137282, 0.7054455, 0.4962658, 0.6973401, 0.8954519, 
    0.9215754, 0.8957287, 0.9350678, 0.9029877, 0.6506115, 0.2867609, 
    0.004127264, 0.06475592, 0.2322361, 0.3238215, 0.4493101, 0.649261, 
    1.153428, 1.473594, 0.8964937, 0.2139257, 0.09250605, 0.0792737, 
    0.0664317, 0.4010997, 0.7056897, 0.5957775, 0.1582287, -0.3364326, 
    -0.7679917, -1.072663, -1.113451, -0.928327, -0.6905015, -0.3800524, 
    -0.145287, -0.01105809, 0.2733004,
  0.730185, 0.7977961, 0.8549736, 0.85901, 0.9339122, 0.8401297, 0.6391206, 
    0.5628512, 0.2904064, -0.2711492, -0.4487529, -0.2158589, -0.1913147, 
    -0.4132059, -0.7466207, -0.9923563, -0.9684467, -0.7802145, -0.5835844, 
    -0.3653061, -0.02606475, 0.2585704, 0.3162527, 0.3155533, 0.4251233, 
    0.5858329, 0.7079684, 0.9382743, 1.332024, 1.321168, 1.16163, 1.218824, 
    1.143385, 1.107708, 1.158489, 1.083262, 0.9574642, 0.638356, 0.5311947, 
    0.4802182, 0.382399, 0.443092, 0.6161876, 0.7231375, 0.7643322, 
    0.9549409, 0.9570406, 0.7926689, 0.6427991, 0.4469007, 0.5455986, 
    0.6973076, 0.7059828, 0.917099, 1.133913, 1.26858, 1.4268, 1.395957, 
    1.104387, 0.7786225, 0.8462334, 1.021461, 0.9435153, 0.8657647, 0.754941, 
    0.7556895, 0.6045992, 0.2894953, 0.05525041, -0.0241766, 0.1811295, 
    0.2884865, 0.3655372, 0.6534277, 0.7928478, 1.238535, 1.491285, 
    0.5933362, 0.0006766021, 0.1310965, 0.3284761, 0.3666108, 0.6018649, 
    0.5146089, -0.07713926, -0.6087797, -1.010635, -1.193219, -1.126797, 
    -0.8751372, -0.5523669, -0.2662506, -0.03252637, 0.1684664, 0.3663342, 
    0.5742769,
  1.105413, 1.076018, 0.9786714, 1.079779, 1.162998, 0.756943, 0.5599702, 
    0.5404065, 0.128525, -0.356908, -0.2413478, 0.1516207, -0.0001859665, 
    -0.3289943, -0.5069566, -0.6806548, -0.4488673, -0.1945869, 0.05951452, 
    0.570273, 0.920094, 0.9851817, 1.028232, 0.946933, 0.8375908, 0.8875255, 
    0.9229262, 0.997324, 1.078526, 1.007806, 1.150758, 1.110556, 0.8140393, 
    0.7332776, 0.6494395, 0.5219657, 0.4920503, 0.3696545, 0.277646, 
    0.1314708, 0.2981702, 0.6492769, 0.5039969, 0.5310965, 0.6380464, 
    0.7338635, 0.7303804, 0.6566662, 0.7554454, 0.7514253, 0.8249604, 
    0.895859, 0.787493, 0.9813407, 1.233994, 1.378167, 1.350595, 1.120664, 
    1.00774, 0.9303805, 0.9670666, 0.7957937, 0.571575, 0.6145765, 0.5913995, 
    0.6541598, 0.4606214, 0.1144302, 0.1213964, 0.101751, 0.1715589, 
    0.2324313, 0.3948336, 0.6524832, 0.7029716, 1.104306, 1.061126, 0.35831, 
    -0.04987678, 0.1604259, 0.4980076, 0.4100353, 0.4080985, 0.1341726, 
    -0.7750554, -1.307428, -1.320758, -1.124437, -0.7023995, -0.2070705, 
    0.1586195, 0.4943126, 0.7014253, 0.8184826, 0.9603935, 1.054388,
  0.9959083, 0.9780209, 1.13917, 1.190765, 0.8050718, 0.3490002, 0.1682384, 
    -0.1002673, -0.20043, -0.2152578, 0.04546845, 0.4432059, -0.02220753, 
    -0.6759989, -0.6727933, -0.5698475, -0.289867, 0.01779896, 0.2619233, 
    0.644264, 0.8551365, 0.8139744, 0.8292902, 0.7786716, 0.5890884, 
    0.5144305, 0.4881611, 0.5138769, 0.6251886, 0.7298274, 0.7938898, 
    0.4507254, 0.2333263, 0.4470633, 0.3031506, 0.1435314, 0.2331961, 
    0.2641693, 0.2653087, 0.006584793, 0.3289318, 0.8147228, 0.5964611, 
    0.6805757, 0.6489189, 0.4812431, 0.4373468, 0.4132905, 0.618499, 
    0.5068779, 0.340911, 0.4255464, 0.4715263, 0.7377208, 0.9705821, 
    0.977353, 0.9668386, 0.9954194, 1.024244, 0.8238211, 0.6721284, 
    0.5641369, 0.447812, 0.6048595, 0.5020925, 0.3968517, 0.241741, 
    0.04771435, 0.1373302, 0.1117444, 0.2157156, 0.3606538, 0.4652112, 
    0.5076917, 0.6183696, 1.011338, 0.5507102, -0.1038969, -0.3112049, 
    0.06343703, 0.7663668, 0.4891369, 0.2189221, -0.1122792, -1.082672, 
    -1.733991, -1.124356, -0.4079658, -0.06857753, 0.3920992, 0.6167247, 
    0.6698498, 0.8064873, 0.9297618, 1.024245, 1.063681,
  0.8690691, 0.8718195, 0.9031835, 0.59166, 0.2126243, 0.121217, 0.02606723, 
    -0.1555569, -0.04100639, -0.04346402, 0.1330985, 0.6447206, 0.0551362, 
    -0.7543681, -0.5075103, -0.3101796, -0.2433988, -0.1424711, 0.1473727, 
    0.3992445, 0.6406507, 0.7360616, 0.6022563, 0.4120708, 0.1793396, 
    0.1448827, 0.1761813, 0.2941666, 0.5061951, 0.5237727, 0.2610283, 
    -0.1023831, -0.07263064, -0.01330447, -0.227562, 0.002971292, 0.295192, 
    0.3353128, 0.2427343, 0.2279227, 0.7516694, 0.9215915, 0.6085551, 
    0.5632911, 0.3301697, 0.1187277, 0.1158133, 0.00474596, -0.005019903, 
    -0.03996444, -0.0114814, 0.2334081, 0.4430598, 0.6239352, 0.713958, 
    0.6857355, 0.9158948, 1.014153, 0.8388764, 0.7370209, 0.7606701, 
    0.7539644, 0.5614513, 0.4983166, 0.3402762, 0.2133231, 0.2320405, 
    0.1628185, 0.1267996, 0.08614209, 0.1340915, 0.143369, 0.1914654, 
    0.3486753, 0.5279064, 0.5682373, 0.1540947, -0.09639382, -0.3539128, 
    0.03716737, 0.46749, 0.08453077, -0.04707736, 0.2202892, -0.3137761, 
    -0.8855532, -0.4554424, 0.2986585, 0.3712658, 0.5241303, 0.6204519, 
    0.6900324, 0.8145115, 0.9448667, 0.9600036, 0.90499,
  0.5376234, 0.4255476, 0.2255297, -0.006158352, 0.136826, -0.05741259, 
    -0.1965728, -0.1801991, -0.03218472, -0.1444894, 0.02297476, 0.3593688, 
    -0.1103098, -0.1927316, -0.1551173, -0.3071194, -0.1749084, -0.06670523, 
    0.1806581, 0.4331155, 0.6172953, 0.5833921, 0.4264581, 0.3129168, 
    0.1437273, 0.07079458, 0.08384752, 0.1378679, 0.1898699, 0.04115534, 
    -0.2609115, -0.5447979, -0.2171285, -0.1070049, -0.06392288, 0.2924414, 
    0.6348242, 0.6760681, 0.3138765, 0.4941499, 0.6701103, 0.4304788, 
    0.2500424, 0.04180646, -0.1646869, -0.2460508, -0.2648661, -0.2612691, 
    -0.2124248, -0.09859037, 0.02030587, 0.1764581, 0.3336356, 0.3789481, 
    0.555283, 0.6610122, 0.8583102, 0.7860121, 0.6573664, 0.8023528, 
    0.6452566, 0.4652924, 0.3340425, 0.1977633, 0.1676525, 0.2273368, 
    0.2293712, 0.1400809, 0.02974582, 0.03472638, 0.08860016, 0.1046326, 
    0.2546482, 0.2529879, 0.06688833, -0.05710602, -0.1631246, -0.06060272, 
    -0.1629298, -0.03015029, -0.03456092, -0.1723215, -0.08955774, 
    -0.02922213, -0.06537139, -0.2944243, 0.03008735, 0.4456148, 0.4593843, 
    0.5156509, 0.5537854, 0.7653909, 0.806895, 0.7968364, 0.7436783, 0.5880308,
  0.3476825, 0.1165299, -0.0717535, -0.1602607, 0.1945082, -0.002708793, 
    -0.09766325, 0.05541301, 0.03750932, -0.1189523, -0.06382531, 
    -0.08568406, -0.3694894, -0.1579654, -0.09165716, -0.2475982, -0.0172596, 
    0.09926081, 0.2626724, 0.4382424, 0.5168228, 0.3982515, 0.2118263, 
    0.03218746, -0.04429388, -0.03814125, 0.06189108, 0.1765723, 0.1037045, 
    -0.2136135, -0.4396877, -0.5053449, -0.3605855, -0.1262438, -0.04754913, 
    0.248708, 0.5506938, 0.5099545, 0.1252372, 0.115391, 0.04848003, 
    -0.0686264, -0.1215887, -0.3754787, -0.4117417, -0.4008203, -0.4026754, 
    -0.09124947, 0.08705425, 0.09553409, 0.1054788, 0.2125585, 0.4787207, 
    0.6396577, 0.7504815, 0.7818942, 0.7219821, 0.584938, 0.5186129, 
    0.4242442, 0.2393811, 0.09021103, 0.01102829, 0.04813743, 0.1456149, 
    0.2126722, 0.1588311, 0.1411393, 0.09125376, 0.09039116, 0.1188087, 
    0.0876565, 0.07481432, -0.05326176, -0.1616278, 0.008473396, 0.3182874, 
    0.08220328, 0.1367607, -0.1599679, -0.08195674, -0.009007692, -0.1309151, 
    -0.2606516, -0.3460194, -0.171117, 0.2974864, 0.4402112, 0.3864679, 
    0.5489686, 0.5658305, 0.6254497, 0.6206639, 0.6190848, 0.6072526, 
    0.4798274,
  0.006877899, -0.1714911, -0.2711816, -0.3843651, -0.1070222, -0.03371468, 
    -0.1249908, 0.0740653, 0.2293875, 0.0758231, -0.1595285, -0.2570546, 
    -0.2260976, -0.1286521, -0.08866215, -0.002301216, 0.06639957, 
    0.08690739, 0.2870049, 0.3214135, 0.2619891, 0.08278942, -0.03158188, 
    -0.08685589, -0.001211166, 0.03459644, 0.05201197, -0.08656263, 
    -0.2761626, -0.4914455, -0.5278544, -0.4352114, -0.4120347, -0.4627184, 
    -0.3617908, -0.1627182, -0.1096094, -0.2041078, -0.1932359, -0.04297543, 
    -0.02092171, -0.2286849, -0.4702868, -0.4828997, -0.4766665, -0.3269267, 
    -0.1027899, 0.1566672, 0.2004006, 0.1147888, 0.2199805, 0.4035578, 
    0.5370537, 0.5709563, 0.4830986, 0.4398369, 0.3868586, 0.2674901, 
    0.2077894, -0.000820756, 0.02850866, -0.03386104, -0.05366874, 
    0.08866525, 0.09942436, 0.05984092, 0.06067085, 0.05718803, -0.01576185, 
    -0.008616447, -0.04844427, -0.1076074, -0.2098374, -0.2076564, 
    -0.3203192, 0.08837247, -0.0201079, 0.1610769, 0.009270251, -0.1371976, 
    -0.1320871, -0.06180713, -0.04289436, 0.05373651, -0.1525131, 0.05108368, 
    0.3292258, 0.3937767, 0.3826764, 0.346755, 0.3654232, 0.369427, 
    0.4708428, 0.4924741, 0.36028, 0.1721454,
  -0.01221371, -0.09572601, -0.1563706, -0.327529, -0.2331287, -0.2276437, 
    -0.3533436, -0.2454498, -0.1076403, -0.06927788, -0.1621, -0.2704, 
    -0.1137276, 0.09385729, 0.1405692, 0.05526686, 0.1134701, 0.1354918, 
    0.1405697, 0.07387066, 0.03829098, -0.1083393, -0.1220117, -0.08073521, 
    -0.07650328, -0.1917548, -0.223249, -0.3403544, -0.4595764, -0.5557513, 
    -0.4475319, -0.4486227, -0.4728901, -0.3933172, -0.3331447, -0.4844307, 
    -0.5210841, -0.5624089, -0.2731678, -0.1247294, -0.5980859, -0.6740952, 
    -0.7438378, -0.6361232, -0.6738672, -0.4247293, -0.3111551, -0.1427472, 
    0.0514586, 0.1946874, 0.3455012, 0.4806409, 0.5287039, 0.4656833, 
    0.384352, 0.2726005, 0.1676526, -0.007005334, -0.1186756, -0.1259021, 
    -0.05309892, -0.03019857, 0.1320252, 0.09055376, 0.07126665, 0.01957393, 
    -0.05335951, -0.1411686, -0.2213445, -0.2617579, -0.3639717, -0.2966046, 
    -0.3893132, -0.4210186, -0.2575417, 0.0217378, 0.02953392, -0.07512093, 
    -0.2416575, -0.2558176, -0.04129931, 0.01862913, 0.1321382, 0.02723902, 
    -0.1733956, 0.1816347, 0.2619243, 0.2628675, 0.3028903, 0.2171812, 
    0.335947, 0.3458428, 0.3636489, 0.249929, 0.1537533, 0.0615983,
  0.008131504, -0.05604434, -0.1130433, -0.1340392, -0.009837627, -0.100967, 
    -0.2173409, -0.2566802, -0.2666737, -0.1756579, -0.1646872, 0.006536484, 
    0.05176783, 0.09607124, 0.2942486, 0.3222103, 0.2374444, 0.04649448, 
    -0.07554388, -0.09885049, -0.1851623, -0.2504945, -0.1766019, -0.1667051, 
    -0.1825099, -0.3484762, -0.599844, -0.4424872, -0.2214746, -0.5963774, 
    -0.4039936, -0.3326557, -0.1879296, -0.4713113, -0.527317, -0.5030334, 
    -0.2935128, -0.2578684, -0.07261443, -0.06948924, -1.12307, -1.057233, 
    -0.7911844, -0.6008849, -0.1261621, 0.3552829, 0.3762792, 0.6408949, 
    0.750237, 0.8230561, 0.7865329, 0.68554, 0.6261488, 0.3978609, 0.2323498, 
    0.05481072, -0.03366578, -0.06159544, -0.1575752, -0.08736014, 
    -0.01651073, 0.008212566, 0.0147562, -0.07904243, -0.004775047, 
    -0.09577417, -0.2127666, -0.288743, -0.3579164, -0.3890848, -0.3502178, 
    -0.340827, -0.3587787, -0.3298728, -0.1889226, 0.1142834, -0.07780647, 
    -0.2323475, -0.1981841, -0.1811268, -0.08187547, 0.01858025, -0.102188, 
    -0.1235098, -0.1273995, -0.2044015, 0.06789756, 0.3195572, 0.2747979, 
    0.3086848, 0.3892999, 0.3488216, 0.3435154, 0.1969824, 0.1177993, 
    0.04353142,
  0.1146748, 0.06963897, -0.0231185, -0.01180708, -0.05666389, -0.1389068, 
    -0.03405645, -0.06421599, -0.1689849, -0.1889877, -0.1047425, 0.1653414, 
    0.2737236, 0.3425226, 0.3471608, 0.3136487, 0.09856129, -0.007948875, 
    -0.1196837, -0.1424866, -0.0253315, -0.003928423, -0.08898711, 
    -0.2171774, -0.5114646, -0.8026755, -0.7085674, -0.06356496, -0.1678944, 
    -0.7570696, -0.2035061, -0.2558174, -0.136042, -1.330866, -1.222207, 
    -0.245759, -0.04662159, 0.008716971, -0.0761463, -0.5497785, -1.296133, 
    -0.789557, -0.2652574, 0.05240226, 0.6251559, 0.9673107, 1.013974, 
    1.194785, 1.121266, 0.9535248, 0.7629161, 0.537135, 0.3810151, 0.2460216, 
    0.1347586, 0.0975516, 0.0275158, 0.02515578, 0.06937784, 0.02927351, 
    -0.02782238, -0.0217191, -0.0336169, 0.08080411, -0.02603197, 
    -0.01856089, 0.01628613, -0.1264222, -0.2250061, -0.267812, -0.2350159, 
    -0.3477762, -0.3544006, -0.4560444, -0.4285222, -0.1448963, -0.07341194, 
    -0.09465218, -0.09074591, -0.02974331, -0.00156951, 0.127467, 0.04483372, 
    -0.3681709, -0.300007, -0.5255599, -0.1992092, 0.03352213, -0.05119419, 
    0.06286836, 0.0631125, 0.1032491, 0.1036236, 0.08685851, 0.115016, 
    0.147438,
  -0.153636, -0.09087563, -0.03446293, -0.03581427, -0.03337288, -0.01393928, 
    0.04115511, 0.05796827, -0.05949599, -0.1409412, 0.01263988, 0.3123798, 
    0.2420998, 0.3925557, 0.3631606, 0.3492775, 0.242425, 0.2582459, 
    0.2820578, 0.2273042, 0.2197368, 0.0816021, -0.1683493, -0.2801006, 
    -0.4803121, -0.6303778, -0.1270576, 0.03438428, -0.4825425, -0.960814, 
    -0.2191802, -0.06748746, -0.06037484, -1.471393, -1.575023, -0.4142159, 
    -0.0002349019, 0.110491, -0.3014872, -1.063727, -1.04859, -0.4103097, 
    -0.2453845, -0.1849842, -0.03397512, -0.1284088, -0.2749093, -0.524307, 
    -0.6671129, -0.7072822, -0.6136787, -0.3871486, -0.2369372, -0.06771517, 
    -0.08133829, -0.04055047, -0.05430365, -0.05331087, -0.02712202, 
    -0.004107714, -0.03395796, -0.03521132, -0.09976196, -0.0385313, 
    -0.1391013, -0.06714463, -0.2689681, -0.331224, -0.2994208, -0.3339252, 
    -0.3341045, -0.3226624, -0.1503804, -0.03854775, 0.1350683, -0.1036203, 
    -0.3090402, -0.2487375, -0.02757859, -0.03221726, -0.3165435, -0.3775135, 
    -0.342178, -0.3527088, -0.3401271, -0.1710346, -0.1409891, -0.4711325, 
    -0.654124, -0.583323, -0.5744691, -0.4265041, -0.3553936, -0.2618062, 
    -0.05462861, -0.05834007,
  -0.04606795, -0.01240849, 0.007789254, 0.001441538, -0.1180409, -0.1147856, 
    -0.1407948, -0.1148019, -0.09331715, -0.1459868, -0.05106461, 0.3301854, 
    0.3671813, 0.3201733, 0.06897068, 0.01150036, 0.1123476, 0.1556249, 
    0.3564708, 0.3803965, 0.2069758, 0.1383891, 0.04276705, -0.1084375, 
    -0.1858947, -0.2275455, -0.01159553, 0.02098909, -0.2386953, -0.620254, 
    -0.2963449, 0.03055942, 0.3406831, -0.6149642, -1.131956, -0.3942451, 
    -0.1356838, -0.3449126, -0.6613836, -0.7903874, -0.582494, -0.3097399, 
    -0.4102773, -0.4637765, -0.295938, -0.5705311, -0.7263254, -0.8543039, 
    -1.085342, -1.299828, -1.370515, -1.273412, -1.094066, -0.9070543, 
    -0.7845773, -0.6608791, -0.5463445, -0.354564, -0.3515198, -0.3146708, 
    -0.4877338, -0.4617085, -0.37709, -0.3241599, -0.3705792, -0.5029356, 
    -0.6592021, -0.5372782, -0.7675192, -0.7284729, -0.7407289, -0.7003486, 
    -0.5547593, -0.2380276, 0.486501, -0.05485725, -0.8631906, -0.5518786, 
    0.03938109, -0.1669992, -0.7222881, -0.7703518, -0.4785225, -0.1733143, 
    -0.0496977, 0.06846631, 0.145989, -0.0008533001, -0.2628001, -0.2595446, 
    -0.2966378, -0.1444566, -0.1851957, -0.2642643, -0.0006905198, 0.02678323,
  -0.08410501, -0.129971, -0.1064848, -0.04488003, 0.004940923, 0.3425714, 
    0.493727, 0.372047, -0.02056384, -0.003099442, 0.0851329, 0.05344439, 
    0.4602957, 0.5294514, 0.4504137, 0.04494762, -0.01885414, -0.004009962, 
    -0.04557997, -0.1353097, -0.01597378, 0.180788, 0.2575784, 0.07917643, 
    -0.07769203, -0.01341796, -0.1334381, -0.1233143, -0.09134793, 
    -0.1149964, 0.02501035, 0.1291597, -0.005345345, -0.191413, -0.2087138, 
    -0.521116, -0.4965072, -0.5146061, -0.6548893, -0.5233955, -0.3894276, 
    -0.2509022, -0.1679757, -0.1899809, 0.105299, -0.07253303, -0.123412, 
    0.03233346, -0.07049859, -0.1891509, -0.2557688, -0.3839586, -0.3431382, 
    -0.3236721, -0.3807523, -0.3240793, -0.3142323, -0.3249256, -0.395173, 
    -0.4079985, -0.5208565, -0.255915, -0.1609932, -0.128099, -0.435033, 
    -0.7272037, -0.5420967, -0.4969954, -0.8649806, -0.7841867, -0.9482492, 
    -0.8128813, -0.8500232, -1.188174, -0.3288644, -0.4634185, -0.6788317, 
    -0.88876, -1.085651, -0.6847558, -0.5449932, -0.5547918, -0.5397857, 
    -0.2908435, -0.2470932, -0.2182525, -0.06392294, -0.0002999306, 
    -0.1300038, -0.01861051, -0.03635144, -0.05659878, 0.04720974, 
    -0.0644275, -0.1034739, -0.02699256,
  0.07331663, 0.2046645, 0.2328873, 0.125107, -0.1072661, -0.1494862, 
    -0.07813199, 0.2254975, 0.1874443, 0.01595998, -0.1632882, -0.05261099, 
    0.1793225, 0.3629334, 1.099584, 0.6931877, 0.2276955, 0.09805703, 
    -0.1621653, -0.3699778, -0.1818592, 0.01796186, 0.2159438, -0.0003318787, 
    -0.1254621, 0.3203228, 0.2435639, 0.04895136, -0.02565803, 0.1874605, 
    0.7352316, 0.7795186, -0.1342511, -0.3984606, 0.1489034, -0.1821675, 
    -0.5309958, -0.674453, -0.8029044, -0.5791086, -0.405606, -0.5071684, 
    -0.5542063, -0.6101307, -0.3992583, -0.3273182, -0.3177967, -0.2963449, 
    -0.2493886, -0.2130116, -0.1519113, -0.03900421, 0.08466136, 0.06722927, 
    -0.1015043, -0.01240921, 0.190488, 0.1320406, -0.03104532, -0.0787015, 
    -0.1188058, 0.1838312, 0.1968844, 0.3030041, 0.07500929, -0.3025135, 
    -0.2918851, -0.2905669, -0.3719309, -0.4555246, -0.6762276, -0.4876047, 
    -0.5277902, -1.136595, -1.153815, -0.9033433, -0.5528389, -1.177285, 
    -1.2982, -0.8048086, -0.7291086, -0.707315, -0.4889226, -0.3205144, 
    -0.302562, -0.1866114, -0.1602437, -0.1148171, -0.0989325, -0.04097366, 
    -0.09167361, -0.3070871, 0.172226, 0.3983003, 0.1981376, 0.1523529,
  0.2122651, 0.06000277, -0.1489491, -0.03386116, -0.1561102, -0.3721583, 
    -0.6735744, -0.4183981, -0.07642293, 0.04301065, -0.5142968, -0.3425362, 
    0.2519137, 0.2067314, 0.8105569, 0.805542, 0.4836364, 0.3304954, 
    -0.1135813, -0.371003, -0.3004953, 0.08077109, 0.3941499, -0.02310228, 
    -0.4052148, 0.04519248, 0.1920828, 0.2340588, 0.2671809, 0.4216087, 
    0.9489675, 1.378476, 0.8249444, 0.02678323, 0.03514957, 0.127419, 
    -0.1910543, -0.5857973, -0.8177475, -0.6357493, -0.352546, -0.5698475, 
    -0.838093, -0.6982818, -0.3608957, -0.2556711, -0.330215, -0.5009835, 
    -0.4973053, -0.5066315, -0.4822007, -0.3477931, -0.2394761, -0.1773994, 
    -0.2351142, -0.1896222, 0.05930352, 0.1852641, -0.002935648, -0.1099997, 
    -0.1711812, 0.03189492, 0.03511763, 0.09867573, 0.09476876, -0.1675847, 
    -0.339216, -0.3247303, -0.3829334, -0.2436919, 0.1050711, 0.318271, 
    -0.02709031, -0.322891, -0.413744, -0.6338612, -0.7683824, -0.7905995, 
    -0.7370837, -0.5979237, -0.4885161, -0.4079658, -0.3048246, -0.2041407, 
    -0.130801, -0.09673476, -0.1134338, -0.03509736, 0.009954453, 0.1011329, 
    0.3018651, -0.02414346, 0.1522555, 0.3798757, 0.3272391, 0.3796316,
  0.2016857, -0.02575569, -0.8059962, -0.8307679, -0.5578845, -0.4029357, 
    -0.2443583, -0.2707911, -0.2410059, 0.3349388, 0.3387308, -0.1273179, 
    0.2421642, 0.3163996, 0.6136321, 0.4638448, 0.08065748, 0.2886326, 
    -0.3700753, -0.6126698, -0.1621327, 0.1469007, 0.293271, 0.127467, 
    -0.0644114, -0.02246797, -0.02943414, -0.0250721, 0.05500615, 0.2427342, 
    0.6992447, 1.222633, 1.559433, 1.358181, 0.9452077, 0.5941341, 0.1941824, 
    -0.2598538, -0.6885163, -0.5469633, -0.09994173, -0.3353423, -0.7011138, 
    -0.6273833, -0.242048, 0.06397402, -0.09173858, -0.3579005, -0.4835517, 
    -0.5549057, -0.4230372, -0.4268945, -0.3631576, -0.2357814, -0.2068754, 
    -0.177204, -0.09037089, 0.1015563, -0.01594019, 0.02645874, 0.09937525, 
    0.2522888, 0.3690691, 0.3121846, 0.2675231, 0.005397558, -0.2361722, 
    -0.01081428, -0.07123096, -0.1712472, -0.2167711, -0.2396388, 0.4473401, 
    0.1859304, -0.5823964, -0.6542876, -0.7250558, -0.7594959, -0.6619211, 
    -0.5446358, -0.4178455, -0.327969, -0.3450428, -0.2705636, -0.1689029, 
    -0.1723206, -0.1417215, -0.1680079, -0.09582376, -0.001845837, 0.1093192, 
    0.1599541, 0.05984092, 0.1998628, 0.1464775, 0.1381115,
  -0.130671, 0.1389253, -0.4803617, -0.8324938, -0.913581, -1.093789, 
    -0.9556053, -0.4915752, -0.2797918, 0.1122499, 0.5691671, 0.4177012, 
    0.5052502, 0.4921807, 0.9195079, 0.8329197, 0.6762139, 0.8981541, 
    -0.116153, -0.6847399, -0.1445709, 0.2054943, 0.1030529, -0.02064496, 
    -0.1226957, 0.01027948, 0.03000602, -0.2924387, -0.3044016, 0.04236054, 
    0.5394633, 0.8537209, 0.9616959, 1.435671, 1.631325, 1.385296, 0.9071544, 
    0.2835382, -0.2980212, -0.2421132, 0.0114677, -0.2449449, -0.2296782, 
    -0.1227935, -0.05510139, 0.2362071, 0.106666, -0.1218327, -0.2733953, 
    -0.4917058, -0.4207261, -0.4577053, -0.4803617, -0.3981514, -0.3099841, 
    -0.179515, -0.1556873, -0.03075147, -0.05402637, 0.08807993, 0.2771585, 
    0.4730406, 0.7348728, 0.6288023, 0.3076763, -0.07249975, -0.1071194, 
    0.2747, 0.3231701, 0.1303966, -0.266397, -0.2840402, 0.3632579, 
    0.1369884, -0.346589, -0.2975655, -0.267113, -0.3011789, -0.3495514, 
    -0.2769927, -0.295173, -0.322354, -0.2759185, -0.1875393, -0.1017808, 
    -0.1141996, -0.1516988, -0.2901266, -0.2656641, -0.2373276, -0.2817779, 
    -0.1505938, -0.07661819, 0.07806993, 0.01184213, -0.2715235,
  0.1576105, 0.223919, -0.06439503, -0.4996977, -0.8056222, -0.9614327, 
    -1.078082, -0.86415, -0.6322823, 0.03749323, 0.110898, 0.3126724, 
    0.4917741, 0.1298604, 0.3859469, 0.5111909, 0.7688735, 1.153818, 
    0.5879978, 0.05275989, 0.003231883, -0.0907948, -0.1725819, -0.2697659, 
    -0.4969144, -0.3361225, -0.2688055, -0.4973369, -0.4414132, -0.2613342, 
    0.01625371, 0.4501567, 0.679323, 1.169508, 1.576084, 1.472454, 1.07719, 
    0.5733654, 0.07727206, -0.1852282, -0.08504927, -0.06960344, 0.05892873, 
    0.3090588, 0.268564, 0.3544689, 0.3285412, 0.1733655, 0.04299462, 
    -0.2872137, -0.4255112, -0.4508369, -0.476553, -0.4268622, -0.3175365, 
    -0.1194407, -0.07931972, -0.06603885, -0.04219365, 0.1385193, 0.3977478, 
    0.6557555, 0.9189224, 0.781878, 0.3156509, 0.2391369, 0.1060477, 
    0.08661407, 0.02419548, 0.04983024, 0.2923921, 0.7703872, 0.5294528, 
    -0.05230191, -0.06568083, -0.2270415, -0.4235745, -0.2283109, -0.2044501, 
    -0.1990792, -0.2051501, -0.2729562, -0.3646228, -0.3933338, -0.2069894, 
    -0.07484436, -0.05550814, -0.1279364, -0.2124572, -0.2233138, -0.2065983, 
    -0.274437, -0.2877674, -0.1973376, 0.2469005, 0.30123,
  0.9949311, 1.081894, 0.8922456, 0.4201102, -0.4956449, -0.9838603, 
    -1.190647, -1.090046, -0.8244534, -0.1464748, -0.2413311, 0.05070925, 
    0.5938736, 0.3054619, 0.1171479, 0.02888274, 0.004762888, 0.428184, 
    0.5577567, 0.8184502, 0.5096936, -0.1742258, -0.3174384, -0.1979076, 
    -0.3678126, -0.4860411, -0.4425032, -0.3445215, 0.1266693, 0.01400673, 
    -0.2899321, -0.1588445, 0.2797954, 0.7487564, 0.9931412, 0.9168878, 
    0.7699474, 0.7164482, 0.5945242, 0.02702737, -0.1446676, 0.04891944, 
    0.1379489, 0.4732356, 0.6359793, 0.527174, 0.5229096, 0.4962658, 
    0.3784272, 0.06325799, -0.2858143, -0.4393299, -0.5652251, -0.662035, 
    -0.5491607, -0.2205962, -0.0528878, -0.05469465, -0.03265655, 0.09097695, 
    0.2662532, 0.4989028, 0.8054137, 0.7290788, 0.4298279, 0.3537691, 
    0.2608328, -0.1842192, -0.01073277, 0.3418388, 0.1880952, 0.1276622, 
    0.1311128, 0.04764926, 0.1606701, -0.0334217, -0.3396391, -0.3130277, 
    -0.2501045, -0.1630927, -0.231078, -0.307559, -0.3772203, -0.50126, 
    -0.4168201, -0.2376535, -0.1132394, -0.0403229, -0.04880238, -0.09455371, 
    -0.1522689, -0.2876692, -0.4445214, -0.3685932, -0.1434956, 0.6238701,
  -0.03154993, 0.1668223, 0.4429455, 0.6197358, 0.1005952, -0.7267969, 
    -1.130312, -1.325983, -0.8216858, -0.2505114, -0.3009174, 0.0483501, 
    0.4785414, 0.09494781, -0.1853259, -0.1201078, -0.2185776, -0.1998112, 
    -0.05274105, 0.3509209, 0.2861909, 0.03156853, 0.1005463, 0.368808, 
    0.3905529, 0.3220796, 0.2092703, 0.1356538, 0.2274344, 0.1111584, 
    -0.01974964, -0.07940125, 0.05471349, 0.3299739, 0.4250915, 0.4500589, 
    0.3428154, 0.2503511, 0.42234, 0.2277111, -0.05873013, -0.0901103, 
    -0.06563139, 0.2116961, 0.5488212, 0.648577, 0.7370863, 0.7462984, 
    0.6615653, 0.3707938, -0.09188525, -0.3180897, -0.498998, -0.769294, 
    -0.8501047, -0.5273995, -0.1933013, -0.1611561, -0.08710003, 0.08750963, 
    0.1687276, 0.2614517, 0.5298109, 0.6544533, 0.3591568, 0.6746025, 
    0.5705495, -0.01620185, 0.07343102, 0.82322, 0.7145923, 0.1587658, 
    -0.05666381, -0.04193407, -0.03846723, 0.03516552, 0.06094679, 
    -0.06763396, -0.07376987, -0.03776705, -0.2424548, -0.4009993, 
    -0.3992254, -0.4869207, -0.5091051, -0.3248278, -0.1583729, -0.1031971, 
    -0.01844776, 0.02776027, -0.02080679, -0.1704819, -0.4805732, -0.784626, 
    -0.6278384, -0.3030014,
  -0.2651274, -0.282575, -0.00425458, 0.2186779, -0.04182014, -0.3573798, 
    -0.6336168, -1.010066, -1.005036, -0.6660711, -0.641836, -0.4308335, 
    -0.2321359, -0.4802802, -0.5045471, -0.2592678, -0.1490952, -0.4479399, 
    -0.5244533, -0.1751368, 0.005884945, 0.08544222, 0.1431409, 0.071868, 
    0.1699962, 0.3495698, 0.1610281, 0.009465665, 0.009286523, 0.1462495, 
    0.1801851, 0.104127, -0.1310618, -0.1079984, 0.07191718, 0.2429621, 
    0.166074, -0.1808664, -0.2160389, -0.1041411, -0.06559956, -0.03534198, 
    -0.03576493, -0.02085614, 0.2140558, 0.5760348, 0.7848238, 0.8235117, 
    0.8206149, 0.6183848, 0.1742607, -0.1860744, -0.3915106, -0.6651925, 
    -0.9612858, -0.894603, -0.4848701, -0.2526759, -0.1181386, 0.002157629, 
    0.01140285, -0.004629135, 0.1795998, 0.3019145, 0.1840587, 0.420631, 
    0.4387302, 0.1456149, -0.02997124, 0.3825778, 0.6658787, 0.4758395, 
    0.1654718, -0.03604198, -0.1195382, -0.008649588, 0.1230074, 0.2516695, 
    0.3519299, 0.3670993, 0.1504165, -0.1346424, -0.3068914, -0.3047917, 
    -0.2558172, -0.2032292, -0.1604884, -0.0973376, -0.03985077, -0.09629606, 
    -0.04390341, 0.09419918, -0.2089586, -0.5797596, -0.6596742, -0.2438872,
  0.1763765, 0.0808363, 0.02893174, -0.06442758, -0.3446522, -0.4085192, 
    -0.3104886, -0.5371326, -0.775902, -0.6578685, -0.3508533, -0.2472726, 
    -0.1130929, -0.2131905, -0.333145, -0.1603749, -0.006224275, -0.2046127, 
    -0.45489, -0.3476307, -0.1539295, -0.02022183, 0.01281853, -0.0574777, 
    -0.1110584, -0.06618538, -0.0193592, 0.04066694, 0.04489875, 0.04253864, 
    0.1588309, 0.2103446, -0.01642952, -0.2102772, -0.1823801, -0.001178868, 
    0.1864514, 0.1411551, -0.03089893, -0.1463774, -0.2507882, -0.2107328, 
    -0.09854198, 0.01846623, 0.110719, 0.3162855, 0.5371677, 0.639609, 
    0.6198502, 0.5425715, 0.3869888, 0.09188759, -0.2112207, -0.3855691, 
    -0.5882549, -0.8342183, -0.7802308, -0.4838767, -0.1780989, 0.114886, 
    0.07663689, -0.1208394, -0.1188376, 0.02912712, 0.0905692, 0.1041108, 
    0.1136323, 0.1057058, 0.1733003, 0.2336844, 0.2331635, 0.1869886, 
    0.1408622, 0.01981735, -0.1156478, -0.1262436, -0.101976, 0.06161439, 
    0.2081312, 0.2850194, 0.2791276, 0.1644304, -0.04461884, -0.1048567, 
    -0.06831694, 0.05044961, 0.1737244, 0.2721131, 0.254746, 0.08843744, 
    0.02224243, 0.1780855, 0.06796193, -0.4033101, -0.3634834, 0.001490414,
  0.1764091, 0.2525972, 0.2061616, 0.1003836, -0.1047433, -0.2613351, 
    -0.2499744, -0.2710683, -0.5171946, -0.6595936, -0.5065336, -0.2629301, 
    -0.1848378, -0.283145, -0.4360259, -0.3572336, -0.1559315, -0.1500071, 
    -0.3144439, -0.441576, -0.487214, -0.3389719, -0.09186897, 0.05010694, 
    -0.0542388, -0.06353238, -0.06208381, 0.01389274, 0.005266443, 
    -0.1183826, -0.07601611, -0.009072751, -0.1269927, -0.2276273, 
    -0.2161852, -0.1394277, 0.004468858, 0.1010509, 0.1178477, 0.1101656, 
    0.1410898, 0.2427669, 0.3420831, 0.4742447, 0.58541, 0.6192317, 
    0.7019627, 0.7916921, 0.6933035, 0.5203873, 0.3904392, 0.1465101, 
    -0.1332254, -0.1917217, -0.2816632, -0.4697659, -0.5785389, -0.4693265, 
    -0.2073629, 0.16168, 0.2570244, 0.05468051, -0.1398345, -0.1092681, 
    0.02930617, 0.1409923, 0.1851981, 0.195631, 0.2267834, 0.2875581, 
    0.2653902, 0.1984303, 0.1360281, 0.006031394, 0.02079368, -0.009658575, 
    0.001832604, 0.05520141, 0.08482409, 0.1108494, 0.03200841, 0.06298208, 
    0.04502988, 0.1029067, 0.0555439, 0.08300161, 0.2205338, 0.2856059, 
    0.3183208, 0.3541281, 0.2874768, 0.3025973, 0.2831473, 0.02911091, 
    -0.1875069, -0.0764392,
  0.4455667, 0.6102967, 0.578753, 0.4811456, 0.3555269, 0.2444103, 0.2155855, 
    0.1532482, -0.1614979, -0.4201729, -0.3396066, -0.1451242, -0.1151437, 
    -0.171052, -0.1127022, -0.08060604, -0.1299058, -0.1135976, -0.06519258, 
    -0.2211659, -0.4774321, -0.6017647, -0.5175035, -0.2565989, -0.1395577, 
    -0.0302642, 0.01941031, 0.09032503, 0.149928, 0.1800874, 0.1240978, 
    0.006194353, -0.07663465, -0.08495167, -0.03447965, -0.007070839, 
    0.05525023, 0.08934838, 0.02709261, 0.03077096, 0.1820568, 0.3618418, 
    0.5226003, 0.7364514, 0.9532484, 1.03152, 0.9852142, 0.965146, 0.8782808, 
    0.6355562, 0.3548923, 0.09594035, -0.05166674, -0.06966758, -0.1025126, 
    -0.2463446, -0.3451724, -0.3070216, -0.07839203, 0.3130307, 0.4482193, 
    0.342474, 0.1989517, 0.169394, 0.2402273, 0.2456801, 0.3033784, 
    0.2871838, 0.2514416, 0.2967541, 0.3073498, 0.292978, 0.322861, 
    0.3528087, 0.2841564, 0.1842214, 0.09921169, 0.06880832, 0.06525993, 
    0.07701123, -0.008714616, -0.07114947, -0.1747785, -0.04453802, 
    -0.1268132, -0.2097235, -0.07140946, 0.1028748, 0.2366149, 0.3572857, 
    0.4092224, 0.404372, 0.4304783, 0.4153903, 0.2888768, 0.2543385,
  0.522162, 0.5157158, 0.4696546, 0.3999606, 0.3731054, 0.3866795, 0.4637299, 
    0.4624767, 0.2708266, 0.05886364, 0.1126233, 0.2833752, 0.3000744, 
    0.2203221, 0.2114025, 0.2024671, 0.1677178, 0.1945409, 0.2250583, 
    0.09554982, -0.1455473, -0.3110743, -0.3600979, -0.3459213, -0.1831284, 
    0.06495082, 0.1532972, 0.1467051, 0.1592052, 0.1929455, 0.165553, 
    0.0580498, -0.04575872, -0.05057675, -0.08934611, -0.1137115, 
    -0.06934279, -0.02756244, -0.01032591, -0.03695357, 0.01587838, 
    0.2185965, 0.3349864, 0.4986258, 0.7684337, 1.040683, 1.164088, 1.14358, 
    1.004632, 0.7308198, 0.3388439, 0.04372668, -0.09798884, -0.1572497, 
    -0.1990783, -0.2766337, -0.3219955, -0.2594471, -0.05451441, 0.2546487, 
    0.3986425, 0.378298, 0.3597596, 0.4859638, 0.5446055, 0.5278088, 
    0.5243094, 0.4463797, 0.3892183, 0.364316, 0.3400809, 0.3222587, 
    0.3428967, 0.3614188, 0.3926037, 0.3552338, 0.4069432, 0.3199966, 
    0.2642999, 0.2162853, 0.1143485, -0.07259814, -0.07582068, -0.1069567, 
    -0.2891181, -0.4558332, -0.3850648, -0.1219625, 0.1196065, 0.2817323, 
    0.3652284, 0.3455994, 0.2690856, 0.3038187, 0.4517841, 0.5215273,
  0.41627, 0.5664971, 0.5661066, 0.4052178, 0.1963149, 0.09958601, 0.2744073, 
    0.5404879, 0.5416433, 0.3900809, 0.3592866, 0.5199474, 0.6587496, 
    0.7702243, 0.7220473, 0.6132743, 0.5173435, 0.5086679, 0.5344659, 
    0.4592544, 0.311891, 0.1756769, 0.04449189, -0.07603192, -0.1132877, 
    -0.0167551, 0.08381498, 0.1450943, 0.2017674, 0.2506766, 0.1566011, 
    -0.02507204, -0.1340076, -0.1271067, -0.1730539, -0.2871163, -0.4107653, 
    -0.4545151, -0.4412179, -0.3604723, -0.2309642, -0.0395903, 0.03749323, 
    0.142148, 0.3448336, 0.5667576, 0.6968358, 0.6944429, 0.6004486, 
    0.4318454, 0.2166923, -0.0001860261, -0.09997444, -0.1592193, -0.2438056, 
    -0.3559151, -0.398314, -0.2566955, -0.08913422, 0.1752539, 0.4086361, 
    0.5902767, 0.6692481, 0.5893331, 0.4795994, 0.5054295, 0.5898858, 
    0.5356378, 0.4207612, 0.3325288, 0.3147717, 0.3568615, 0.1058198, 
    0.007431209, 0.04024369, 0.1972749, 0.2948334, 0.2043225, 0.1258394, 
    0.1079032, 0.09507763, 0.02587187, 0.01827097, -0.005036287, -0.240388, 
    -0.6086332, -0.8777901, -0.8631903, -0.6309147, -0.2972069, 0.02007842, 
    0.0968039, 0.01127315, -0.06983042, 0.02460313, 0.2397888,
  -0.09826446, 0.1778586, 0.358376, 0.2963798, 0.08941358, -0.08828825, 
    -0.041641, 0.1240655, 0.2207451, 0.2116629, 0.1992281, 0.2967703, 
    0.4913504, 0.6154715, 0.7272554, 0.8311455, 0.8601981, 0.8950614, 
    0.9077729, 0.8846285, 0.7530854, 0.602418, 0.4519948, 0.3171321, 
    0.2404231, 0.2065363, 0.1829358, 0.2251232, 0.2948827, 0.3251233, 
    0.2771903, 0.2094168, 0.1602632, 0.1044852, -0.005931467, -0.1744374, 
    -0.2910389, -0.355687, -0.3045805, -0.2860581, -0.2559803, -0.2198634, 
    -0.01952171, 0.2380465, 0.5119885, 0.6778256, 0.7171488, 0.7156842, 
    0.583262, 0.3305278, 0.006568432, -0.1756254, -0.1430082, -0.05018602, 
    0.00233674, -0.09502655, -0.1840077, -0.1642325, -0.02990592, -0.0574441, 
    0.1364028, 0.2733819, 0.3513122, 0.2925224, 0.2697684, 0.3128839, 
    0.4195406, 0.4452406, 0.3868583, 0.3089774, 0.2976004, 0.2148694, 
    0.1562757, 0.08267546, 0.06016588, 0.1003184, 0.2139741, 0.1791434, 
    0.04401988, 0.01623631, 0.02373981, 0.01825488, 0.06384385, 0.1727632, 
    -0.01517636, -0.4108468, -0.8904366, -1.25087, -1.343952, -1.134479, 
    -0.7511462, -0.4362533, -0.323493, -0.3495183, -0.356566, -0.2675359,
  -0.3645902, -0.2713928, -0.1340718, -0.05236685, -0.09066439, -0.1667711, 
    -0.2811757, -0.2507232, -0.2072336, -0.1399647, -0.05493864, -0.0121001, 
    0.1038179, 0.2822521, 0.5245699, 0.7402925, 0.8757417, 0.8831636, 
    0.8686941, 0.8559989, 0.8814058, 0.8871026, 0.7838308, 0.5875421, 
    0.4238216, 0.3301529, 0.250644, 0.2113538, 0.2752208, 0.3420177, 
    0.3726493, 0.358896, 0.3219819, 0.2179292, 0.06498325, -0.06945687, 
    -0.09779344, -0.05443406, 0.008505374, -0.05824274, -0.1334866, 
    -0.1763417, -0.1262274, -0.03187513, 0.1034596, 0.2913343, 0.5871189, 
    0.9211855, 1.096755, 1.010345, 0.6765721, 0.3718684, 0.1749117, 
    0.1675874, 0.2184989, 0.1951754, 0.09865838, 0.01792914, 0.00982368, 
    -0.04997456, -0.0737375, -0.0454008, 0.02894813, 0.1356701, 0.240146, 
    0.3131766, 0.3634696, 0.3695731, 0.3238699, 0.3340424, 0.3995697, 
    0.394329, 0.3380628, 0.264739, 0.2296643, 0.4213959, 0.4674085, 
    0.4693616, 0.268792, 0.1536553, 0.1904391, 0.2468355, 0.2649995, 
    0.1486258, 0.1024018, -0.1459703, -0.2580464, -0.6770902, -0.865566, 
    -0.9110096, -0.8302639, -0.6969634, -0.6271718, -0.5500884, -0.4994371, 
    -0.4505115,
  -0.5441151, -0.519587, -0.5007558, -0.4761624, -0.5193751, -0.5642644, 
    -0.6360257, -0.6544667, -0.6118559, -0.5268461, -0.4591216, -0.4306222, 
    -0.3381906, -0.1887765, 0.09484978, 0.3132905, 0.4178966, 0.4333913, 
    0.4718029, 0.5149018, 0.6012462, 0.6823498, 0.6927502, 0.6126561, 
    0.4592545, 0.3005956, 0.1426688, 0.06299764, 0.01014924, 0.08747673, 
    0.2652762, 0.3994234, 0.4924409, 0.5488212, 0.4696545, 0.3888765, 
    0.2878023, 0.2338634, 0.2055432, 0.1773693, 0.164153, 0.1286877, 
    0.02323526, -0.1619537, -0.3000233, -0.2772693, -0.06125391, 0.3346289, 
    0.7191346, 0.5632257, 0.8693125, 0.8168397, 0.6315038, 0.5849214, 
    0.4555756, 0.3607678, 0.3335216, 0.3737398, 0.3671155, 0.4231701, 
    0.3938895, 0.4132091, 0.4176362, 0.4441987, 0.4830334, 0.4755952, 
    0.4268159, 0.4223074, 0.4533784, 0.4758718, 0.5344331, 0.4426525, 
    0.2859631, 0.3639417, 0.2878672, 0.2344335, 0.4996511, 0.5452895, 
    0.4022555, 0.3833425, 0.3697358, 0.3098074, 0.1786228, 0.04353154, 
    0.04242468, -0.03228247, -0.04763055, -0.07544613, -0.02959633, 
    0.1301532, -0.1619849, -0.3941302, -0.5117255, -0.5933011, -0.5762277, 
    -0.5514556,
  -0.2993071, -0.3680572, -0.4533599, -0.5662667, -0.6966215, -0.810082, 
    -0.9073639, -0.9853747, -1.015811, -0.9774321, -0.8954985, -0.8012928, 
    -0.6597401, -0.4740304, -0.2848214, -0.1027088, -0.05702204, -0.05132526, 
    -0.007607996, 0.2549734, 0.3683848, 0.4204845, 0.484124, 0.4823336, 
    0.4029064, 0.2954031, 0.168027, 0.07639274, 0.02836213, 0.04222934, 
    0.1448335, 0.2686779, 0.4002534, 0.493271, 0.5256766, 0.4432873, 
    0.487021, 0.4574963, 0.4853771, 0.4255628, 0.2431735, 0.1806571, 
    0.06753856, -0.0605213, -0.1304595, -0.1684477, -0.1876373, -0.1367909, 
    -0.1245348, -0.06180704, -0.01371145, 0.09232712, 0.1996351, 0.2453868, 
    0.2129325, 0.1883069, 0.1510835, 0.1378022, 0.164625, 0.274456, 
    0.3735118, 0.4074312, 0.4483654, 0.4931245, 0.468922, 0.4798107, 
    0.5288991, 0.5966729, 0.6465427, 0.7309339, 0.6420181, 0.5144627, 
    0.5037529, 0.3425548, 0.3707128, 0.4146582, 0.4980397, 0.4386648, 
    0.5748141, 0.655592, 0.4342703, 0.1681083, -0.03405619, -0.09181952, 
    -0.1361721, -0.1034734, 0.0408947, 0.1591402, 0.2923279, 0.4002209, 
    0.187201, 0.1118584, 0.1580989, 0.04921198, -0.0627836, -0.190518,
  0.1508232, -0.01564819, -0.1419178, -0.2877023, -0.4441313, -0.5885161, 
    -0.7266508, -0.8091216, -0.8996489, -0.9443591, -0.9553782, -0.923054, 
    -0.8937245, -0.8776438, -0.7742093, -0.6852284, -0.5956774, -0.4857492, 
    -0.3622304, -0.256013, -0.1284739, -0.05397838, 0.07321893, 0.09488232, 
    0.1267345, 0.1012463, 0.03606072, -0.00954476, -0.01745491, 0.02608351, 
    0.05396436, 0.03625603, 0.1417736, 0.2325125, 0.323577, 0.3816825, 
    0.3901135, 0.358424, 0.316204, 0.3073172, 0.3066011, 0.2340099, 
    0.1667573, 0.1225027, 0.1137626, 0.115146, 0.1262951, 0.1317476, 
    0.1705984, 0.2434663, 0.3188733, 0.3755139, 0.3552991, 0.305885, 
    0.2282644, 0.1776298, 0.1479911, 0.1538341, 0.1721121, 0.2003835, 
    0.2396742, 0.2246837, 0.1766531, 0.1392019, 0.04367787, 0.1961356, 
    0.2240979, 0.2673274, 0.2822523, 0.3069756, 0.3427666, 0.3096611, 
    0.2928644, 0.2225192, 0.2394136, 0.2965913, 0.3513765, 0.5234143, 
    0.3650972, 0.2614188, 0.3084402, 0.2291108, 0.1261163, -0.006826401, 
    -0.1322169, -0.181322, -0.104548, 0.00583601, 0.111891, 0.2607036, 
    0.3013773, 0.1572852, -0.1776428, -0.02746367, 0.144899, 0.2933526,
  0.2370862, 0.1419201, -0.06504606, -0.2890369, -0.4553944, -0.6215565, 
    -0.7512603, -0.8207915, -0.8808339, -0.8821359, -0.8704659, -0.8490629, 
    -0.8757394, -0.8808013, -0.9059478, -0.8734933, -0.7884185, -0.6760324, 
    -0.6492584, -0.6197662, -0.5711009, -0.4662506, -0.398477, -0.3508371, 
    -0.3500233, -0.4366769, -0.4090239, -0.2997791, -0.276065, -0.237214, 
    -0.1887765, -0.08836962, -0.02474658, 0.01760368, 0.02356072, 0.05658481, 
    0.07769482, 0.09621697, 0.1017508, 0.1164481, 0.1263928, 0.1445894, 
    0.154713, 0.1592703, 0.159661, 0.1752046, 0.1925874, 0.2249605, 
    0.2614351, 0.2927339, 0.3199474, 0.3220471, 0.3186454, 0.3252697, 
    0.3302176, 0.3296642, 0.3181408, 0.2851493, 0.2550061, 0.2311617, 
    0.1928966, 0.1490816, 0.1109631, 0.05886352, 0.0224213, -0.002350569, 
    0.004940987, 0.02011037, 0.05863571, 0.077223, 0.08016884, 0.06312793, 
    0.172926, 0.1752697, 0.1812267, 0.235898, 0.2707125, 0.3091242, 
    0.3652437, 0.3759861, 0.3234966, 0.2285583, 0.1533144, 0.03869772, 
    -0.009560704, 0.005787194, 0.05832634, 0.1058201, 0.1617281, 0.1768486, 
    0.2271421, 0.2738218, 0.3127701, 0.4066337, 0.4089127, 0.3321709,
  0.2485119, 0.1177502, -0.01177457, -0.1350981, -0.264509, -0.3693429, 
    -0.4768787, -0.5680408, -0.6449614, -0.7081776, -0.765339, -0.8414132, 
    -0.8965402, -0.9422271, -0.9874418, -1.011612, -1.017113, -0.999535, 
    -0.9724516, -0.9452218, -0.91905, -0.8906482, -0.8577707, -0.8141834, 
    -0.7597075, -0.7431711, -0.7106027, -0.6902902, -0.644994, -0.59016, 
    -0.5413807, -0.4749907, -0.4199452, -0.3485259, -0.2830962, -0.2246815, 
    -0.1753976, -0.1373442, -0.1080148, -0.07738329, -0.04611702, 
    -0.01896858, 0.01543896, 0.06010043, 0.1030203, 0.1480399, 0.1860933, 
    0.2217378, 0.2554455, 0.2800223, 0.2967215, 0.3125581, 0.3309501, 
    0.3478608, 0.3519136, 0.3640718, 0.3656017, 0.3693126, 0.3630463, 
    0.352467, 0.3324963, 0.3068126, 0.2838634, 0.2667086, 0.2589449, 
    0.2323335, 0.2099216, 0.1823336, 0.1434502, 0.1054944, 0.06057245, 
    -0.0002999604, -0.07549528, -0.1143625, -0.1761952, -0.2069405, 
    -0.2225004, -0.202904, -0.09513998, -0.09906256, -0.04382169, 
    -0.02481151, -0.01359749, -0.02674848, -0.02500707, -0.007933408, 
    0.02453728, 0.05801709, 0.1190197, 0.2282645, 0.3262953, 0.4127211, 
    0.4707451, 0.4840752, 0.4316988, 0.3605886,
  0.06770134, 0.003557459, -0.05301806, -0.1167388, -0.179727, -0.2483306, 
    -0.3186268, -0.3854237, -0.4537342, -0.5189035, -0.5740467, -0.6318755, 
    -0.6860259, -0.7405018, -0.7944406, -0.8425525, -0.8852772, -0.9233143, 
    -0.9506906, -0.9664295, -0.9694244, -0.9568266, -0.9360096, -0.9079171, 
    -0.8744861, -0.8338937, -0.7922108, -0.7449126, -0.6925688, -0.6412668, 
    -0.5816802, -0.5252186, -0.4721099, -0.4065662, -0.3499419, -0.2950103, 
    -0.2404855, -0.1801502, -0.125186, -0.0732329, -0.02077523, 0.02818312, 
    0.07386996, 0.1181245, 0.1609956, 0.2029878, 0.2374116, 0.2704032, 
    0.3011649, 0.3316499, 0.364967, 0.3939546, 0.4133068, 0.4293061, 
    0.4408296, 0.4440686, 0.4453381, 0.4490001, 0.4433198, 0.4384044, 
    0.4368907, 0.4245698, 0.4146251, 0.4007742, 0.3858002, 0.3667735, 
    0.342099, 0.3134207, 0.279241, 0.2464448, 0.2102469, 0.1744722, 
    0.1330008, 0.09869093, 0.06218376, 0.03555616, 0.01166293, -0.001895014, 
    -0.012979, -0.01908251, -0.01379281, -0.006582513, 0.002776206, 
    0.0154878, 0.0381766, 0.06119092, 0.08309847, 0.1033784, 0.1232352, 
    0.1397717, 0.1484142, 0.1551851, 0.1570568, 0.147812, 0.1279064, 0.1028576,
  0.1631947, 0.1519809, 0.1401968, 0.128428, 0.1159763, 0.1022234, 
    0.08751011, 0.07071304, 0.05119991, 0.03033352, 0.007025242, -0.0167532, 
    -0.04214382, -0.06759977, -0.09229088, -0.1164443, -0.1393449, 
    -0.1619201, -0.1843157, -0.2071348, -0.2310768, -0.2562233, -0.2839251, 
    -0.3134173, -0.344358, -0.3757545, -0.4057839, -0.433274, -0.456923, 
    -0.4752011, -0.4881401, -0.4952202, -0.4967332, -0.4926162, -0.4832416, 
    -0.4697957, -0.4529338, -0.4328666, -0.4105191, -0.3864636, -0.3612347, 
    -0.3358126, -0.3103075, -0.285862, -0.2615929, -0.2388391, -0.2188692, 
    -0.2156301, -0.1990285, -0.1773973, -0.1601448, -0.1501832, -0.1543837, 
    -0.1591034, -0.1847553, -0.1450253, -0.139751, -0.122386, -0.1735411, 
    -0.1360245, -0.1024306, -0.08584571, -0.05168223, -0.04224181, 
    -0.02837467, -0.01520753, -0.001226425, 0.01060653, 0.02219486, 
    0.05256605, 0.07854271, 0.1057074, 0.1314723, 0.1450627, 0.1834414, 
    0.2076437, 0.2272732, 0.233458, 0.2615993, 0.2719505, 0.2792261, 
    0.2839949, 0.2865827, 0.285541, 0.2811627, 0.2764915, 0.2704043, 
    0.263422, 0.2546817, 0.2448184, 0.2341576, 0.2225368, 0.2108505, 
    0.1984971, 0.1862087, 0.1741805,
  0.08568811, 0.1033154, 0.1261001, 0.1487751, 0.1635356, 0.1664171, 
    0.1595325, 0.1440699, 0.1226015, 0.09859467, 0.07639432, 0.05544662, 
    0.03316498, 0.008034468, -0.01973248, -0.04922462, -0.07832611, 
    -0.1024961, -0.1179258, -0.127903, -0.1338763, -0.1390033, -0.1454649, 
    -0.1536843, -0.1697811, -0.1937722, -0.2231989, -0.2557836, -0.2870498, 
    -0.3144588, -0.3366108, -0.350739, -0.3549366, -0.3475142, -0.3282437, 
    -0.2977104, -0.2567921, -0.2065639, -0.1494837, -0.09333134, -0.05221939, 
    0.001670837, 0.04003429, 0.1006131, 0.1157503, 0.1252384, 0.1289821, 
    0.117116, 0.1143827, 0.1115344, 0.1120546, 0.0838809, 0.1022403, 
    0.09377694, 0.07745183, 0.1151798, 0.1111107, 0.08145571, 0.08270896, 
    0.07121807, 0.03772199, 0.001019478, -0.03001881, -0.0548234, 
    -0.08289981, -0.107672, -0.1225808, -0.1296772, -0.1297585, -0.1034727, 
    -0.0571509, -0.01566339, 0.0218854, 0.06485438, 0.08425546, 0.1047311, 
    0.09839964, 0.101069, 0.06125736, 0.09286523, 0.07976317, 0.08710337, 
    0.1089622, 0.1401147, 0.1579694, 0.175629, 0.1938418, 0.1971784, 
    0.1906846, 0.1732204, 0.1508088, 0.1260366, 0.1017356, 0.08353949, 
    0.07128382, 0.07180452,
  0.3279238, 0.3274851, 0.3086693, 0.2606063, 0.189024, 0.09735739, 
    0.005007148, -0.06178972, -0.07380146, -0.03018165, 0.05743229, 
    0.1599226, 0.2503524, 0.3076117, 0.3283148, 0.3170843, 0.2771266, 
    0.219249, 0.1505964, 0.0746361, 0.003005186, -0.05467713, -0.08804291, 
    -0.09154236, -0.06571226, -0.02568948, -0.01218033, -0.03472269, 
    -0.0928607, -0.1801, -0.2827857, -0.3790421, -0.4502823, -0.4859266, 
    -0.4882536, -0.4621148, -0.4052463, -0.3251514, -0.2279029, -0.1260309, 
    -0.02720261, 0.1127706, 0.1664176, 0.2401962, 0.2082949, 0.2081647, 
    0.2015729, 0.221918, 0.256651, 0.2799746, 0.2819928, 0.2657981, 
    0.2462018, 0.2349063, 0.2348086, 0.2183047, 0.1801049, 0.1449324, 
    0.1149356, 0.08671284, 0.04769945, -0.01147985, -0.08939314, -0.1623745, 
    -0.2247291, -0.2693903, -0.2899473, -0.2851132, -0.265761, -0.2447324, 
    -0.2383847, -0.2495172, -0.25912, -0.2695689, -0.3227262, -0.3580132, 
    -0.4334683, -0.4640999, -0.4187226, -0.3438048, -0.2479224, -0.1349504, 
    -0.001812458, 0.07756573, 0.2004824, 0.2675072, 0.3070742, 0.309841, 
    0.3022239, 0.3394964, 0.2833276, 0.2695584, 0.2540479, 0.2513785, 
    0.2736607, 0.3059516,
  0.5712832, 0.5039167, 0.4284284, 0.3624453, 0.284353, 0.176931, 0.06999755, 
    -0.00549078, -0.02621007, 0.02605247, 0.1373634, 0.26894, 0.3901153, 
    0.494884, 0.5724721, 0.5662861, 0.4890568, 0.3284938, 0.1561302, 
    0.02178774, -0.04102147, -0.01733947, 0.0432725, 0.08628988, 0.08803129, 
    0.1068464, 0.146397, 0.167491, 0.108995, 0.003118992, -0.1084368, 
    -0.1831602, -0.2096087, -0.2076719, -0.1870664, -0.1673887, -0.1533751, 
    -0.1254776, -0.06159401, 0.01819181, 0.1052513, 0.1745563, 0.3057404, 
    0.4236765, 0.5269313, 0.6302354, 0.4711044, 0.4963648, 0.5029407, 
    0.4570253, 0.3718691, 0.304942, 0.2591739, 0.2341252, 0.2100202, 
    0.1789655, 0.08422279, -0.006988287, -0.1169492, -0.1433653, -0.1337298, 
    -0.1394265, -0.1307025, -0.1382057, -0.2260799, -0.3565651, -0.4407773, 
    -0.5023167, -0.5313857, -0.5285211, -0.5150928, -0.5174851, -0.5426326, 
    -0.5907443, -0.659348, -0.7347062, -0.7330461, -0.6700091, -0.5169492, 
    -0.4635471, -0.3049862, -0.08184183, 0.1076602, 0.2530378, 0.3554465, 
    0.4321067, 0.475336, 0.4539329, 0.4547956, 0.4863385, 0.4694115, 
    0.4803002, 0.6179142, 0.6725852, 0.6699159, 0.6347922,
  0.2858179, 0.2026799, 0.1522729, 0.09654379, 0.02385569, -0.0324111, 
    -0.1450572, -0.2184615, -0.06753445, -0.08691835, -0.01981306, 
    0.03596449, 0.1128199, 0.174099, 0.2418239, 0.2522736, 0.1362906, 
    0.050776, -0.01327133, -0.08724546, -0.1832741, -0.1090388, 0.03218842, 
    0.1404893, 0.2358991, 0.3518984, 0.3533635, 0.2295027, 0.0879674, 
    -0.03410387, -0.1399636, -0.1916234, -0.1992245, -0.1995177, -0.1995988, 
    -0.2177954, -0.2390833, -0.2555389, -0.233079, -0.164784, -0.04658699, 
    0.1226516, 0.2913699, 0.4122505, 0.4231553, 0.4588978, 0.3802841, 
    0.3274357, 0.2426698, 0.140554, 0.04830146, 0.008864641, 0.04154688, 
    0.1126406, 0.1608827, 0.164252, 0.0957298, -0.008518249, -0.1094135, 
    -0.1388406, -0.1408426, -0.1140032, -0.1038632, -0.1115291, -0.1823789, 
    -0.273069, -0.3226132, -0.3501197, -0.364931, -0.3822486, -0.2734271, 
    -0.264166, -0.3038307, -0.4098365, -0.5272194, -0.5839739, -0.6052142, 
    -0.4663796, -0.3817767, -0.2289445, -0.06291282, 0.1198183, 0.2648379, 
    0.3496199, 0.4069928, 0.4501732, 0.4497826, 0.4364036, 0.4389753, 
    0.4861596, 0.5694115, 0.5664167, 0.5227481, 0.4918886, 0.4191673, 
    0.3584903,
  0.1326602, 0.05132884, -0.02004153, -0.04601824, -0.0303607, 0.007774115, 
    0.03952909, 0.128917, 0.07118559, 0.05687904, 0.05388415, 0.04680389, 
    0.03939843, 0.08921957, 0.1660264, 0.2020297, -0.00182724, -0.06436014, 
    0.02458763, 0.1193628, 0.1891544, 0.1895449, 0.2008893, 0.2330996, 
    0.2723253, 0.2571878, 0.1760693, 0.0661726, -0.0443573, -0.1297898, 
    -0.209934, -0.2536027, -0.251096, -0.241672, -0.2179909, -0.2374401, 
    -0.261138, -0.2815008, -0.2748747, -0.1741095, 0.00188303, 0.11448, 
    0.2393661, 0.2979441, 0.211827, 0.2035425, 0.1440861, 0.02222729, 
    -0.1266661, -0.2700906, -0.3192929, -0.2808164, -0.1652403, -0.01117125, 
    0.07056704, 0.05712302, -0.01003194, -0.09349543, -0.1759987, -0.2439511, 
    -0.2734922, -0.3111387, -0.368349, -0.4424213, -0.4851296, -0.5117409, 
    -0.4984923, -0.4724994, -0.4290913, -0.4205951, -0.4724669, -0.5511941, 
    -0.6642475, -0.7360572, -0.7017473, -0.584267, -0.4300189, -0.2471738, 
    -0.09336527, 0.04940818, 0.169444, 0.3023867, 0.4271588, 0.4970156, 
    0.4927838, 0.4727155, 0.4562441, 0.4410423, 0.4897076, 0.5556419, 
    0.560541, 0.5059349, 0.425108, 0.3181908, 0.252924, 0.1944115,
  0.06288475, -0.04084247, -0.1214089, -0.1586972, -0.1663633, -0.1594949, 
    -0.1612037, -0.2118223, -0.2615131, -0.2636452, -0.212278, -0.1702533, 
    -0.1328184, -0.1026589, -0.1595598, -0.2908912, -0.434413, -0.4574111, 
    -0.3475645, -0.1964574, -0.09243751, -0.01761651, 0.02551496, 0.00997138, 
    -0.01548433, -0.007297516, -0.06636333, -0.1307673, -0.1965553, 
    -0.2084043, -0.2281146, -0.264703, -0.2680722, -0.2745502, -0.3998103, 
    -0.4460831, -0.4602757, -0.4042702, -0.3531635, -0.287392, -0.2253802, 
    -0.2148659, -0.2009661, -0.172955, -0.1507871, -0.1833066, -0.2512266, 
    -0.3589089, -0.491754, -0.5754779, -0.6034239, -0.4918027, -0.3515033, 
    -0.308502, -0.2942604, -0.3560443, -0.4016009, -0.4028217, -0.3963275, 
    -0.4184955, -0.4933164, -0.5902565, -0.6909727, -0.7126685, -0.6778055, 
    -0.5945047, -0.5278217, -0.5052468, -0.6153217, -0.6916889, -0.7923887, 
    -0.8617246, -0.9267638, -0.8930561, -0.6593646, -0.3314838, -0.05462825, 
    0.05780679, 0.06879282, 0.08314842, 0.1285098, 0.1975853, 0.2721784, 
    0.3153262, 0.3062604, 0.2704533, 0.2258895, 0.1990989, 0.2225202, 
    0.2756452, 0.2919538, 0.2357526, 0.1281679, 0.07260154, 0.1041933, 
    0.1130312,
  -0.1579485, -0.1924375, -0.2232969, -0.2585996, -0.2919654, -0.3077695, 
    -0.3570209, -0.4336645, -0.4915097, -0.5447487, -0.5678607, -0.5360736, 
    -0.5104389, -0.5080788, -0.5713601, -0.6390195, -0.6769426, -0.6581438, 
    -0.5594296, -0.4740618, -0.4296445, -0.4005756, -0.4234759, -0.4689674, 
    -0.5096738, -0.5475644, -0.5992083, -0.6786191, -0.7489153, -0.7829811, 
    -0.8085019, -0.8988014, -1.021148, -1.16957, -1.311985, -1.209544, 
    -0.9092833, -0.7590715, -0.5781797, -0.5419493, -0.6347389, -0.6878802, 
    -0.7859596, -0.8565489, -0.9438047, -0.9296445, -0.9280981, -0.9314834, 
    -0.8623757, -0.8423073, -0.7333879, -0.6301653, -0.5419167, -0.4522195, 
    -0.5573465, -0.6557676, -0.7008034, -0.7470599, -0.5459205, -0.5721738, 
    -0.8038307, -0.9231015, -1.042617, -0.9979063, -0.9826556, -0.996474, 
    -0.9559141, -1.028408, -1.099778, -1.139134, -1.134934, -1.136562, 
    -1.163645, -1.073329, -0.8443255, -0.5981992, -0.4618223, -0.5780821, 
    -0.6366433, -0.5384336, -0.5049049, -0.4101784, -0.2769265, -0.04909444, 
    0.06158268, 0.1719505, 0.2258079, 0.2033633, 0.1198834, 0.06242919, 
    0.05248439, 0.01836979, -0.04636002, -0.08763593, -0.1154356, -0.1240131,
  -0.3997618, -0.4180073, -0.4488339, -0.5070208, -0.5698137, -0.465403, 
    -0.4281307, -0.519765, -0.6652403, -0.9460181, -1.056158, -1.108649, 
    -1.140126, -1.072337, -1.058697, -1.10707, -1.155377, -1.139133, 
    -1.004384, -0.8850645, -0.8313372, -0.7344786, -0.7533913, -0.796181, 
    -0.795058, -0.7473041, -0.7657123, -0.7798562, -0.7962624, -0.8723366, 
    -1.015045, -1.238271, -1.318105, -1.187945, -0.9589572, -0.7616918, 
    -0.6336482, -0.5987036, -0.7214572, -1.012521, -1.316688, -1.548084, 
    -1.59981, -1.54701, -1.476731, -1.44382, -1.375543, -1.331923, -1.292665, 
    -1.324094, -1.286513, -1.188238, -1.194358, -1.282932, -1.363255, 
    -1.330068, -1.185455, -0.9712298, -0.79081, -0.672711, -0.6721412, 
    -0.7933977, -0.8449277, -0.777675, -0.6671282, -0.6584044, -0.7861712, 
    -0.9926815, -1.197451, -1.298557, -1.314979, -1.289589, -1.287343, 
    -1.288303, -1.265452, -1.217698, -1.108485, -0.975087, -0.816949, 
    -0.6724015, -0.5014381, -0.2965878, -0.1140684, 0.04006577, 0.0805769, 
    0.04600656, 0.0562768, 0.05167067, 0.02932358, -0.02277613, -0.04217708, 
    -0.06252217, -0.1134011, -0.2307676, -0.3206764, -0.3710182,
  -1.175575, -1.024664, -0.9731989, -0.9001195, -0.7631567, -0.6775608, 
    -0.759413, -0.924387, -1.092762, -1.115614, -1.052398, -1.082818, 
    -1.195237, -1.293658, -1.364036, -1.400885, -1.350396, -1.157639, 
    -0.9619526, -0.9486549, -1.095628, -1.188905, -1.255361, -1.154531, 
    -0.9917539, -0.798362, -0.8117898, -0.9303119, -0.9526262, -0.9229711, 
    -0.9647353, -1.023166, -0.9593639, -0.775461, -0.666688, -0.7216687, 
    -0.8684297, -1.079953, -1.340126, -1.594748, -1.758794, -1.777886, 
    -1.744731, -1.629514, -1.444634, -1.354741, -1.451372, -1.623019, 
    -1.737717, -1.709576, -1.519911, -1.244927, -1.162555, -1.261774, 
    -1.18871, -0.9067929, -0.6124568, -0.4146218, -0.2642148, -0.1937721, 
    -0.2870013, -0.5264869, -0.6244035, -0.5113502, -0.3923073, -0.4771216, 
    -0.7246312, -0.9827368, -1.167681, -1.224371, -1.175185, -1.171246, 
    -1.271425, -1.394293, -1.439507, -1.341216, -1.058859, -0.6997936, 
    -0.3930395, -0.2088113, -0.18399, -0.05352116, 0.1030376, 0.1454697, 
    0.1323998, 0.1533308, 0.1856225, 0.08171606, -0.1085997, -0.1995827, 
    -0.2839414, -0.4352435, -0.6183652, -0.8584043, -1.075445, -1.160178,
  -1.014508, -0.8196833, -0.7303767, -0.6328669, -0.5665095, -0.6074438, 
    -0.760422, -0.8146539, -0.7344458, -0.671783, -0.7242894, -0.8790257, 
    -1.054644, -1.154872, -1.14579, -1.060748, -0.9342501, -0.8127172, 
    -0.7772355, -0.7804258, -0.7051816, -0.5763404, -0.5009011, -0.4624245, 
    -0.465403, -0.5696999, -0.7412817, -0.8184135, -0.8015356, -0.7833874, 
    -0.8341525, -0.7996793, -0.6642303, -0.5967011, -0.6929412, -0.871408, 
    -1.034755, -1.14395, -1.252984, -1.382037, -1.448654, -1.417258, 
    -1.437114, -1.472271, -1.432443, -1.450949, -1.663628, -1.860292, 
    -1.724224, -1.405783, -1.015208, -0.6307349, -0.5150933, -0.6396701, 
    -0.5417049, -0.09940362, 0.2537863, 0.2935164, 0.1954043, 0.0007429123, 
    -0.1770892, -0.3084531, -0.2695858, -0.1528215, -0.1837461, -0.3392308, 
    -0.4363015, -0.5786839, -0.8463597, -1.059608, -1.168072, -1.255735, 
    -1.310129, -1.268772, -1.124354, -0.8999724, -0.6012096, -0.323313, 
    -0.1543188, -0.1612363, -0.1942606, -0.1255918, 0.01034594, 0.1107366, 
    0.1675072, 0.217263, 0.2321882, 0.1311953, -0.04212832, -0.1450416, 
    -0.2500709, -0.4817441, -0.7691302, -1.001666, -1.184267, -1.204042,
  -0.6791396, -0.5854874, -0.521848, -0.4911678, -0.5091367, -0.4676814, 
    -0.300559, -0.1035213, -0.04954982, -0.1449926, -0.3249893, -0.5231011, 
    -0.7249892, -0.7994034, -0.7402887, -0.6783745, -0.7167861, -0.7656794, 
    -0.7236059, -0.5653539, -0.3999245, -0.3594947, -0.4265032, -0.4838762, 
    -0.5637424, -0.6387913, -0.6112852, -0.556695, -0.5724008, -0.6062875, 
    -0.5690808, -0.4541068, -0.3945031, -0.4957085, -0.608778, -0.6542206, 
    -0.7347217, -0.8475637, -0.8835664, -0.984494, -1.18163, -1.164833, 
    -1.073655, -1.151877, -1.179709, -1.065338, -1.115582, -1.235585, 
    -1.070139, -0.6261938, -0.1987526, 0.05837631, 0.1605411, 0.2359316, 
    0.4906843, 0.8391054, 0.8319278, 0.5375432, 0.2990341, 0.1525168, 
    0.115961, 0.1427839, 0.1906517, 0.1358178, -0.003244638, -0.1424537, 
    -0.2406309, -0.4518285, -0.8111873, -1.024924, -0.9618709, -0.8120499, 
    -0.7269914, -0.6983778, -0.5814836, -0.2482963, 0.1224232, 0.2321885, 
    0.2567649, 0.1252708, -0.08376193, -0.1073461, 0.1152124, 0.3715436, 
    0.4794374, 0.4472597, 0.34337, 0.2016217, 0.0003033876, -0.1777564, 
    -0.3619524, -0.6577045, -0.8869687, -0.9628475, -0.9781468, -0.8536189,
  -0.3106663, -0.2691948, -0.178391, -0.1283422, -0.07287359, 0.2462347, 
    0.5337994, 0.5563908, 0.3475204, 0.01950908, -0.3070209, -0.6249245, 
    -0.8220271, -0.8586806, -0.8187068, -0.7863991, -0.786562, -0.7249407, 
    -0.5846087, -0.5412657, -0.5985899, -0.6621966, -0.6922419, -0.652854, 
    -0.642242, -0.5644591, -0.4004774, -0.3411021, -0.2673879, -0.06870651, 
    0.123579, 0.1664338, 0.03782082, -0.1555552, -0.2381072, -0.2138724, 
    -0.2124243, -0.291477, -0.3027561, -0.3568418, -0.6127009, -0.704514, 
    -0.6339738, -0.7560766, -0.8724827, -0.7322649, -0.5839083, -0.6414773, 
    -0.6548724, -0.2420306, 0.2782819, 0.6688094, 0.8186952, 0.863959, 
    0.9895449, 1.046592, 0.7620385, 0.4696068, 0.4049745, 0.3738223, 
    0.3969342, 0.4485943, 0.4151309, 0.3451765, 0.2250593, 0.06864643, 
    -0.1193089, -0.2811904, -0.3769586, -0.3752172, -0.3349991, -0.2810278, 
    -0.2278214, -0.1585505, 0.0409286, 0.64114, 1.172065, 0.9138775, 
    0.3560489, 0.04512763, -0.1792865, -0.05910397, 0.3513614, 0.6306094, 
    0.7470319, 0.8001407, 0.7074487, 0.4494734, 0.09844792, -0.1781471, 
    -0.3103086, -0.4227598, -0.4168679, -0.3926491, -0.4687722, -0.4087462,
  -0.1072974, 0.01609135, 0.1584251, 0.285167, 0.5157819, 0.7576114, 
    0.6330996, 0.3726993, 0.08736396, -0.5201719, -1.089312, -1.353505, 
    -1.262799, -1.00619, -0.8981503, -0.8311908, -0.7340389, -0.6282933, 
    -0.500494, -0.5508847, -0.5684626, -0.4309785, -0.3338597, -0.2700901, 
    -0.1974828, -0.03822184, 0.1700139, 0.3216579, 0.5852644, 0.772439, 
    0.6713159, 0.4582949, 0.2025168, 0.1474876, 0.2500591, 0.2628198, 
    0.3159933, 0.335655, 0.1950626, -0.05160069, -0.3968971, -0.7176166, 
    -0.6355364, -0.5472715, -0.5681698, -0.3727597, -0.1087135, -0.01060152, 
    0.06251049, 0.26308, 0.7765239, 1.186827, 1.271544, 1.198871, 1.04892, 
    0.891075, 0.6760033, 0.5203229, 0.4359154, 0.43642, 0.591612, 0.7089136, 
    0.7197858, 0.6902937, 0.4962833, 0.308718, 0.2425399, 0.2173283, 
    0.1788354, 0.06553817, 0.02935624, 0.020437, 0.1372013, 0.4327253, 
    0.717377, 1.353721, 1.903607, 1.17877, 0.159597, -0.1853737, -0.05433524, 
    0.3265404, 0.7953392, 0.9827253, 0.9977155, 0.9194929, 0.5386823, 
    0.1643659, -0.1182839, -0.303082, -0.3097714, -0.2711159, -0.2078508, 
    -0.2377663, -0.4308001, -0.3392146,
  0.3722923, 0.4964623, 0.6161075, 0.7049583, 0.885834, 0.8394473, 0.5980736, 
    0.4688093, -0.07253188, -0.842226, -0.9697809, -0.6636126, -0.5228574, 
    -0.4546933, -0.4391003, -0.2051978, 0.06304789, 0.0818789, 0.165082, 
    0.2611107, 0.2922467, 0.3663353, 0.3774682, 0.4426212, 0.5288841, 
    0.7448672, 1.045372, 1.216498, 1.259223, 1.120811, 0.9508241, 0.7345481, 
    0.4274192, 0.4046491, 0.4911237, 0.4048607, 0.3694115, 0.2443138, 
    -0.07389891, -0.3304095, -0.543707, -0.7717344, -0.5668353, -0.1998268, 
    0.01812565, 0.2205182, 0.2459251, 0.2366966, 0.4200137, 0.7417423, 
    1.322732, 1.648952, 1.444542, 1.192198, 0.9978783, 0.8237898, 0.6473249, 
    0.413959, 0.3171979, 0.4982364, 0.8948184, 1.059288, 1.014057, 0.9343204, 
    0.6375105, 0.508588, 0.4815861, 0.3935652, 0.3408797, 0.2700299, 
    0.3717226, 0.3243756, 0.2784284, 0.6538028, 0.9208925, 1.362852, 
    1.599881, 0.6722761, -0.2123919, -0.1497129, 0.4411236, 0.8076113, 
    1.094444, 1.125255, 0.8813906, 0.5671979, 0.04861069, -0.1523496, 
    -0.1635312, -0.3592018, -0.373899, -0.2328835, -0.1547911, -0.1450742, 
    -0.09424412, 0.1256614,
  0.595746, 0.605707, 0.6381127, 0.8394315, 0.9783802, 0.7646267, 0.530349, 
    0.3971132, -0.08431578, -0.492226, -0.2831438, -0.05632102, -0.3312883, 
    -0.3070371, 0.03614318, 0.3487898, 0.6086855, 0.6423119, 0.7539167, 
    0.8444278, 0.7464622, 0.7074323, 0.7378848, 0.8393984, 0.8183372, 
    0.9184999, 1.089756, 1.143663, 1.102387, 1.124409, 1.155203, 0.7605246, 
    0.3650169, 0.3873313, 0.2717389, 0.1473574, 0.1218854, -0.03905207, 
    -0.3600808, -0.6187559, -0.4810931, -0.2384987, 0.01999742, 0.3186139, 
    0.3785911, 0.4372337, 0.4606549, 0.5102805, 0.9162213, 1.268354, 
    1.574864, 1.540766, 1.028949, 0.800222, 0.7596459, 0.6086205, 0.3552513, 
    0.197097, 0.5023867, 0.8848087, 1.157302, 1.234532, 1.12947, 0.9704369, 
    0.6322044, 0.5543076, 0.5274682, 0.4243269, 0.4897403, 0.3610455, 
    0.3118269, 0.212429, 0.2617942, 0.6524681, 0.8390243, 1.119999, 
    0.8612099, 0.02872133, -0.2328836, 0.2440859, 0.8942814, 0.9052513, 
    0.8727643, 0.7350364, 0.3117618, 0.01529372, -0.1999896, -0.2392306, 
    -0.3067441, -0.4308326, -0.286936, 0.06368232, 0.238959, 0.2165307, 
    0.3342878, 0.5204368,
  0.6380804, 0.5854113, 0.6839471, 0.9017363, 0.7818308, 0.3989687, 
    -0.03968689, -0.2557676, 0.009792328, 0.1647403, 0.06234763, 0.133653, 
    -0.3122455, -0.5747452, 0.06934619, 0.5817326, 0.7464297, 0.8037539, 
    0.8468855, 0.6363874, 0.3713159, 0.3088158, 0.3237084, 0.3918724, 
    0.4290631, 0.5964297, 0.7107854, 0.7643988, 0.7783637, 0.9062777, 
    0.8880162, 0.2982202, 0.003900528, 0.1507266, -0.03060484, -0.01729103, 
    -0.06320572, -0.2320207, -0.3814999, -0.4673398, 0.04784572, 0.6596622, 
    0.6569765, 0.8058209, 0.7425885, 0.623513, 0.7452741, 0.7772077, 
    0.9150332, 0.9617454, 0.8963482, 0.6920188, 0.3036562, 0.2371849, 
    0.2759057, 0.24433, 0.2910097, 0.433897, 0.8429303, 1.071674, 1.077224, 
    1.073155, 0.9101342, 0.7488548, 0.5314558, 0.4932234, 0.4660912, 
    0.3231551, 0.3343365, 0.186013, 0.1042096, 0.1925071, 0.3397566, 
    0.5252707, 0.6448517, 0.7482367, 0.1454539, -0.3018938, -0.2249408, 
    0.2100527, 0.8220811, 0.6652774, 0.4947207, 0.4115826, 0.02751696, 
    -0.3235407, -0.5223684, -0.4850645, -0.4345596, -0.1140521, 0.1598249, 
    0.2839948, 0.405349, 0.3732363, 0.4267357, 0.5854108,
  0.5740023, 0.4956656, 0.6255808, 0.5944777, 0.1522729, -0.05205667, 
    -0.1583718, -0.03610611, 0.3368105, 0.1866477, -0.1887428, 0.4005315, 
    0.0592227, -0.5840552, 0.1210227, 0.5448997, 0.6199323, 0.5505149, 
    0.4535749, 0.1665957, 0.008181095, 0.06975317, 0.07839584, 0.182986, 
    0.2381291, 0.3640404, 0.4205513, 0.5006294, 0.558198, 0.5563111, 
    0.4336386, -0.023736, -0.1935606, -0.1719947, -0.2534075, -0.08133733, 
    -0.1134174, -0.2726622, -0.280914, -0.04605079, 0.6517683, 1.004698, 
    0.7715604, 0.7736275, 0.810997, 0.7807233, 0.848074, 0.6122992, 
    0.3617618, 0.3344179, 0.165375, -0.07717049, -0.1860572, -0.03908467, 
    0.2494895, 0.5141218, 0.8043561, 1.007888, 1.044607, 0.9873477, 
    0.8406354, 0.761371, 0.7100528, 0.6931093, 0.5077578, 0.2877057, 
    0.2440534, 0.1903912, 0.2000756, 0.1151471, 0.09970117, 0.1572044, 
    0.1920514, 0.3310328, 0.4874949, 0.5114202, -0.02878094, -0.1093808, 
    -0.2488339, 0.001328766, 0.6768987, 0.4173444, 0.3411074, 0.4483177, 
    0.2220156, -0.4029675, -1.079156, -0.5983293, -0.2619524, 0.02873778, 
    0.2475364, 0.230186, 0.2420839, 0.2941511, 0.4135685, 0.5223415,
  0.3806591, 0.2647896, 0.2591906, -0.01416492, 0.01576567, -0.05731383, 
    -0.07248306, 0.1449975, 0.08747786, -0.08587827, -0.2840553, 0.07258558, 
    -0.1768938, -0.007151067, 0.6093041, 0.4517845, 0.4224224, 0.3845487, 
    0.2482204, 0.05665112, 0.03422284, 0.08279061, -0.01084566, 0.01096439, 
    0.05744934, 0.112967, 0.1428661, 0.2076941, 0.2190704, 0.2218223, 
    0.1387968, -0.2205627, -0.1991594, -0.1904192, -0.209446, -0.1814349, 
    -0.1485247, -0.06141543, 0.04094464, 0.4496036, 0.7799584, 0.7935655, 
    0.6327584, 0.6132598, 0.6647575, 0.565506, 0.415066, 0.06002045, 
    -0.2071183, -0.2459207, -0.3148496, -0.2251848, 0.09919643, 0.5143332, 
    0.9620222, 1.174538, 1.177859, 1.147553, 1.01614, 0.9363059, 0.8093692, 
    0.7669212, 0.7652448, 0.5859316, 0.3096295, 0.1958437, 0.1944766, 
    0.1899356, 0.1841738, 0.1564395, 0.1758244, 0.2168889, 0.2819934, 
    0.2893829, 0.1658149, 0.1072054, -0.2481503, -0.04878515, -0.1506406, 
    -0.03578061, 0.2833927, 0.1512637, 0.1706322, 0.147862, 0.07510817, 
    -0.4943255, -1.061496, -0.3464251, -0.05068946, 0.1735782, 0.3337669, 
    0.4230736, 0.4649844, 0.4631779, 0.4851835, 0.3899689,
  0.1338983, -0.006629944, -0.1095591, -0.293478, 0.2386172, 0.1483502, 
    -0.09258401, 0.07152736, -0.07168564, -0.04040302, -0.2130267, 
    -0.4293027, -0.4640032, 0.1160749, 0.6747508, 0.3816674, 0.3994412, 
    0.3087349, 0.1129827, -0.009592056, -0.0400281, -0.07822752, -0.1220107, 
    -0.1751513, -0.1280975, -0.09316921, -0.05451298, 0.02296066, 0.02063274, 
    -0.0052948, -0.04111814, -0.09881687, -0.2838597, -0.2790911, -0.1094785, 
    0.033409, -0.03615499, -0.1273007, 0.268386, 0.7409127, 0.6532497, 
    0.5358992, 0.5658321, 0.4813099, 0.3608184, 0.2712183, 0.08756018, 
    -0.2481339, -0.2689025, -0.04082584, 0.117377, 0.4952579, 0.8485943, 
    1.143875, 1.290505, 1.232644, 1.115229, 0.9858013, 0.7539979, 0.5499128, 
    0.4521263, 0.4088646, 0.3494245, 0.2383894, 0.1688092, 0.2279564, 
    0.216856, 0.1862247, 0.1515405, 0.1905868, 0.234386, 0.2051864, 
    0.1963005, 0.09019661, 0.07702923, 0.2308383, 0.2683861, -0.01600504, 
    -0.09030533, -0.2671283, 0.001426458, 0.1303327, 0.1311302, -0.06042254, 
    -0.3616107, -0.5283262, -0.4751686, 0.007806599, 0.08139074, 0.3090762, 
    0.3223412, 0.3275661, 0.3365664, 0.2485299, 0.2257113, 0.1339784,
  -0.09263229, -0.1446338, -0.154139, -0.3350477, -0.02757746, -0.1937884, 
    -0.4703833, -0.1765195, -0.1172585, -0.09946877, -0.3397684, -0.4356179, 
    -0.2032285, 0.2059348, 0.5209422, 0.3512321, 0.2613068, 0.05173635, 
    -0.07743025, -0.2392631, -0.3526249, -0.4366269, -0.3842168, -0.2994676, 
    -0.2277722, -0.2446985, -0.1964087, -0.2350311, -0.2278042, -0.2072005, 
    -0.256125, -0.2811255, -0.3198953, -0.3555723, -0.1724179, -0.01576111, 
    0.1196555, -0.01371002, 0.2814558, 0.6261344, 0.4300566, 0.3995719, 
    0.4232044, 0.1367788, -0.08244324, -0.03796101, -0.2367568, -0.4550188, 
    -0.1755593, 0.2391706, 0.4417911, 0.6373314, 0.740489, 0.9097598, 
    0.9110944, 0.7584903, 0.683002, 0.5738386, 0.3768171, 0.1729759, 
    0.1169212, 0.1138288, 0.1165957, 0.2054466, 0.1581647, 0.09758568, 
    0.0401473, 0.03217196, 0.0212183, 0.07608557, 0.03004074, 0.03420639, 
    0.02507591, 0.01047707, 0.03384876, 0.1240501, -0.05604431, 0.0362246, 
    -0.08954024, -0.251959, -0.07765886, -0.1082416, -0.04142841, -0.1990619, 
    -0.4828998, -0.2544654, -0.08638281, 0.05289125, 0.08340883, 0.1670353, 
    0.1673281, 0.2094996, 0.1971464, 0.1182404, 0.07587433, -0.02083826,
  -0.1864953, -0.1194878, -0.1405168, -0.3040423, -0.2252663, -0.4168353, 
    -0.525722, -0.4021705, -0.3726784, -0.1665912, -0.1576231, -0.2295792, 
    0.06322718, 0.3490996, 0.3685493, 0.10146, -0.02292156, -0.1396537, 
    -0.2219453, -0.4287002, -0.5311418, -0.4598203, -0.4095268, -0.3523171, 
    -0.3434949, -0.3169322, -0.1698949, -0.2281637, -0.231158, -0.2846899, 
    -0.2141819, -0.2081275, -0.1655169, -0.09767818, -0.1012591, -0.1675352, 
    0.01661193, -0.02679586, -0.0003802776, 0.1540632, 0.03326273, 
    -0.001242161, -0.1896868, -0.3925838, -0.1240616, 0.01797938, -0.1677957, 
    0.1153587, 0.4302512, 0.5695417, 0.6705996, 0.7532168, 0.7565046, 
    0.7368757, 0.6470319, 0.5346783, 0.4333112, 0.2830508, 0.1246523, 
    0.1174909, 0.1383893, 0.1911075, 0.1532171, 0.05787206, 0.005805016, 
    -0.01650953, -0.1111877, -0.1068416, -0.07557535, -0.03057146, 
    -0.1203175, -0.06419849, -0.1271381, -0.1756568, -0.02845645, -0.1294981, 
    -0.03836858, -0.02655214, 0.03630596, -0.03003517, -0.0303607, 
    -0.1062071, -0.03255796, -0.3080299, -0.5838926, -0.1192604, 0.05626035, 
    0.01573348, 0.1468043, 0.0783143, 0.098351, 0.07103968, -0.01035786, 
    -0.04339695, -0.1489792, -0.2147503,
  -0.05656481, -0.04443908, -0.07874942, -0.09357691, -0.01481718, 
    -0.2476621, -0.08228123, -0.0589087, -0.2487363, -0.1681046, 0.02558041, 
    0.1082144, 0.2167907, 0.250319, 0.1549911, 0.106782, 0.04336977, 
    -0.0836482, -0.244895, -0.3279841, -0.3977759, -0.3796444, -0.4035537, 
    -0.46135, -0.4041889, -0.3786352, -0.5027394, -0.3867397, -0.174078, 
    -0.5710669, -0.2440004, -0.07510352, 0.02642632, -0.1839411, -0.1527238, 
    -0.04938698, -0.0836482, -0.112636, -0.02611274, 0.005137444, -0.3165579, 
    -0.2053113, -0.4046116, -0.3633034, 0.3577741, 0.7756776, 0.8642356, 
    1.263275, 1.315066, 1.220958, 1.162901, 1.016042, 0.9364362, 0.8619733, 
    0.7460553, 0.6039492, 0.4403098, 0.352761, 0.2396101, 0.2534283, 
    0.181537, 0.1819766, 0.174099, 0.1694932, 0.1500597, 0.07335067, 
    0.03345776, 0.1058049, 0.03510189, 0.008392572, 0.0350852, -0.003195524, 
    -0.08449435, -0.1640029, -0.1711318, 0.03194399, 0.005625635, 0.05124737, 
    0.02115297, 0.01127341, -0.03346944, -0.01427997, -0.2200905, -0.3603249, 
    -0.4127337, -0.6706439, -0.2286516, 0.07880282, 0.05888081, 0.04994559, 
    0.08358812, -0.0166235, -0.01310778, -0.04183531, -0.1060441, -0.06514263,
  -0.08395743, -0.07604742, -0.06449151, 0.04439515, -0.03589455, -0.1508523, 
    0.001231104, 0.02748436, -0.03446226, -0.0720762, -0.02497339, 0.4119582, 
    0.4490032, 0.399652, 0.2714627, 0.4661727, 0.295372, 0.02852607, 
    -0.1827532, -0.2229388, -0.1558164, -0.1826068, -0.3404031, -0.6392474, 
    -0.8445532, -0.9000709, -0.6169329, -0.09443948, -0.1596413, -0.6671271, 
    -0.1444719, -0.1260312, -0.07500589, -0.6866422, -0.6803446, -0.1740618, 
    -0.08268817, 0.003135383, -0.02803323, -0.1389866, -0.1925011, 
    0.06947684, 0.05222392, 0.2770937, 0.7430605, 0.9850689, 1.103966, 
    1.076996, 0.9807559, 0.887543, 0.7753686, 0.658474, 0.5240339, 0.4355736, 
    0.3747337, 0.344444, 0.278526, 0.2653261, 0.2813093, 0.2992455, 
    0.2497175, 0.2492292, 0.2293398, 0.2583927, 0.1472924, 0.1693954, 
    0.2401474, 0.2281194, 0.1376569, 0.03646874, -0.05907154, -0.2084205, 
    -0.2991431, -0.4257381, -0.4487852, -0.07883078, 0.03139061, 0.07390362, 
    -0.008957699, -0.02328062, 0.02206443, 0.06280351, -0.1283424, 
    -0.3804746, -0.4651263, -1.082574, -0.6762265, -0.3234756, -0.3340716, 
    -0.1694229, -0.1828835, -0.1583064, -0.07621002, -0.1536839, -0.09751534, 
    -0.08455968,
  -0.07427311, -0.1197972, -0.09496033, -0.009983093, 0.04120506, 0.06649803, 
    0.08558983, 0.09099349, 0.2212994, 0.09480206, -0.07262945, 0.3884385, 
    0.5038848, 0.6790638, 0.5174422, 0.6683372, 0.6059023, 0.4904889, 
    0.49669, 0.3186791, -0.01908135, -0.4323952, -0.6728899, -0.8472064, 
    -0.869993, -0.6974992, -0.08740819, 0.03655011, -0.3541237, -0.7204812, 
    -0.1989317, -0.02080666, -0.0401426, -0.7586647, -0.9363339, -0.4322324, 
    -0.140403, -0.02272724, -0.1804259, -0.2128637, -0.03032804, 0.1701927, 
    0.06848371, 0.1187929, 0.0691022, -0.02691019, -0.1573951, -0.4273984, 
    -0.406793, -0.2943906, -0.2965716, -0.2252338, -0.1823138, -0.1323951, 
    -0.1571184, -0.1986876, -0.1950579, -0.2188859, -0.1807675, -0.158632, 
    -0.1226618, -0.07402897, -0.1245661, -0.2234595, -0.3456438, -0.2777078, 
    -0.272727, -0.235878, -0.2801979, -0.2833717, -0.2956111, -0.2812231, 
    -0.231272, -0.2495661, -0.2169656, -0.04784116, -0.1538145, -0.05490506, 
    -0.00127542, 0.01106182, -0.1896706, -0.2195534, -0.2590717, -0.3183489, 
    -0.4153216, -0.485862, -0.4176002, -0.5172911, -0.5355691, -0.4490943, 
    -0.4875872, -0.3700902, -0.3211811, -0.4607317, -0.1556046, -0.124615,
  0.01474035, -0.08970284, 0.04092854, 0.1236432, 0.1353945, 0.1685162, 
    0.02328512, -0.01012957, 0.02076226, -0.1035703, -0.03639913, 0.1421816, 
    0.4011662, 0.8688102, 0.6171656, 0.3976178, 0.6216412, 0.8619571, 
    0.9119896, 0.6231549, 0.2265403, -0.278082, -0.628033, -0.733681, 
    -0.5940814, -0.310569, -0.05477476, -0.013987, -0.2366107, -0.677252, 
    -0.6659563, -0.2140196, 0.08570376, -0.1538144, -0.4126687, -0.3686256, 
    -0.282981, -0.2420957, -0.209088, -0.1640195, -0.1127661, -0.1262266, 
    -0.2079812, -0.1609759, -0.241819, -0.3365619, -0.5152891, -0.8931699, 
    -1.107151, -1.082428, -1.133583, -1.240891, -1.283062, -1.334186, 
    -1.346279, -1.3308, -1.216282, -1.036594, -0.8433814, -0.8002827, 
    -0.7494361, -0.7517798, -0.7816629, -0.7426164, -0.6748269, -0.699892, 
    -0.6680722, -0.3562396, -0.4325577, -0.3098041, -0.1794003, -0.178082, 
    -0.1342018, 0.007611275, -0.1659725, -0.05884376, -0.3900123, 
    -0.07830989, 0.233767, -0.07240158, -0.2279027, -0.4468157, -0.41358, 
    -0.5225808, -0.3917865, -0.209446, -0.1447324, -0.1136289, -0.06711197, 
    -0.1067114, -0.2310117, -0.2309303, -0.28469, -0.4368547, -0.03888929, 
    0.0146426,
  0.2122501, 0.2003196, 0.1464134, 0.1324811, 0.1621361, 0.4874942, 
    0.6306908, 0.5717064, 0.224636, 0.06667709, 0.1527937, 0.3549094, 
    0.5110292, 1.011616, 1.465213, 1.005609, 0.7302839, 0.833295, 0.7623314, 
    0.2579206, 0.08964258, -0.2403542, -0.9455462, -0.9900286, -0.6099505, 
    -0.3944069, -0.3933978, -0.1037819, 0.233002, -0.1650938, -0.7163307, 
    -0.7167703, -0.3733783, 0.02395245, -0.01110613, -0.4314675, -0.5412494, 
    -0.4773332, -0.3656634, -0.2463275, -0.05630472, -0.04622985, -0.1534564, 
    0.08837302, 0.08998437, 0.1019147, 0.1932884, 0.03327864, -0.07912374, 
    -0.2084694, -0.3454486, -0.4050514, -0.4002825, -0.5044492, -0.5982969, 
    -0.556207, -0.4780332, -0.3849342, -0.3087786, -0.4406796, -0.5095761, 
    -0.5437722, -0.6935443, -0.8016986, -0.6174863, -0.4631731, -0.3919655, 
    -0.1963763, -0.1916888, -0.06987893, 0.02533592, 0.1112246, -0.1243222, 
    -0.2134172, -0.1931699, -0.4078346, -0.4460996, -0.4854387, -0.6392472, 
    -0.3103087, -0.1010799, -0.1490295, -0.4067279, -0.3766985, -0.4177141, 
    -0.4315814, -0.3340229, -0.202203, -0.116884, -0.04600191, -0.05036396, 
    -0.0980202, 0.1451601, 0.1573834, 0.2333602, 0.1875267,
  0.3100527, 0.2858014, 0.1194277, 0.01776755, -0.2487686, -0.1638894, 
    0.0181582, 0.2740014, 0.06957436, -0.1593158, -0.154791, 0.08952868, 
    0.2380475, 0.3572208, 1.192393, 1.24088, 0.9926699, 0.8972924, 0.980528, 
    0.5398053, 0.2290305, 0.1561138, -0.7559792, -1.240696, -0.8309629, 
    -0.2516822, -0.04426038, -0.04076093, 0.1397402, 0.1578066, -0.09491134, 
    -0.2306861, -0.2703021, -0.08569924, 0.1224713, -0.2168516, -0.4895077, 
    -0.5618223, -0.524778, -0.3284075, -0.02555928, 0.1989687, 0.06690492, 
    0.05341209, -0.01091087, -0.01584244, 0.1350201, 0.03199291, 0.1450137, 
    0.1915468, 0.1432395, 0.08277404, 0.1899194, 0.3515568, 0.3057234, 
    0.1732037, 0.0804956, 0.1189232, 0.2329206, 0.1314719, 0.08436918, 
    0.1986759, 0.01955795, -0.3884823, -0.4330951, -0.2538633, -0.2350157, 
    -0.3412656, -0.3697976, -0.1811257, 0.0554468, 0.3198673, 0.1571393, 
    0.05136156, -0.1158097, -0.3980201, -0.4891498, -0.8606016, -0.7354388, 
    -0.2391009, -0.07067645, -0.1989478, -0.1988666, -0.1821349, -0.2667537, 
    -0.1925349, -0.1805398, -0.1565158, -0.04974508, 0.0522244, 0.09805751, 
    0.01228261, 0.3393985, 0.4304955, 0.4548281, 0.3288352,
  0.1062604, -0.1446999, -0.3988665, -0.1995662, -0.1329973, -0.2190485, 
    -0.3633361, -0.08996248, -0.04121637, -0.1614957, -0.4120007, -0.1980039, 
    0.04708071, 0.1033795, 0.367735, 0.2023216, 0.7642357, 0.9329693, 
    0.8031842, 0.7676538, 0.5028912, 0.9108666, 0.5028099, -0.4856666, 
    -0.9472064, -0.5694069, 0.08163476, 0.1818464, 0.3852646, 0.6991477, 
    0.219347, 0.1834736, 0.4434023, 0.3436954, 0.1799421, -0.1114642, 
    -0.4775124, -0.6051328, -0.4534563, -0.2776425, -0.1330137, 0.259955, 
    0.2819602, 0.08604553, 0.06565171, 0.05347741, 0.1292422, 0.04939187, 
    0.1239036, 0.2671329, 0.2525496, 0.08635473, -0.04974556, -0.0655818, 
    -0.0770731, -0.2286677, -0.3800187, -0.3127825, -0.107867, -0.04038644, 
    -0.08472252, 0.03897524, 0.04350042, -0.2399147, -0.4412165, -0.4781145, 
    -0.4312398, -0.4701557, -0.4452207, -0.09474856, 0.2520123, 0.2324486, 
    0.1733828, 0.7711856, 0.4488876, -0.02590106, -0.2621315, -0.3639545, 
    -0.2319395, -0.08761983, -0.02448499, -0.008501887, 0.08316469, 
    -0.02272725, -0.09878516, -0.1236873, -0.1971412, -0.1448624, 
    -0.05918503, 0.0464468, 0.1284456, 0.06854916, 0.1532981, 0.1954369, 
    0.2157167, 0.2763451,
  0.3483829, 0.09421617, -0.5357155, -0.6300673, -0.354856, -0.2644914, 
    -0.1944392, 0.03417349, 0.0170517, 0.2311954, 0.3981714, -0.1715228, 
    -0.1044655, 0.2308536, 0.4953068, -0.01294529, -0.00461185, 0.508588, 
    0.3098086, 0.4392519, 0.5007103, 0.6173282, 0.5315859, 0.2170026, 
    -0.04097268, -0.1184466, -0.04622984, 0.01234763, 0.2038193, 0.531652, 
    0.3737741, 0.1295848, 0.3664837, 0.6099229, 0.4595649, 0.1407819, 
    -0.3624895, -0.7808653, -0.7030658, -0.3943418, -0.2291888, 0.09989646, 
    0.3178489, 0.1914004, 0.1725365, 0.1919212, 0.230984, 0.1790795, 
    0.2144147, 0.3296002, 0.2803328, 0.2542424, 0.2846947, 0.2481713, 
    0.283767, 0.1201601, -0.1959367, -0.1497614, -0.002268076, 0.03249764, 
    -0.03895378, -0.08019733, -0.03794479, -0.01317263, 0.005625725, 
    -0.3207905, -0.6409239, -0.4262429, -0.13067, -0.05742764, 0.07823324, 
    -0.09087491, 0.1568626, 0.6328878, 0.154763, -0.1489968, -0.3147357, 
    -0.4081276, -0.2116433, -0.06956968, 0.02245505, 0.08020243, 0.08391345, 
    0.03334379, -0.01836526, -0.1334367, -0.1469295, -0.1546934, -0.1889048, 
    -0.1609421, -0.1881394, -0.02243376, 0.2054791, 0.1698997, -0.03226495, 
    0.1777449,
  0.05697656, 0.2149355, -0.3223203, -0.6440651, -0.5396217, -0.6402402, 
    -0.6411026, -0.4005587, -0.3331752, 0.1254339, 0.5726342, 0.1599713, 
    0.3003033, 0.4741967, 0.7169701, 0.2583112, 0.1069604, 0.7388939, 
    0.16308, -0.1529191, 0.2948672, 0.3445907, 0.2714785, 0.1549258, 
    -0.0559628, 0.0150983, -0.03135353, -0.3025286, -0.08268797, 0.233686, 
    0.3802843, 0.2212515, 0.08070803, 0.3810492, 0.4337835, 0.2876573, 
    -0.02668214, -0.439752, -0.5974343, -0.5831114, -0.4602109, -0.1245827, 
    0.3448021, 0.3771588, 0.2375267, 0.2572532, 0.2739525, 0.2449487, 
    0.2488223, 0.2795677, 0.2977319, 0.3166122, 0.2884545, 0.1621523, 
    0.1066837, -0.04185152, -0.3376684, -0.3169327, -0.1254449, -0.0966363, 
    -0.1210833, -0.1182346, -0.1314831, -0.08608818, 0.05896282, -0.0346899, 
    -0.2894427, -0.05772072, 0.2389915, 0.0887962, 0.1513614, 0.5366806, 
    0.5309513, 0.4146264, 0.05294025, -0.06338477, -0.2525775, -0.3777891, 
    -0.2361224, -0.08413655, 0.09550193, 0.1977806, 0.2211204, 0.1887799, 
    0.01832098, -0.1694394, -0.2026099, -0.1808, -0.1517959, -0.2048879, 
    -0.3379769, -0.3333211, -0.045578, 0.08663154, -0.3019589, -0.3437395,
  0.01789784, 0.2379987, 0.1164818, -0.3287331, -0.5297911, -0.5219948, 
    -0.4782773, -0.2834368, -0.3471079, 0.05061293, 0.2068789, 0.07414782, 
    0.3209741, 0.4045352, 0.2820255, 0.140733, 0.1792748, 0.6997501, 
    0.4364851, 0.1991479, 0.4095318, 0.2065371, 0.06918359, 0.09883848, 
    -0.3024955, -0.3005915, -0.05130792, -0.319504, -0.1417212, -0.02365494, 
    0.04328918, 0.2587347, 0.1446729, 0.1943474, 0.2898388, 0.2367296, 
    0.1444442, -0.06302643, -0.3757381, -0.6659564, -0.8018777, -0.5317603, 
    0.107123, 0.2737897, 0.1895775, 0.1783145, 0.1378847, 0.1886172, 
    0.293386, 0.3364362, 0.3840924, 0.4750267, 0.6164654, 0.5618756, 
    0.3555931, 0.155593, -0.1526101, -0.2689512, -0.1399148, -0.07760978, 
    -0.05485582, -0.02230358, -0.1137576, -0.2604384, -0.2415748, 0.1212509, 
    0.1939557, 0.1715761, 0.2368105, 0.4497988, 0.7571394, 1.159678, 1.00408, 
    0.4616152, 0.1283307, 0.02766335, -0.2580788, -0.3931862, -0.4081277, 
    -0.4035377, -0.2186419, -0.04837823, 0.005479246, 0.03407617, 
    -0.01776303, -0.2078346, -0.3791237, -0.3301491, -0.2094786, -0.2530818, 
    -0.266835, -0.4152236, -0.2063527, 0.04333758, 0.04794332, -0.03382754,
  0.3850364, 0.605463, 0.7813418, 0.492963, -0.343121, -0.8283262, 
    -0.7920631, -0.6041887, -0.4943733, -0.1015029, -0.02070892, -0.3224016, 
    -0.05894136, 0.187901, 0.06028059, 0.02318764, -0.05985296, 0.1940696, 
    0.4224225, 0.3931582, 0.2663515, 0.08295304, -0.4201717, -0.4473202, 
    -0.4414444, -0.5625215, -0.4792049, -0.3543839, 0.3204206, 0.3078555, 
    -0.1048398, 0.00281024, 0.07449007, 0.2220163, 0.3290634, 0.216043, 
    0.203738, 0.1359482, -0.05124283, -0.3360246, -0.7988665, -0.8092019, 
    -0.4164772, -0.3076555, -0.2378802, -0.02873302, 0.02295959, 0.06361723, 
    0.1613874, 0.3254986, 0.3756614, 0.3712018, 0.5209903, 0.5269636, 
    0.3856224, 0.149099, -0.2151588, -0.3903704, -0.4141332, -0.3784889, 
    -0.203017, -0.02082276, -0.06535482, -0.2733774, -0.1740124, 0.1645775, 
    0.4432071, 0.2364363, 0.243028, 0.5718691, 0.6452415, 0.533181, 
    0.5243269, 0.3280705, 0.2288028, 0.3365338, 0.1828229, -0.03719664, 
    -0.1951393, -0.2858946, -0.2279518, -0.1447487, -0.1540585, -0.2233782, 
    -0.220237, -0.2986712, -0.465517, -0.4047258, -0.2299863, -0.1464413, 
    -0.01769781, -0.0921278, -0.2904029, -0.237294, -0.1409401, 0.1192324,
  -0.03366474, -0.0115456, 0.1580019, 0.3767357, -0.01362893, -0.5250872, 
    -0.8703346, -0.8599989, -0.3642147, -0.09460205, -0.1173886, -0.1132221, 
    0.0288353, 0.1130801, -0.1463438, -0.1359758, -0.1217831, -0.175136, 
    0.06807685, 0.1423771, 0.09499738, 0.2935163, 0.3206646, 0.2049583, 
    0.3297304, 0.3796166, 0.2223575, 0.1802675, 0.5021752, 0.4032168, 
    -0.05734634, -0.2083879, -0.2061579, -0.07080674, -0.04888296, 
    -0.1130104, -0.06390572, -0.0339576, -0.003065586, -0.007687807, 
    -0.3296933, -0.5088437, -0.3641497, -0.3274308, -0.3329324, -0.3284237, 
    -0.2798073, -0.2148333, -0.1925026, -0.07524991, 0.05175209, 0.1570254, 
    0.2245058, 0.1994082, 0.2566673, 0.1508242, -0.1939186, -0.3759824, 
    -0.4625709, -0.5473855, -0.4073301, -0.1326718, -0.09932137, -0.2331758, 
    -0.04780841, 0.2835391, 0.4404889, 0.4223901, 0.536534, 0.7769961, 
    0.7926699, 0.556407, 0.440554, 0.2925559, 0.09542055, 0.0581159, 
    0.1556582, 0.2834902, 0.2549909, 0.07315505, 0.03672922, 0.06861401, 
    -0.1114968, -0.3908262, -0.4847878, -0.373492, -0.4190487, -0.4748594, 
    -0.4065651, -0.2286191, 0.04942441, 0.1672142, 0.1221623, 0.01047587, 
    -0.2074928, -0.2095599,
  0.0616966, 0.1580021, 0.03648496, -0.08965424, -0.282851, -0.5675839, 
    -0.8771542, -1.231598, -0.7905169, -0.412864, -0.4408098, -0.3558002, 
    -0.2721251, -0.2765033, -0.3226621, -0.2564349, -0.2954323, -0.5546283, 
    -0.01463804, 0.4600853, 0.223204, 0.09641337, 0.3848411, 0.3918724, 
    0.4783959, 0.6270449, 0.6436302, 0.128054, -0.03055602, 0.08239972, 
    0.03983787, -0.2254941, -0.4985737, -0.3830463, -0.1998594, -0.4428277, 
    -0.4619688, -0.2562884, -0.2068092, -0.06865788, -0.09123302, -0.185211, 
    -0.202903, -0.03682229, 0.1653914, 0.1383731, 0.07265031, 0.1233015, 
    0.1107688, 0.03697336, -0.006483674, 0.030056, 0.08489001, 0.07997465, 
    0.1210554, -0.01807225, -0.3607643, -0.5376199, -0.6135638, -0.6157448, 
    -0.4649798, -0.1633523, 0.07086027, 0.00058043, -0.03757098, 0.03646873, 
    0.2959251, 0.4643822, 0.4434187, 0.4232038, 0.6303327, 0.7258893, 
    0.6248964, 0.4627057, 0.2763777, 0.09405339, 0.05621156, 0.1305117, 
    0.2224713, 0.2707461, 0.4283796, 0.6093529, 0.4908144, 0.04543686, 
    -0.3054583, -0.3635474, -0.3941466, -0.4425677, -0.4328997, -0.2896706, 
    0.01475647, 0.2277936, 0.3379987, 0.380528, 0.06635171, -0.07987242,
  0.34975, 0.7373639, 0.4901634, -0.0647357, -0.3962624, -0.3699929, 
    -0.5032611, -0.9398984, -1.055198, -0.7420794, -0.3176003, -0.1387266, 
    -0.08044201, -0.08625257, -0.1541075, -0.1514219, -0.1923887, -0.4176167, 
    -0.1947813, 0.2331647, 0.1168399, -0.1009011, -0.01138285, -0.1600808, 
    -0.3877663, -0.1687233, 0.1503034, 0.08567122, -0.05301678, -0.02640557, 
    0.09984761, -0.1030658, -0.4161028, -0.4341367, -0.3227598, -0.4219785, 
    -0.5978249, -0.5022844, -0.4682675, -0.6388241, -0.5331113, -0.3164772, 
    -0.2027565, -0.04292572, 0.198985, 0.3670188, 0.425808, 0.4662539, 
    0.4910424, 0.4834576, 0.3277123, 0.1682396, 0.1125267, 0.02494526, 
    -0.08552027, -0.217454, -0.4192767, -0.7087297, -0.8836155, -0.8700902, 
    -0.7071021, -0.2838438, 0.2168888, 0.2934186, 0.1478945, 0.0334903, 
    0.2134056, 0.424278, 0.4329694, 0.2860944, 0.3572695, 0.4751407, 
    0.5317161, 0.4647403, 0.3465111, 0.1991804, 0.02678454, -0.05404234, 
    -0.09622985, -0.1034401, -0.01107341, 0.2706647, 0.5094993, 0.4269636, 
    0.1800072, -0.01427984, -0.1274636, -0.2285051, -0.3819232, -0.4476783, 
    -0.1578834, 0.1956323, 0.4719179, 0.6061465, 0.376866, 0.1846623,
  0.2622337, 0.3216901, 0.3090599, 0.1110455, -0.1624896, -0.2296933, 
    -0.3177468, -0.4505756, -0.7129615, -0.8294655, -0.6127011, -0.3036028, 
    -0.1124245, -0.02485937, -0.161155, -0.2780169, -0.2507546, -0.2116269, 
    -0.2419167, -0.1362038, 0.08160222, 0.2498313, 0.3808049, 0.2379498, 
    -0.008420594, 0.07922587, 0.2194277, 0.2399519, 0.184597, 0.125987, 
    0.1375104, 0.181765, 0.05928776, -0.158388, -0.3063535, -0.3774961, 
    -0.3795632, -0.5472226, -0.7837461, -1.080019, -1.179758, -1.014394, 
    -0.7332088, -0.4490292, -0.1329648, 0.208344, 0.5232201, 0.7357855, 
    0.8455997, 0.8696393, 0.7383244, 0.5389428, 0.3723252, 0.1566024, 
    -0.02178335, -0.1054094, -0.3366268, -0.6699605, -0.8445532, -0.8824763, 
    -0.8984916, -0.6250701, -0.03475475, 0.3262639, 0.3225691, 0.1914659, 
    0.1888616, 0.24975, 0.4300397, 0.5649518, 0.4638776, 0.3190045, 
    0.2745709, 0.3309023, 0.2487409, 0.1546652, 0.07784247, 0.04966867, 
    -0.0133847, -0.2207904, -0.4368712, -0.3593158, -0.2286024, -0.1608784, 
    -0.07070887, 0.07017636, 0.06854892, -0.08508062, -0.3521545, -0.5252664, 
    -0.3810933, -0.03892183, 0.2600366, 0.5556744, 0.6725206, 0.4189236,
  0.3688745, 0.2106552, 0.2471786, 0.3552188, 0.4260684, 0.2025495, 
    -0.1194232, -0.3286518, -0.4500547, -0.6152239, -0.5840878, -0.4556537, 
    -0.4207253, -0.3289121, -0.2190163, -0.2658751, -0.3222226, -0.2034401, 
    -0.03084886, -0.04165626, -0.1035378, 0.0547471, 0.2608342, 0.3064559, 
    0.4205019, 0.3734317, 0.4202904, 0.3901797, 0.4070254, 0.3717389, 
    0.3376732, 0.3956485, 0.3688905, 0.1620548, -0.05747658, -0.2054421, 
    -0.2736386, -0.3126199, -0.5129615, -0.8101785, -1.067258, -1.138108, 
    -1.099583, -0.9857317, -0.7286681, -0.2766008, 0.2007265, 0.6464136, 
    1.016824, 1.273464, 1.318565, 1.211599, 1.030544, 0.7384219, 0.4180768, 
    0.116189, -0.1965387, -0.4664447, -0.6072805, -0.705328, -0.8110232, 
    -0.6281457, -0.1175838, 0.1129012, 0.2450466, 0.1629987, 0.2358179, 
    0.2594668, 0.3153262, 0.4450951, 0.464903, 0.3462181, 0.2879337, 
    0.2983015, 0.3060651, 0.307058, 0.2081321, 0.1328717, 0.0265404, 
    -0.1148168, -0.2859107, -0.3321183, -0.4942278, -0.658209, -0.64081, 
    -0.3763566, -0.03371358, -0.009706259, -0.2558978, -0.4683814, 
    -0.4320536, -0.2048237, 0.1159775, 0.5283146, 0.7406197, 0.6353457,
  0.4505312, 0.2967389, -0.01486564, -0.1861384, -0.1037169, 0.0244571, 
    0.0385685, -0.1285865, -0.3259987, -0.4693906, -0.4315976, -0.3655658, 
    -0.474957, -0.5506079, -0.4322813, -0.3386127, -0.3591529, -0.3253152, 
    -0.1221085, 0.03249741, 0.04608786, 0.07764745, 0.2047138, 0.2700791, 
    0.2224228, 0.2451115, 0.2524194, 0.2402285, 0.2910913, 0.3734967, 
    0.3980898, 0.3960391, 0.4602318, 0.4768984, 0.3591574, 0.1751895, 
    0.063959, 0.04450917, -0.1687882, -0.5669003, -0.751487, -0.5966042, 
    -0.4167865, -0.659153, -0.7665424, -0.6102598, -0.266819, 0.1418073, 
    0.6463482, 1.075808, 1.282579, 1.303998, 1.300922, 1.145388, 0.7636663, 
    0.222211, -0.2109108, -0.4339576, -0.56091, -0.6727586, -0.7337451, 
    -0.4759326, -0.1406627, 0.08472776, -0.01644421, -0.05083585, 0.1218691, 
    0.2146426, 0.225629, 0.2566185, 0.3554792, 0.4977643, 0.6122009, 
    0.6104594, 0.5807883, 0.5891544, 0.4472597, 0.32322, 0.2626407, 
    0.1681907, -0.01966734, -0.2615619, -0.5216367, -0.795595, -0.8553118, 
    -0.615338, -0.1609759, 0.09670639, 0.1188254, -0.01761651, -0.04543233, 
    0.04016376, 0.1831975, 0.3162217, 0.4174912, 0.4603946,
  0.3322697, 0.4480085, 0.338552, 0.05461669, -0.198427, -0.2783751, 
    -0.2344949, -0.1438372, -0.1581764, -0.2548236, -0.3035377, -0.3467506, 
    -0.4301165, -0.5303605, -0.4848366, -0.3593482, -0.3091367, -0.3244687, 
    -0.2579812, -0.08818936, 0.100987, 0.3052027, 0.4480901, 0.470958, 
    0.4458277, 0.4593854, 0.4169869, 0.3416444, 0.3784122, 0.4574159, 
    0.4520287, 0.4092389, 0.467312, 0.5617292, 0.511713, 0.3592227, 
    0.3529401, 0.3042583, 0.03362131, -0.3473034, -0.3835506, -0.07612896, 
    0.1592389, 0.01714945, -0.2282445, -0.256516, -0.1304581, 0.1040633, 
    0.4731225, 0.9048933, 1.197634, 1.28393, 1.321479, 1.211094, 0.8290795, 
    0.3299583, -0.1289935, -0.3570696, -0.4102108, -0.4657607, -0.5113499, 
    -0.4324112, -0.120285, -0.1978571, -0.1424048, -0.02915633, 0.08360422, 
    0.1091738, 0.1384056, 0.199457, 0.2997338, 0.5052187, 0.5987734, 
    0.7392356, 0.8971948, 0.9850202, 0.9335878, 0.6293561, 0.4465438, 
    0.3741803, 0.1595809, -0.08275324, -0.3379126, -0.6303607, -0.8082416, 
    -0.7835345, -0.5939837, -0.3744525, -0.1624408, 0.0066185, 0.1538842, 
    0.3070905, 0.4111757, 0.3854108, 0.2729435, 0.2338812,
  0.3244896, 0.2491484, 0.2587185, 0.1947861, 0.02413154, -0.1308165, 
    -0.1212136, -0.04592049, 0.01613998, 0.01128972, -0.04227471, -0.1265032, 
    -0.1922909, -0.2563535, -0.3183327, -0.4145566, -0.436806, -0.4159075, 
    -0.3179095, -0.1950254, -0.02808201, 0.1540956, 0.2961856, 0.4171166, 
    0.4317813, 0.4565372, 0.4424584, 0.444086, 0.4891218, 0.5248965, 
    0.5103945, 0.3655541, 0.2288678, 0.1719179, 0.1396426, 0.04883853, 
    -0.02637303, -0.1776752, -0.4567277, -0.6373594, -0.5128636, -0.2523167, 
    -0.07498932, -0.2261612, -0.4198949, -0.4221895, -0.2820358, 0.04826927, 
    0.3980098, 0.823318, 1.11116, 1.129356, 0.9375429, 0.7282006, 0.609711, 
    0.3911563, 0.1863548, -0.02300376, -0.01248956, -0.09670138, -0.1067603, 
    -0.2089903, -0.3578994, -0.3409563, -0.2156634, -0.06001562, -0.03950787, 
    -0.04084241, 0.03728247, 0.1905867, 0.3548281, 0.4346133, 0.4444929, 
    0.5559838, 0.7762963, 1.01002, 1.082514, 0.901052, 0.7194766, 0.6096784, 
    0.49114, 0.3358828, 0.1337184, -0.08226466, -0.3340716, -0.5065488, 
    -0.6272032, -0.5842996, -0.4025612, -0.1432838, 0.1214622, 0.3782818, 
    0.591368, 0.7082785, 0.6877221, 0.5161889,
  0.5720644, 0.5252218, 0.4920192, 0.4541607, 0.3890243, 0.2600691, 
    0.1539817, 0.2061791, 0.2160261, 0.1723738, 0.08111393, 0.01718163, 
    -0.02555919, -0.1011451, -0.2035052, -0.3394427, -0.4335996, -0.4559141, 
    -0.4148984, -0.2467507, -0.08156508, 0.04437888, 0.1486269, 0.2280215, 
    0.2220156, 0.2327904, 0.2515403, 0.3047467, 0.539903, 0.8085554, 
    0.8940697, 0.8173608, 0.600808, 0.3154075, 0.1526634, 0.09481834, 
    -0.01745379, -0.2118223, -0.4110411, -0.5963275, -0.746246, -0.5316463, 
    -0.3600643, -0.3087461, -0.3899636, -0.5459855, -0.5573137, -0.2953172, 
    0.1866646, 0.8856716, 1.321821, 1.434468, 1.030073, 0.578998, 0.3084089, 
    0.2928327, 0.324457, 0.2804303, 0.2652774, 0.1977805, 0.1560488, 
    0.166905, 0.13961, 0.1298932, 0.09787828, 0.06812567, 0.0945254, 
    0.07035547, 0.04716212, 0.1030214, 0.2214296, 0.3399192, 0.3879825, 
    0.3813583, 0.3631778, 0.5400007, 0.666498, 0.6396751, 0.5396101, 
    0.5762311, 0.689903, 0.5901146, 0.3229921, 0.09856183, 0.01620507, 
    -0.1356828, -0.2619197, -0.4307175, -0.2443247, 0.1398709, 0.5545353, 
    0.787071, 0.9223087, 0.9312441, 0.8176212, 0.6816835,
  0.5680609, 0.4342064, 0.4027936, 0.4200786, 0.4186954, 0.4491155, 
    0.4692161, 0.4417261, 0.4106387, 0.3221784, 0.196739, -0.02982354, 
    -0.175836, -0.2669817, -0.2497294, -0.3395891, -0.3937396, -0.4379452, 
    -0.438287, -0.3550352, -0.250185, -0.09500909, 0.02977931, 0.06054115, 
    0.05901122, -0.009917974, -0.01686788, 0.01270586, 0.1610944, 0.3669049, 
    0.5525007, 0.6451601, 0.6313906, 0.5440859, 0.3984641, 0.3318463, 
    0.2032982, -0.06917904, -0.2559792, -0.4495177, -0.4940815, -0.2965553, 
    -0.0220924, 0.1332461, 0.1315696, -0.1767961, -0.3626848, -0.4086645, 
    0.06561995, -0.1863666, 0.8579698, 1.364871, 1.159939, 0.7995546, 
    0.4467227, 0.4016218, 0.4309675, 0.5100853, 0.5761661, 0.5928653, 
    0.5469016, 0.475987, 0.3521263, 0.2897239, 0.1666282, 0.08692446, 
    0.0529238, 0.06267317, 0.1183372, 0.1641868, 0.3530866, 0.3828718, 
    0.3229596, 0.2898217, 0.1512474, 0.07095778, 0.3084253, 0.452273, 
    0.5475041, 0.6458601, 0.5816835, 0.3909284, 0.1860619, 0.06265688, 
    -0.03623638, -0.1640846, -0.3150771, -0.5043831, -0.2189984, 0.01249504, 
    0.743453, 1.233817, 1.458784, 1.402061, 1.1546, 0.8437929,
  0.7217552, 0.3776634, 0.1210881, -0.0310604, -0.05324459, 0.02987731, 
    0.198204, 0.3858993, 0.5218694, 0.5576605, 0.4757754, 0.285948, 
    0.06161523, -0.1312396, -0.2740291, -0.2973365, -0.2194882, -0.1721087, 
    -0.1024798, -0.1706276, -0.1126687, -0.1122617, -0.1321511, -0.1543678, 
    -0.1370502, -0.1373105, -0.1381569, -0.1142962, -0.04066344, 0.09473696, 
    0.1966575, 0.2529726, 0.2532168, 0.2712182, 0.2591739, 0.3414329, 
    0.2444114, 0.04047264, -0.2364479, -0.4067768, -0.5018613, -0.4260801, 
    -0.2748268, -0.2022682, -0.1571673, -0.1971087, -0.3170954, -0.3938372, 
    -0.3777235, -0.3394752, -0.2397521, 0.00479579, 0.206342, 0.2470319, 
    0.2094668, 0.2145774, 0.2711368, 0.3610293, 0.4406028, 0.5334089, 
    0.6063256, 0.6084415, 0.5170839, 0.3281191, 0.2221295, 0.2079857, 
    0.2486269, 0.3839135, 0.4777611, 0.599929, 0.4985619, 0.36697, 0.2221133, 
    0.05456769, 0.02396876, 0.05987382, 0.2622501, 0.2663516, 0.5499616, 
    0.6611595, 0.5791119, 0.2861595, 0.09599042, 0.07429433, 0.0172956, 
    -0.0961647, -0.1894264, -0.211936, -0.2312226, -0.0731988, 0.1640244, 
    -0.1540084, 0.4335561, 1.151264, 1.336762, 1.086615,
  0.8935164, 0.7680442, 0.5792584, 0.3914491, 0.2389752, 0.1592552, 
    0.1825299, 0.280886, 0.3532493, 0.434369, 0.4148052, 0.267621, 0.132009, 
    0.0379173, 0.01138735, -0.1109434, -0.1647845, -0.1296771, -0.0565652, 
    0.04652733, 0.1700787, 0.2018496, 0.1399355, 0.02798897, -0.06525636, 
    -0.2119524, -0.2164609, -0.1859597, -0.1593158, -0.1259336, -0.1099505, 
    -0.1690651, -0.1428281, -0.1074929, -0.05568624, -0.03361592, 
    -0.05759053, -0.07970965, -0.1000873, -0.1588926, -0.2359434, -0.2796446, 
    -0.2779844, -0.2594459, -0.2444394, -0.2408586, -0.2315325, -0.230865, 
    -0.2073789, -0.1857969, -0.1520892, -0.1152401, -0.09341407, -0.08739197, 
    -0.09609962, -0.064345, -0.007313848, 0.05494201, 0.118207, 0.1780866, 
    0.2403425, 0.3210228, 0.3840111, 0.4242943, 0.4761172, 0.4696718, 
    0.4699323, 0.5256127, 0.5508894, 0.5349551, 0.4984479, 0.3015567, 
    0.1301212, 0.03238344, 0.0107038, -0.09875262, -0.1073301, 0.1471133, 
    0.1521588, 0.1465275, 0.1111758, 0.1351831, 0.2406032, 0.3488064, 
    0.3179467, 0.1935488, 0.1060488, 0.03650129, -0.09959912, -0.06777859, 
    -0.1225324, 0.04807425, -0.2245493, -0.007183075, 0.1377223, 0.5701931,
  0.2913352, 0.3678977, 0.4459577, 0.4195743, 0.3646914, 0.3606549, 
    0.3801211, 0.4226829, 0.4015241, 0.3478294, 0.2898704, 0.2366803, 
    0.1447044, 0.05725323, -0.04346291, -0.1289284, -0.1510801, -0.153196, 
    -0.1576882, -0.1433164, -0.1680235, -0.2053119, -0.251308, -0.3002012, 
    -0.3440489, -0.4522682, -0.4515685, -0.448541, -0.4313698, -0.4424701, 
    -0.4321348, -0.4194395, -0.4048236, -0.370416, -0.3358946, -0.2785704, 
    -0.2312071, -0.1958229, -0.1552142, -0.130084, -0.1105039, -0.09712501, 
    -0.06838152, -0.04110295, -0.01764905, -0.008306623, -0.006744087, 
    -0.01919526, -0.024306, -0.0333392, -0.03244382, -0.01818621, 
    0.004535198, 0.02986068, 0.05559307, 0.09299546, 0.1273053, 0.1618106, 
    0.211713, 0.2790794, 0.3501895, 0.4200137, 0.4662702, 0.4857038, 
    0.4914167, 0.4770938, 0.4426374, 0.4265241, 0.3923282, 0.3342878, 
    0.2618594, 0.3148216, 0.2290469, 0.166677, 0.1256614, 0.05767643, 
    0.01085031, -0.02552676, -0.08875895, -0.09800363, -0.0463438, 
    -0.01937437, 0.08786869, 0.1197209, 0.1455833, 0.1694766, 0.1859642, 
    0.1499453, 0.1062768, 0.00503993, -0.04133058, -0.02474523, -0.07020402, 
    0.04864359, 0.1529727, 0.2307236,
  -0.05547464, -0.05267513, -0.05835545, -0.04260021, -0.01818633, 
    -0.02666605, -0.02860287, -0.03595969, -0.03154886, -0.02941674, 
    -0.03947532, -0.05762312, -0.08195576, -0.1033262, -0.1243386, 
    -0.1451068, -0.1715554, -0.2046445, -0.2422096, -0.2974017, -0.3429095, 
    -0.3849505, -0.4308164, -0.4686582, -0.4997292, -0.5221087, -0.5544167, 
    -0.5779193, -0.5869688, -0.5790586, -0.5429258, -0.4964577, -0.4410866, 
    -0.3899473, -0.3372455, -0.2879453, -0.2390196, -0.1988666, -0.1695046, 
    -0.1400775, -0.1094623, -0.0796771, -0.04865497, -0.0174538, 0.00367251, 
    0.009304017, 0.008408815, 0.001621723, -0.001177847, -0.002024055, 
    -0.003407598, 0.001670599, 0.0118106, 0.03466225, 0.07318765, 0.131179, 
    0.1864362, 0.2639264, 0.3490013, 0.4223737, 0.4833438, 0.5470644, 
    0.5932233, 0.618793, 0.6354923, 0.6317325, 0.6147403, 0.5837018, 
    0.5494408, 0.5082461, 0.4603945, 0.4124128, 0.3598736, 0.2989526, 
    0.197211, 0.1950136, 0.1942812, 0.1901472, 0.2228945, 0.2434187, 
    0.2358502, 0.1892031, 0.1602806, 0.1339297, 0.1182396, 0.07671937, 
    0.03340883, -0.02373633, -0.07855403, -0.04123306, -0.05259371, 
    -0.0601784, -0.0490129, -0.04981053, -0.04243755, -0.04502535,
  -0.1108457, -0.1382709, -0.1548561, -0.1735899, -0.1915912, -0.210862, 
    -0.2298399, -0.2388731, -0.2533262, -0.2678119, -0.2858295, -0.3127663, 
    -0.3342995, -0.359153, -0.3895241, -0.4176654, -0.4479551, -0.4784076, 
    -0.5141335, -0.5575091, -0.5860736, -0.6096575, -0.6360409, -0.6561745, 
    -0.6760475, -0.6823789, -0.6853899, -0.6867245, -0.6780983, -0.6584694, 
    -0.6404192, -0.6098691, -0.5714902, -0.5334369, -0.4896543, -0.4412168, 
    -0.3931211, -0.3360573, -0.2858457, -0.2398822, -0.1964089, -0.1528867, 
    -0.1071673, -0.06108987, -0.02009051, 0.01845115, 0.05865297, 0.09761782, 
    0.1320579, 0.1640566, 0.1967064, 0.2349225, 0.2698021, 0.2997664, 
    0.3358015, 0.370502, 0.407351, 0.4483829, 0.4833438, 0.5207461, 
    0.5672957, 0.6091738, 0.6410912, 0.6608991, 0.6797467, 0.6921166, 
    0.699392, 0.7028587, 0.6928978, 0.6815534, 0.666612, 0.6505802, 
    0.6287539, 0.6069766, 0.5839785, 0.5583437, 0.5289817, 0.4999453, 
    0.4701276, 0.4341901, 0.3978457, 0.360362, 0.3254661, 0.2913841, 
    0.255707, 0.2183535, 0.1834902, 0.1495384, 0.1204368, 0.0926536, 
    0.06571677, 0.0410423, 0.01036194, -0.02100199, -0.04854104, -0.08202085,
  -0.08417344, -0.09358096, -0.1011987, -0.1065047, -0.1083603, -0.1081161, 
    -0.1050725, -0.1006286, -0.09457397, -0.0869894, -0.07948589, 
    -0.07199907, -0.06368256, -0.05686307, -0.05079174, -0.04514384, 
    -0.04073322, -0.03811276, -0.03702217, -0.03873104, -0.04205135, 
    -0.04890355, -0.05842495, -0.06853271, -0.08070719, -0.09374428, 
    -0.1078558, -0.1198676, -0.1327088, -0.1423116, -0.151654, -0.1588635, 
    -0.163878, -0.166254, -0.16396, -0.1596127, -0.15237, -0.1408305, 
    -0.1272244, -0.1112413, -0.09314203, -0.07426167, -0.05492544, 
    -0.03790092, -0.02193403, -0.008100033, 0.003472805, 0.009429932, 
    0.01895189, 0.03014946, 0.02723575, 0.03858018, 0.04352808, 0.03187466, 
    0.03914928, 0.04067922, 0.04616427, 0.04543209, 0.05859923, 0.06125247, 
    0.04507411, 0.05645108, 0.05490482, 0.06286371, 0.07088792, 0.07987225, 
    0.08996344, 0.09852457, 0.1112525, 0.1220273, 0.1326392, 0.1408423, 
    0.1437393, 0.160634, 0.1503475, 0.1513891, 0.1506892, 0.1438534, 
    0.1453019, 0.1400611, 0.1314348, 0.122532, 0.1116758, 0.1009011, 
    0.0908588, 0.07884708, 0.06597286, 0.05234945, 0.03802645, 0.0224669, 
    0.006874084, -0.009857655, -0.02675223, -0.0439229, -0.05923867, 
    -0.07221079,
  -0.169492, -0.2232358, -0.2674911, -0.3001082, -0.3169861, -0.3224061, 
    -0.315733, -0.3041773, -0.2902451, -0.2733341, -0.2572371, -0.2406681, 
    -0.2233667, -0.2037216, -0.1820743, -0.1599388, -0.1376568, -0.1155377, 
    -0.09026098, -0.06417048, -0.03881241, -0.01587945, 0.005051613, 
    0.0193581, 0.02808189, 0.03254151, 0.0301652, 0.01709533, -0.004583836, 
    -0.03588319, -0.07365942, -0.1119733, -0.1430779, -0.1635032, -0.1707788, 
    -0.163569, -0.1385527, -0.09836674, -0.04968548, 0.007492542, 0.06805611, 
    0.1139054, 0.1629453, 0.2266011, 0.2427959, 0.2221742, 0.2510478, 
    0.2414451, 0.2266173, 0.1862686, 0.1811577, 0.1424534, 0.102854, 
    0.08831954, 0.06066686, 0.05267531, 0.02305283, -0.00227271, -0.01490295, 
    -0.03917062, -0.07230866, -0.1171818, -0.1595974, -0.1947536, -0.2280382, 
    -0.2512641, -0.2458601, -0.2080996, -0.128998, -0.03057674, 0.05925083, 
    0.1474178, 0.210797, 0.2558813, 0.2516983, 0.2263565, 0.1883194, 
    0.1493709, 0.088238, 0.03801024, 0.02290606, 0.02549398, 0.05933225, 
    0.08403915, 0.1356017, 0.1795957, 0.2139868, 0.2334858, 0.2363665, 
    0.220253, 0.1873596, 0.1403058, 0.08259034, 0.022434, -0.040277, -0.106276,
  -0.2164657, -0.2984641, -0.3518331, -0.3639097, -0.351264, -0.3322535, 
    -0.308832, -0.2933046, -0.2834413, -0.2635032, -0.2256942, -0.1794702, 
    -0.1236107, -0.05901146, -0.002598763, 0.03669167, 0.05080318, 
    0.04191649, 0.02085561, 0.0006569922, -0.02011125, -0.05049872, 
    -0.08248097, -0.1091248, -0.1187115, -0.1072043, -0.07898176, 
    -0.05232179, -0.0357039, -0.02982831, -0.03308368, -0.04551792, 
    -0.07243848, -0.1048448, -0.1347921, -0.1493425, -0.1515231, -0.1352806, 
    -0.1091576, -0.06677437, -0.003314018, 0.03791356, 0.1059794, 0.1425354, 
    0.1628149, 0.1808813, 0.1853409, 0.1912326, 0.195497, 0.1729875, 
    0.1325741, 0.08542258, 0.05415636, 0.04598577, 0.03815699, 0.03058869, 
    0.0333879, 0.02637315, 0.01735592, -0.01190829, -0.0617938, -0.1445088, 
    -0.2471945, -0.3334737, -0.3837829, -0.405496, -0.3817486, -0.3139263, 
    -0.1853457, -0.02907956, 0.1171441, 0.2161682, 0.2449279, 0.2333558, 
    0.1726944, 0.09704328, -0.01705122, -0.1603293, -0.1963811, -0.2131779, 
    -0.1733176, -0.0908308, 0.005539894, 0.09600204, 0.2186258, 0.3335997, 
    0.4076068, 0.4461972, 0.4515033, 0.4232805, 0.358876, 0.2627015, 
    0.1751361, 0.08776665, -0.009581089, -0.1143336,
  -0.01081753, -0.02979577, -0.03030026, -0.02299213, -0.02463597, 
    -0.03635472, -0.05059624, -0.04426515, -0.007448673, 0.05838776, 
    0.1326392, 0.1890516, 0.2316625, 0.2726457, 0.2990615, 0.2988663, 
    0.2517958, 0.1642797, 0.06089437, -0.02219458, -0.08822668, -0.1042426, 
    -0.07082725, -0.01809287, 0.01406837, 0.01790929, 0.01374292, 
    -0.002777398, -0.03187907, -0.05287492, -0.07374108, -0.09452558, 
    -0.1028427, -0.09141684, -0.0687443, -0.03619254, 0.01115489, 0.06642818, 
    0.1104066, 0.1571186, 0.2000554, 0.2308822, 0.2771714, 0.3149807, 
    0.3572977, 0.3855853, 0.3950255, 0.4004939, 0.4264215, 0.3997779, 
    0.3281797, 0.2384011, 0.1269754, 0.03854762, -0.02810276, -0.03949594, 
    -0.03186274, -0.0152775, -0.04898512, -0.106521, -0.09149837, 
    -0.08764058, -0.08386448, -0.06853247, -0.05173558, -0.01745844, 
    0.05853462, 0.1172907, 0.1688209, 0.2009501, 0.208307, 0.165159, 
    0.07183242, -0.0457294, -0.196902, -0.3324814, -0.4429306, -0.4852479, 
    -0.4434837, -0.3879335, -0.2670516, -0.07294345, 0.09258401, 0.2357807, 
    0.3395079, 0.4314187, 0.4813211, 0.483388, 0.425608, 0.3327206, 
    0.2182674, 0.1919981, 0.1105363, 0.09040284, 0.0625546, 0.02419186,
  0.02043247, 0.0481503, 0.09242117, 0.1327202, 0.1766497, 0.2263403, 
    0.2648499, 0.2567444, 0.2165916, 0.1377177, 0.07463169, 0.04554605, 
    0.08021402, 0.1462134, 0.1762917, 0.1114483, -0.01581383, -0.1201925, 
    -0.2521267, -0.2351828, -0.1636171, -0.05684662, 0.08452749, 0.2125542, 
    0.2660539, 0.2680887, 0.216542, 0.1229718, 0.01281548, -0.08062553, 
    -0.1439559, -0.1509058, -0.1053653, -0.03082108, 0.06478477, 0.1549051, 
    0.2396226, 0.3090718, 0.3702044, 0.408762, 0.4076719, 0.351666, 
    0.2755427, 0.1823459, 0.09043598, 0.1166892, 0.1585999, 0.2815323, 
    0.4019749, 0.4021868, 0.3112201, 0.1900125, 0.05788355, -0.03309952, 
    -0.08598039, -0.06631893, -0.02206437, -0.03708715, -0.0538352, 
    -0.04991267, -0.04304418, -0.01259172, 0.01898378, 0.03976828, 
    0.04575771, -0.005169988, -0.09110761, -0.2084415, -0.3523218, 
    -0.4242293, -0.4544865, -0.4643335, -0.5178002, -0.6011986, -0.6772078, 
    -0.710655, -0.7032657, -0.5715599, -0.4728295, -0.367377, -0.2024682, 
    -0.01493561, 0.168349, 0.337278, 0.4428445, 0.5216368, 0.5209044, 
    0.4549538, 0.3811908, 0.3029194, 0.2226296, 0.06966752, -0.006276488, 
    -0.0320904, -0.01358455, 0.005800217,
  -0.1276145, -0.1271424, -0.062787, -0.06999737, -0.0476017, -0.06929791, 
    -0.05681372, 0.03574777, -0.026443, -0.1017358, -0.131163, -0.1656191, 
    -0.1803, -0.1048118, -0.03285563, -0.01417041, -0.07833004, -0.1495376, 
    -0.223366, -0.2455997, -0.1290796, -0.03622448, 0.04240504, 0.08182561, 
    0.04074466, -0.03529668, -0.1138287, -0.1569114, -0.1702902, -0.1981871, 
    -0.2291286, -0.2290633, -0.185704, -0.1151469, -0.04166007, 0.04434204, 
    0.09457016, 0.09422803, 0.09613228, 0.0832417, 0.06442666, 0.01799107, 
    -0.07072949, -0.1545999, -0.1580341, -0.02458739, 0.1885312, 0.3772842, 
    0.4853085, 0.468821, 0.3186095, 0.1197651, 0.03143498, 0.008306742, 
    -0.0001080632, -0.03596401, -0.09190476, -0.1668722, -0.2277446, 
    -0.2335877, -0.2364849, -0.2470969, -0.316205, -0.4214459, -0.5495546, 
    -0.6628358, -0.74044, -0.7985618, -0.8511497, -0.8594667, -0.8167095, 
    -0.7228618, -0.6455345, -0.602468, -0.5901308, -0.6162701, -0.6468853, 
    -0.6259869, -0.5086855, -0.3655702, -0.1928977, -0.1105411, 0.002333522, 
    0.1587136, 0.3132546, 0.4107156, 0.4070209, 0.2806374, 0.1765359, 
    0.1026264, 0.05814396, -0.001393795, -0.03724992, -0.09979874, 
    -0.1511822, -0.1542909,
  -0.5458274, -0.4986106, -0.501817, -0.5490174, -0.6251406, -0.6675724, 
    -0.6530375, -0.5625591, -0.4436954, -0.3231388, -0.2594178, -0.251996, 
    -0.3132753, -0.3377057, -0.2929956, -0.2850366, -0.2585881, -0.3099554, 
    -0.4129825, -0.5317978, -0.5256124, -0.4226831, -0.3560816, -0.3391056, 
    -0.3814396, -0.4615666, -0.4988221, -0.4448671, -0.3880801, -0.3067489, 
    -0.2737895, -0.2614524, -0.2417908, -0.1665144, -0.2341902, -0.2241968, 
    -0.2641053, -0.20058, -0.1437116, -0.07453859, -0.08337641, -0.1790959, 
    -0.3167423, -0.3732202, -0.2551374, -0.06475645, 0.1216368, 0.2397195, 
    0.2290913, 0.1084859, -0.04805726, -0.1489524, -0.2109967, -0.2309023, 
    -0.233539, -0.3375755, -0.4886661, -0.5959088, -0.6172141, -0.5122011, 
    -0.4211043, -0.4560976, -0.5660585, -0.7168398, -0.7698183, -0.76072, 
    -0.7838808, -0.7853293, -0.7570417, -0.7208436, -0.6994406, -0.6456158, 
    -0.6396262, -0.6272076, -0.621983, -0.7387799, -0.8234804, -0.804535, 
    -0.6806418, -0.4693463, -0.335134, -0.3803488, -0.3222597, -0.184776, 
    -0.03744522, 0.01105738, -0.05420955, -0.1331321, -0.2083111, -0.23572, 
    -0.2882102, -0.3375754, -0.3666933, -0.4325299, -0.5087831, -0.5610129,
  -0.7924745, -0.8405864, -0.8638451, -0.9014101, -0.9393983, -0.9744406, 
    -0.8990827, -0.757416, -0.6236268, -0.4792258, -0.4164817, -0.4111431, 
    -0.4955507, -0.5928651, -0.6597272, -0.6504499, -0.5762799, -0.643858, 
    -0.8954367, -1.044167, -1.109581, -1.053477, -0.9934836, -0.9813254, 
    -0.9793886, -0.9626405, -0.879063, -0.7364198, -0.6088157, -0.4996848, 
    -0.5293723, -0.6412864, -0.7239036, -0.7290305, -0.7064719, -0.6488059, 
    -0.5645449, -0.4599712, -0.3373964, -0.2946067, -0.4034609, -0.6048117, 
    -0.8684348, -1.064626, -0.8886497, -0.6507916, -0.4629498, -0.4385682, 
    -0.4634055, -0.4734484, -0.4762965, -0.49962, -0.5542259, -0.6180447, 
    -0.7624294, -0.8085229, -0.9148059, -0.9179468, -0.8025011, -0.6140729, 
    -0.5934678, -0.6944278, -0.8960068, -0.9934676, -1.01767, -0.9758079, 
    -0.9947859, -1.021137, -1.03559, -1.017328, -1.026687, -1.05932, 
    -1.140277, -1.18157, -1.244704, -1.322716, -1.404568, -1.289838, -1.0553, 
    -0.846153, -0.7366152, -0.8314394, -0.741254, -0.5109479, -0.2772564, 
    -0.2351991, -0.2808371, -0.2565858, -0.2483339, -0.3186951, -0.442035, 
    -0.5411235, -0.577354, -0.5738385, -0.6285911, -0.6969992,
  -0.761664, -0.9403424, -1.018565, -1.082595, -1.063568, -1.004079, 
    -0.9752707, -0.9646266, -0.9493271, -0.9382919, -0.9600366, -1.028363, 
    -1.143093, -1.288129, -1.360232, -1.369704, -1.387022, -1.494476, 
    -1.650548, -1.730561, -1.730447, -1.662266, -1.587185, -1.408849, 
    -1.269786, -1.127729, -0.7934517, -0.5419705, -0.4090602, -0.4726344, 
    -0.539708, -0.6680772, -0.8045516, -0.8797147, -0.8928654, -0.8553169, 
    -0.7870878, -0.7605252, -0.9246036, -1.19791, -1.432497, -1.584727, 
    -1.687592, -1.659499, -1.464871, -1.238178, -1.067117, -1.017507, 
    -1.034874, -1.01225, -0.9875753, -1.059727, -1.170616, -1.216449, 
    -1.112836, -1.000939, -0.9489038, -0.8930445, -0.9113876, -0.9782821, 
    -0.9917589, -0.9885037, -1.090815, -1.234972, -1.292898, -1.310297, 
    -1.402338, -1.564008, -1.666157, -1.620274, -1.581716, -1.667638, 
    -1.813129, -1.920828, -1.978819, -2.037429, -1.948269, -1.678494, 
    -1.334581, -1.06404, -0.9415793, -0.8099713, -0.6284121, -0.4620383, 
    -0.4138287, -0.4250429, -0.4088157, -0.3783796, -0.3994408, -0.5091576, 
    -0.6060327, -0.6557235, -0.6932884, -0.6559024, -0.6616803, -0.6934512,
  -0.6635851, -0.8626249, -0.9682884, -0.9795024, -1.00836, -1.135606, 
    -1.229633, -1.218223, -1.202208, -1.227761, -1.254877, -1.298253, 
    -1.464561, -1.625694, -1.64879, -1.525336, -1.396593, -1.386908, 
    -1.510867, -1.620844, -1.589154, -1.467784, -1.267637, -1.092198, 
    -0.9523543, -0.7273871, -0.4549098, -0.2521918, -0.2331326, -0.3771749, 
    -0.530072, -0.6720479, -0.841742, -0.9882588, -1.06225, -1.119786, 
    -1.161241, -1.263731, -1.486876, -1.759727, -1.881, -1.874782, -1.826427, 
    -1.740651, -1.637103, -1.513991, -1.386533, -1.297292, -1.280885, 
    -1.276329, -1.349522, -1.474228, -1.494964, -1.300092, -1.080088, 
    -1.023675, -1.038552, -1.023871, -0.9780865, -0.9429301, -0.9386983, 
    -0.9486268, -1.09529, -1.334337, -1.512006, -1.644167, -1.793728, 
    -1.879942, -1.776215, -1.628949, -1.652989, -1.817995, -1.939073, 
    -1.988568, -1.981423, -1.858392, -1.569655, -1.247047, -1.006439, 
    -0.8218859, -0.724604, -0.5714626, -0.4209253, -0.3780869, -0.4619086, 
    -0.5448999, -0.5364691, -0.5202093, -0.5249945, -0.4989041, -0.3816026, 
    -0.3309513, -0.4447207, -0.5675076, -0.5724068, -0.5793566,
  -0.5769796, -0.7523701, -0.8871677, -0.9933853, -1.129388, -1.28598, 
    -1.344883, -1.260215, -1.215179, -1.307138, -1.39975, -1.408213, 
    -1.37322, -1.225775, -1.028575, -0.9242942, -0.9533956, -1.021885, 
    -1.073773, -1.035833, -0.8236425, -0.6044698, -0.5822041, -0.6080182, 
    -0.49018, -0.2768819, -0.1220481, -0.1300395, -0.3423111, -0.5551202, 
    -0.6040299, -0.6312273, -0.7617612, -0.912884, -1.049538, -1.182806, 
    -1.247829, -1.258294, -1.373724, -1.60429, -1.703314, -1.685004, 
    -1.610964, -1.549538, -1.476816, -1.402711, -1.252517, -1.149912, 
    -1.194248, -1.285459, -1.405576, -1.447633, -1.30831, -1.052159, 
    -0.8684022, -0.8247173, -0.799587, -0.6590271, -0.6199646, -0.7188091, 
    -0.8121033, -0.8602643, -1.079616, -1.355756, -1.502582, -1.565879, 
    -1.631781, -1.540424, -1.322064, -1.264333, -1.400564, -1.522568, 
    -1.520632, -1.483441, -1.417474, -1.177387, -0.7852974, -0.400645, 
    -0.22602, -0.230479, -0.2232528, -0.1442652, -0.05826259, -0.03565502, 
    -0.09122157, -0.2095158, -0.2940047, -0.3094507, -0.2698022, -0.1517519, 
    -0.01550531, -0.03362083, -0.2223089, -0.3497827, -0.3809509, -0.4172304,
  -0.6290624, -0.7066178, -0.7236423, -0.7796319, -0.8738544, -0.8814061, 
    -0.7865169, -0.6979589, -0.6798766, -0.6596782, -0.5438254, -0.4179301, 
    -0.3370056, -0.2919536, -0.2867615, -0.3890727, -0.5003357, -0.4422302, 
    -0.3539164, -0.2766864, -0.1878195, -0.1734803, -0.2809348, -0.2733011, 
    -0.1466575, -0.07278037, -0.1292744, -0.2695088, -0.3801696, -0.3542418, 
    -0.2783141, -0.3585229, -0.5548449, -0.7405534, -0.8553646, -0.9105077, 
    -0.9748468, -1.078363, -1.216058, -1.31334, -1.364187, -1.357432, 
    -1.34459, -1.203412, -0.9948175, -0.8398044, -0.715781, -0.6731222, 
    -0.7467711, -0.8077414, -0.7816672, -0.7741151, -0.6619406, -0.4770284, 
    -0.3986592, -0.4012959, -0.2966084, -0.2082133, -0.2726176, -0.4296327, 
    -0.4857197, -0.5802186, -0.8455505, -1.095274, -1.077484, -1.031016, 
    -0.9613547, -0.7900167, -0.6111269, -0.6870055, -0.8380637, -0.8706157, 
    -0.8344502, -0.7071555, -0.3964782, 0.02054644, 0.2863021, 0.3855529, 
    0.3418677, 0.3102762, 0.304986, 0.3696182, 0.3965714, 0.3394425, 
    0.3154514, 0.264931, 0.1252174, 0.04403257, 0.03831935, 0.04382086, 
    -0.003265858, -0.08948016, -0.2008083, -0.3114197, -0.4198506, -0.5211854,
  -0.04437852, -0.02357745, 0.008291006, -0.05473018, -0.1343203, 0.01698208, 
    0.2336318, 0.280328, 0.1992732, 0.1166236, 0.04551351, -0.03502035, 
    -0.1701927, -0.3303816, -0.4155543, -0.3814886, -0.2816186, -0.1358504, 
    -0.009222984, 0.01935792, -0.006195068, -0.05336308, -0.03389668, 
    0.02303672, -0.02168989, -0.07688236, -0.06128979, -0.008457184, 
    0.1323628, 0.2822819, 0.2806377, 0.193691, 0.07959604, -0.1073833, 
    -0.2761006, -0.327826, -0.3791442, -0.4708598, -0.4728787, -0.3931587, 
    -0.4885036, -0.667817, -0.6802843, -0.5310159, -0.3268168, -0.217751, 
    -0.1988871, -0.1992941, -0.3414333, -0.4019637, -0.4082627, -0.4211531, 
    -0.3045349, -0.226068, -0.2355087, -0.09577894, 0.09984279, 0.2098851, 
    0.1571183, 0.05610895, -0.124018, -0.3482692, -0.5243266, -0.4996684, 
    -0.2860453, -0.1652284, -0.06804395, 0.05682588, 0.08037734, -0.06273794, 
    -0.1687112, -0.09932709, 0.02069235, 0.2367244, 0.5937885, 1.097581, 
    1.375836, 1.149387, 0.6898173, 0.3636287, 0.2745503, 0.3823136, 
    0.5258361, 0.537913, 0.5769266, 0.5732645, 0.4005754, 0.2682512, 0.24107, 
    0.1974015, 0.1102271, -0.0001571178, -0.1162212, -0.1869407, -0.1802185, 
    -0.09257197,
  0.5262756, 0.5278869, 0.5206437, 0.4621477, 0.5536519, 0.7391496, 
    0.7178768, 0.4829484, 0.228912, -0.01579833, -0.2694441, -0.4482529, 
    -0.454031, -0.3570417, -0.2719669, -0.1217556, 0.04220939, 0.1312723, 
    0.202008, 0.2551005, 0.3102763, 0.3817277, 0.4350803, 0.4312885, 
    0.4008355, 0.5195534, 0.6315322, 0.692796, 0.8434789, 0.8935442, 
    0.7595274, 0.6245013, 0.4172423, 0.1734595, 0.06584227, 0.1122453, 
    0.2749569, 0.3788634, 0.3856829, 0.1719787, -0.1255147, -0.4028751, 
    -0.2377061, -0.1361597, -0.09426522, 0.06305909, 0.1874895, 0.1259007, 
    -0.006325722, -0.1987247, -0.2058702, -0.1165633, 0.04370689, 0.1288631, 
    0.1991916, 0.4036841, 0.5804259, 0.6144102, 0.4985087, 0.2730691, 
    0.058339, -0.05490959, -0.01024818, 0.1837945, 0.3752339, 0.4451065, 
    0.4477756, 0.4437718, 0.3928277, 0.3148167, 0.3142638, 0.3748921, 
    0.6030004, 0.9776101, 1.254124, 1.869619, 2.468837, 1.678993, 0.3741759, 
    -0.14822, 0.102952, 0.5168026, 0.9926002, 1.093463, 0.8742408, 0.6929746, 
    0.4386288, 0.3407773, 0.2814025, 0.1565814, 0.04946852, -0.07222748, 
    -0.08695674, 0.0927794, 0.3055725, 0.4901266,
  0.6659403, 0.7023332, 0.7885637, 0.9842833, 1.333827, 1.296083, 0.9527235, 
    0.6120659, 0.113987, -0.3390566, -0.3091903, -0.005576968, 0.1634337, 
    0.2574116, 0.264166, 0.3633194, 0.4528866, 0.4593804, 0.5047095, 0.59343, 
    0.6851618, 0.7712946, 0.8442113, 0.9033909, 0.9495499, 1.027577, 
    1.034902, 1.072011, 1.149469, 1.074762, 0.9301976, 0.6590387, 0.3252823, 
    0.296067, 0.4267474, 0.5349017, 0.6491433, 0.5664773, 0.2542051, 
    0.1058328, -0.07406631, -0.3789821, -0.3972275, -0.266482, -0.005625725, 
    0.2713114, 0.2693091, 0.1245174, -0.03100014, -0.03646898, 0.1459044, 
    0.2542865, 0.3794332, 0.5022033, 0.6665586, 0.8678121, 0.9305233, 
    0.8923887, 0.7269752, 0.4830299, 0.3416072, 0.2754616, 0.3900286, 
    0.6110574, 0.8141497, 0.7529031, 0.633665, 0.6180561, 0.5830139, 
    0.5477761, 0.7325577, 0.814752, 0.908258, 1.212962, 1.483632, 2.047305, 
    2.19343, 0.9083557, -0.3760357, -0.1661073, 0.7295633, 1.03067, 1.24374, 
    1.020416, 0.3928445, 0.1767474, 0.01276612, -0.06306362, -0.06802797, 
    -0.1507592, -0.09457445, -0.005381823, 0.1965876, 0.4516006, 0.639117, 
    0.7258196,
  0.5908425, 0.6944395, 0.8433487, 1.156956, 1.259299, 0.9184632, 0.4610732, 
    0.3166723, 0.004579514, -0.3382919, -0.06239665, 0.4157287, 0.3566791, 
    0.2349016, 0.3327045, 0.4495177, 0.49317, 0.5476297, 0.7103087, 
    0.8636451, 0.968642, 1.004791, 1.042828, 1.144342, 1.127545, 1.024046, 
    0.9559954, 0.9651747, 0.9040747, 0.8621488, 0.808176, 0.5966048, 
    0.3797094, 0.5213597, 0.5182674, 0.4641982, 0.5167534, 0.3386611, 
    0.1014055, 0.07674748, -0.1177351, -0.4900167, -0.3479114, 0.1339413, 
    0.4281471, 0.4527892, 0.2649799, 0.2477598, 0.3146707, 0.3347553, 
    0.4027728, 0.4540587, 0.5981505, 0.8277076, 0.8919005, 0.8866434, 
    0.889394, 0.8372293, 0.7398171, 0.5817442, 0.4752338, 0.4515685, 
    0.5222391, 0.76983, 0.9074278, 0.8281473, 0.7321672, 0.7818256, 
    0.7801003, 0.7454159, 0.8982317, 0.9640847, 0.9662979, 1.114507, 
    1.284772, 1.469684, 0.8166232, -0.1659117, -0.2448997, 0.5416563, 
    1.059967, 0.7784727, 0.7487202, 0.4209532, -0.2396753, -0.2670516, 
    -0.2564397, -0.2502387, -0.08952904, -0.009076357, 0.160862, 0.3422745, 
    0.5135313, 0.5860735, 0.6176163, 0.6606666,
  0.3070204, 0.4811754, 0.5962772, 0.7479882, 0.3953834, -0.03737998, 
    -0.4111757, -0.3562446, -0.1319767, -0.0754171, 0.1479226, 0.4594295, 
    0.07057869, -0.3321397, -0.08412504, 0.1820694, 0.2988827, 0.5559956, 
    0.6446023, 0.5493224, 0.68456, 0.7462624, 0.6759012, 0.679075, 0.5979389, 
    0.549973, 0.5214412, 0.4270086, 0.4027076, 0.6987362, 0.5769587, 
    0.2379622, 0.2794817, 0.4486061, 0.2604878, 0.3449928, 0.3540096, 
    0.06042242, -0.1271265, -0.3540956, -0.3275498, 0.1947811, 0.636806, 
    0.8545632, 0.7472227, 0.4624246, 0.347532, 0.4085508, 0.400722, 
    0.1992409, 0.1984271, 0.3564675, 0.5551164, 0.7343971, 0.7597064, 
    0.7719948, 0.8484759, 0.8264057, 0.6114479, 0.4370824, 0.5310931, 
    0.6523008, 0.7950417, 0.9298074, 0.9917701, 1.035195, 0.9927955, 
    0.9133521, 0.9122781, 0.9656147, 0.9965553, 0.9138888, 0.8385965, 
    0.8232162, 0.903863, 0.9178762, 0.08981657, -0.3738061, -0.1687766, 
    0.1852761, 0.4786676, 0.178082, 0.08438095, -0.00227271, -0.3339458, 
    -0.2434833, -0.1229436, -0.02369165, 0.06847882, 0.1876522, 0.3046443, 
    0.316591, 0.3616759, 0.2789447, 0.2727273, 0.296832,
  0.2957907, 0.3795304, 0.3354549, 0.3064365, 0.002382755, -0.2419862, 
    -0.2461204, -0.04918024, 0.1180398, 0.1753477, 0.1960832, 0.2581117, 
    0.01880455, -0.5056423, -0.1961851, 0.2293028, 0.2604226, 0.3040261, 
    0.2880757, 0.342112, 0.6028868, 0.6112199, 0.4324111, 0.3469945, 
    0.2832901, 0.2959044, 0.3655014, 0.3556376, 0.3434291, 0.4348855, 
    0.1911688, 0.198704, 0.3254129, 0.2195209, -0.03441787, 0.04347897, 
    0.03439689, -0.3392849, -0.5648054, -0.420242, 0.3731014, 1.150299, 
    0.95733, 0.7633193, 0.5592666, 0.285439, 0.2435114, 0.0816462, 
    -0.03026772, -0.05907631, 0.02510345, 0.240631, 0.460943, 0.6612196, 
    0.843446, 0.9303277, 0.9106989, 0.7832574, 0.6979873, 0.7581111, 
    0.9217507, 1.031435, 1.041331, 1.082265, 1.113011, 1.100657, 0.868463, 
    0.749062, 0.7204649, 0.6846247, 0.7327862, 0.6641011, 0.7126367, 
    0.7077041, 0.6736546, 0.6135826, -0.04639721, -0.236599, -0.23266, 
    -0.1416933, 0.04800367, -0.05435604, -0.04976624, 0.1797911, 0.278554, 
    0.08314347, -0.3668728, -0.1591573, 0.03472233, 0.06530523, 0.06068303, 
    -0.02535214, 0.001242757, 0.01006424, 0.1461971, 0.2028055,
  0.207346, 0.1389213, 0.02323151, 0.1486225, 0.1997452, -0.03628963, 
    -0.03864968, 0.1304096, 0.1417703, 0.1890033, -0.0955019, -0.3950462, 
    -0.08586633, -0.08744526, -0.01589584, 0.1009662, 0.175673, 0.2636123, 
    0.3079644, 0.5181535, 0.5597875, 0.3651423, 0.2218158, 0.1013246, 
    0.1239319, 0.1952047, 0.2044005, 0.1884494, 0.140419, 0.1261287, 
    0.1432347, 0.07588482, 0.1803768, -0.175092, -0.4222599, -0.276996, 
    -0.3292747, -0.5334738, -0.2164329, 0.385699, 0.8859923, 0.914036, 
    0.5624573, 0.4707911, 0.1493225, -0.1594834, -0.0122335, -0.1247334, 
    -0.25141, -0.02305746, 0.273329, 0.5841856, 0.8617575, 1.048476, 1.22219, 
    1.227708, 1.100949, 1.052528, 1.079432, 1.107151, 1.061204, 1.019195, 
    0.9391335, 0.9226296, 0.8817116, 0.8502175, 0.6190326, 0.6389543, 
    0.678635, 0.6669981, 0.7569404, 0.6481347, 0.6991749, 0.5033588, 
    0.3764052, 0.3875713, -0.006667137, -0.04161203, -0.07727271, -0.1540308, 
    -0.2834251, -0.1046655, 0.1301166, 0.2632056, 0.2934953, -0.1826277, 
    -0.8115993, -0.3686633, -0.1097434, -0.09299535, -0.03796595, 
    -0.00686276, 0.1087136, 0.1374569, 0.2533264, 0.1776104,
  0.1531143, 0.07855415, 0.02897739, 0.101536, -0.03796637, -0.3643007, 
    -0.2546327, 0.1448302, 0.1165099, 0.1899148, -0.2329042, -0.5687277, 
    -0.2292911, -0.2556093, -0.02527118, 0.03989816, 0.1938045, 0.4494522, 
    0.3942442, 0.4462464, 0.3295796, 0.2572007, 0.1795144, -0.0006775856, 
    0.01618481, 0.08565044, 0.06211424, 0.04722261, 0.04225826, -0.03433704, 
    -0.04880619, -0.1984639, -0.4232852, -0.6348411, -0.5898704, -0.2460226, 
    -0.3400819, -0.4135845, 0.1219785, 0.7453021, 0.7029362, 0.3956761, 
    0.2315984, 0.03076792, -0.1196551, -0.1064234, 0.07207656, 0.08078432, 
    0.2040913, 0.5879614, 0.9223524, 1.06716, 0.9644909, 1.024045, 1.262652, 
    1.26275, 1.069911, 0.965956, 0.9316136, 0.8321998, 0.7285703, 0.6711159, 
    0.6147195, 0.6929908, 0.6400613, 0.6386774, 0.6174858, 0.6396708, 
    0.5333557, 0.5456936, 0.5768621, 0.4848204, 0.5197158, 0.2911677, 
    0.4203839, 0.4059954, 0.3220108, 0.0112527, -0.09162867, -0.2116642, 
    -0.142035, 0.02069247, 0.08822209, 0.1188046, -0.1852645, -0.4978298, 
    -0.634727, -0.2266705, -0.04356501, 0.03644776, 0.1219132, 0.1210179, 
    0.1997783, 0.151536, 0.2012429, 0.108583,
  -1.096725e-005, -0.01566887, -0.1596127, -0.1798608, -0.267914, -0.2103131, 
    0.06769782, 0.1169819, -0.0964296, -0.01822323, -0.3237898, -0.2281027, 
    -0.07055062, -0.3187606, 0.02840757, 0.1303446, 0.3424377, 0.5233622, 
    0.3451557, 0.2358949, 0.1216695, 0.05794883, -0.1047955, -0.08199239, 
    -0.02899742, -0.06807709, -0.03336048, -0.110867, -0.2070255, -0.3063745, 
    -0.3125758, -0.4072697, -0.4902287, -0.4842228, -0.3820092, -0.2630151, 
    -0.2534283, -0.1522241, 0.117242, 0.3692279, 0.3348527, 0.01659155, 
    0.1475492, 0.009885073, 0.06694961, 0.06755161, 0.05969, 0.3479548, 
    0.5911512, 0.7850482, 0.8399311, 0.8407934, 0.7011778, 0.9077042, 
    1.067047, 0.8444883, 0.6236713, 0.5451718, 0.545481, 0.5388243, 
    0.4652891, 0.4174213, 0.3597385, 0.4620172, 0.4244684, 0.4006572, 
    0.4100971, 0.4006736, 0.374095, 0.4057033, 0.380393, 0.4292212, 
    0.3584857, 0.2609591, 0.3686581, 0.1754286, -0.1017681, 0.05134034, 
    -0.004014492, -0.03677791, 0.01261988, -0.08106501, 0.005865321, 
    0.117877, -0.2798606, -0.2533306, -0.2231711, -0.1773706, 0.009348154, 
    0.06118727, 0.1008687, 0.0767312, 0.07896113, 0.02634048, 0.03861332, 
    0.0167861,
  -0.06194067, 0.0108459, -0.1702905, -0.1742128, -0.01600969, 0.07446873, 
    0.131223, -0.02670324, -0.08251363, -0.04346734, -0.01369846, 0.2587461, 
    0.3707575, 0.5065334, 0.6672106, 0.460325, 0.5634983, 0.4684627, 
    0.2106664, 0.08176017, 0.03612256, 0.1093485, -0.04486704, -0.1073017, 
    -0.09859467, 0.01154542, 0.02910709, -0.1483183, -0.2541447, -0.3085067, 
    -0.3128197, -0.2948347, -0.3430607, -0.3221623, -0.1791445, -0.2007757, 
    -0.2431093, 0.007590771, 0.08607316, 0.126682, 0.06190395, -0.0808208, 
    0.3557515, 0.2338274, 0.2788792, 0.2439022, 0.4158261, 0.9039447, 
    0.8384336, 0.6599506, 0.7332743, 0.7636615, 0.6628314, 0.8166562, 
    0.747711, 0.5610085, 0.5499896, 0.5552468, 0.4869525, 0.4400939, 
    0.3913144, 0.4385308, 0.4837292, 0.4227107, 0.3830791, 0.4073303, 
    0.3674052, 0.3385479, 0.3289616, 0.3214259, 0.2788315, 0.27984, 
    0.1612525, 0.274436, 0.2120178, -0.1128521, 0.005051494, 0.008892596, 
    0.110211, 0.07474552, 0.03836857, 0.04616481, 0.04128198, -0.09421611, 
    -0.502696, -0.368142, -0.09542072, -0.07608473, 0.07809854, -0.004291296, 
    0.05405879, 0.06939101, 0.04050088, 0.03960586, -0.01350307, 0.00702095,
  -0.02403426, -0.03127718, -0.2016054, -0.07409883, -0.04558325, -0.1805118, 
    -0.04120529, -0.07688212, -0.1037213, -0.1076601, 0.2985575, 0.7726617, 
    0.6392796, 0.4896538, 0.4152886, 0.2844619, 0.1994687, 0.1308162, 
    0.1729549, 0.1930559, 0.1372616, 0.02585208, -0.181879, -0.2302027, 
    -0.1088154, 0.09188437, -0.1182225, -0.1832132, -0.2100037, -0.5017844, 
    -0.5174422, -0.2515244, -0.121853, -0.3538516, -0.215017, 0.1134009, 
    0.05700445, 0.1156958, 0.02713811, 0.05693948, 0.06638002, 0.3321187, 
    0.5389051, 0.2510962, 0.260097, 0.3938861, 0.8576557, 1.439492, 1.389752, 
    1.144553, 1.190696, 1.184055, 1.039443, 1.044488, 0.8773171, 0.8069394, 
    0.7107319, 0.5818419, 0.5002013, 0.5224505, 0.5836322, 0.6123106, 
    0.6418513, 0.6203179, 0.626047, 0.6059468, 0.5922263, 0.6034892, 
    0.4829326, 0.4250712, 0.3550518, 0.1902246, 0.2015367, 0.06299448, 
    -0.1564555, 0.03161402, 0.03369734, 0.03817326, 0.05576766, 0.08268824, 
    0.1117898, 0.0384825, -0.1360943, -0.2214948, -0.2427677, -0.6540471, 
    -0.4168398, -0.1555281, -0.0640893, 0.004823446, 0.09564424, 0.0610733, 
    0.06743765, 0.1076233, 0.03713179, 0.09157515,
  -0.185118, -0.1545191, -0.2551863, -0.04423225, -0.08248106, -0.07214575, 
    0.009397224, -0.03204158, -0.01672583, 0.06965113, 0.1433328, 0.5423719, 
    0.602821, 0.5848692, 0.2519265, 0.08906853, 0.04528588, 0.2373921, 
    0.3601947, 0.09647399, -0.05007559, -0.1978621, -0.3217227, -0.2056421, 
    -0.1111759, -0.009857535, -0.009987831, -0.03117895, -0.1623151, 
    -0.34127, -0.1029238, -0.07771218, -0.1091411, -0.5832789, -0.5348086, 
    -0.06532615, -0.04815488, -0.04867572, -0.09747125, -0.2234155, 0.110162, 
    0.5228735, 0.4428932, 0.2804097, 0.0746967, 0.01703069, 0.5867083, 
    0.8350807, 0.7291398, 0.577545, 0.5019589, 0.5081113, 0.4319232, 
    0.3757546, 0.2841856, 0.225299, 0.1595274, 0.1327208, 0.1293028, 
    0.1452696, 0.2288634, 0.2826557, 0.2843645, 0.3187717, 0.3677626, 
    0.3861873, 0.2941461, 0.1937723, 0.1571839, 0.07941675, -0.03918648, 
    -0.2424581, -0.2254984, -0.4465108, -0.5012637, -0.1158306, 0.009429771, 
    0.08356714, 0.03778262, 0.06483342, -0.06695369, -0.2928652, -0.2902941, 
    -0.3125429, -0.2952256, -0.7605572, -0.6667258, -0.4552349, -0.3898868, 
    -0.2614686, -0.2379988, -0.1997826, -0.1150661, -0.115001, -0.1153591, 
    -0.1277776,
  -0.2895777, -0.2361594, -0.296023, -0.02593808, 0.05952743, 0.05999944, 
    0.03330673, 0.06205022, 0.256321, 0.2288308, 0.1648985, 0.2847065, 
    0.4002013, 0.65108, 0.3492246, 0.3847065, 0.6107319, 0.4910216, 
    0.4015684, 0.1301166, -0.1879823, -0.3171327, -0.4009055, -0.4986106, 
    -0.4612896, -0.3098085, 0.02162063, -0.1036236, -0.7158468, -0.4314557, 
    -0.01780021, 0.01047144, -0.0247499, -0.2219667, -0.4839133, -0.4382592, 
    -0.3061955, -0.1760682, -0.1838644, -0.1694927, 0.1930886, 0.3009825, 
    0.1273009, -0.05796932, -0.4224713, -0.7342225, -0.6949484, -0.8550396, 
    -0.9280866, -0.7924095, -0.6811628, -0.4552839, -0.323269, -0.2671005, 
    -0.2308699, -0.3222271, -0.3772238, -0.4848249, -0.5252382, -0.5104923, 
    -0.5214295, -0.4938421, -0.4502547, -0.479454, -0.4680607, -0.4186468, 
    -0.364512, -0.2999456, -0.1775661, -0.1559188, -0.1009057, -0.1094507, 
    -0.2394311, -0.3424749, -0.1502056, 0.0291075, -0.07196674, -0.02095759, 
    0.04046819, 0.03306258, -0.4735945, -0.3134872, -0.2295845, -0.3144469, 
    -0.4035262, -0.4408795, -0.4414655, -0.4419864, -0.4254174, -0.3423934, 
    -0.2911076, -0.1947371, -0.1788843, -0.2292587, -0.1121037, -0.2382758,
  0.1501848, 0.1052139, 0.1079, 0.1176004, 0.2114155, 0.4011127, 0.4531472, 
    0.4976133, 0.3771543, 0.02730087, -0.00551188, 0.1813211, 0.2559955, 
    0.5112364, 0.2003474, 0.2069393, 0.5539934, 0.3763403, 0.1625547, 
    0.1876199, -0.008441329, -0.1854921, -0.224278, -0.5143332, -0.5433862, 
    -0.5268497, -0.06244516, -0.05062884, -0.6941347, -0.8294699, -0.8110452, 
    -0.2844992, 0.03254151, 0.1725645, -0.3652447, -0.6639426, -0.3886985, 
    -0.08417375, -0.01241267, -0.07750055, 0.02870061, -0.004632682, 
    0.05425397, 0.01888627, -0.1574973, -0.6230898, -1.146999, -1.465261, 
    -1.579649, -1.665814, -1.749783, -1.74949, -1.610118, -1.577045, 
    -1.581846, -1.551377, -1.439496, -1.423562, -1.297374, -1.140847, 
    -0.9926372, -0.8842877, -0.8014101, -0.7528261, -0.6437442, -0.5411727, 
    -0.3862085, -0.1980735, -0.06905332, 0.113922, 0.1432514, 0.177545, 
    0.1015521, -0.1377382, -0.2767196, -0.03891007, -0.1978949, -0.1451114, 
    -0.1080509, -0.279812, -0.2022562, -0.3210876, -0.361095, -0.4838488, 
    -0.3930119, -0.3353783, -0.268842, -0.1616477, -0.08739632, -0.1123477, 
    -0.1026633, -0.1601666, -0.2623476, -0.2369081, 0.07774031, 0.1400287,
  0.2036844, 0.09622988, -0.1004175, -0.2731553, -0.3791933, -0.04052174, 
    0.4022031, 0.6066625, 0.6240778, 0.4373432, 0.1319395, 0.1662169, 
    0.3492898, 0.7484272, 0.769505, 0.4612198, 0.3710183, 0.4393289, 
    0.2108618, 0.1009499, 0.1604388, -0.08790123, -0.1893172, -0.4853297, 
    -0.6100529, -0.8365343, -0.4514917, -0.06827235, -0.20263, -0.420681, 
    -0.593256, -0.6418879, -0.839268, -0.01775128, -0.05147514, -0.6811789, 
    -0.6624941, -0.3046001, 0.000429213, -0.2113059, -0.1987571, -0.1477485, 
    -0.09542072, 0.06486571, 0.1386614, 0.001356363, -0.1378524, -0.3047791, 
    -0.3834736, -0.4784281, -0.5759218, -0.6855083, -0.6368592, -0.6657653, 
    -0.8733664, -0.9065533, -0.8262959, -0.7754009, -0.6773376, -0.6539657, 
    -0.5002873, -0.3578392, -0.3407661, -0.3920031, -0.334418, -0.1794212, 
    -0.003867745, 0.08980095, 0.1156145, 0.3182023, 0.3659074, 0.6325741, 
    0.7534237, 0.1632547, -0.196332, -0.2509382, -0.2774032, -0.3189886, 
    -0.5374289, -0.2408309, -0.08742929, -0.1741152, -0.4356389, -0.3833928, 
    -0.3781188, -0.3453226, -0.1670187, -0.1225362, 0.03937793, 0.1427464, 
    0.2374898, 0.2615781, 0.29164, 0.2419656, 0.2608947, 0.2220274,
  -0.0003685951, 0.02580321, -0.2080023, -0.2623806, -0.4228449, -0.6555271, 
    -0.4252217, -0.2963479, -0.07855844, 0.03219962, 0.06701437, 0.2263243, 
    0.16192, 0.1611547, 0.4570048, 0.6562724, 0.5017314, 0.5592666, 
    0.5993224, 0.4369524, 0.3596413, 0.228961, 0.2140355, -0.05936921, 
    -0.23227, -0.3474548, -0.3270934, -0.2457626, -0.2489359, -0.3776469, 
    -0.002322197, 0.04398441, -0.882839, -0.5263128, -0.08930099, -0.546446, 
    -0.7550884, -0.4098736, -0.06343807, -0.3570907, -0.450336, -0.3596785, 
    -0.2631128, -0.02956784, 0.0287981, -0.02081156, -0.07728934, -0.2084091, 
    -0.08458066, -0.06509805, -0.02738643, 0.08294868, 0.2017965, 0.2630758, 
    0.2354555, 0.2740622, 0.417031, 0.4038472, 0.2649474, -0.01192427, 
    -0.1838968, -0.2620707, -0.3385355, -0.3146913, -0.2996526, -0.1964461, 
    -0.1094995, -0.1251732, -0.1578554, 0.08678961, 0.6360735, 0.8724177, 
    0.6898494, 0.340045, 0.1806369, 0.1422582, -0.1086041, -0.1763941, 
    -0.1491317, -0.06501704, -0.1506454, -0.2879337, -0.2493761, -0.2262146, 
    -0.2111917, -0.1332133, -0.03814483, -0.03148746, 0.1354227, 0.2495675, 
    0.4237528, 0.4946995, 0.3816301, 0.3047749, 0.06281495, -0.04149818,
  -0.1152124, -0.1889105, -0.3320582, -0.3058863, -0.1267035, -0.3705177, 
    -0.6983504, -0.3897235, -0.264008, -0.1959085, -0.1113715, 0.05366806, 
    -0.01706763, -0.03560621, 0.2298071, 0.352268, 0.4951391, 0.639117, 
    0.6344292, 0.3702204, 0.2655333, 0.4643288, 0.6901591, 0.2392147, 
    -0.1776308, -0.05694392, 0.02280879, -0.07590568, -0.2056251, -0.5082626, 
    -0.5520782, -0.03672981, -0.1210895, -0.3750105, -0.4070899, -0.5396423, 
    -0.7240666, -0.3626407, 0.01447517, -0.1040958, -0.2593367, -0.2595483, 
    -0.113943, 0.09250236, 0.1936091, 0.09453702, -0.02575946, -0.170779, 
    -0.20351, -0.2736104, -0.2011333, -0.06436586, 0.01691675, 0.04930639, 
    0.09732056, 0.06574512, 0.1598849, 0.2814672, 0.2559631, 0.07857037, 
    -0.1163507, -0.1625586, -0.3177514, -0.3384862, -0.3890402, -0.367393, 
    -0.1656685, -0.07707739, -0.1728293, -0.1015567, 0.3992407, 0.2879939, 
    0.2859595, 0.9818587, 0.7270079, 0.7375872, 0.5311095, 0.3002013, 
    0.1541564, 0.03690386, -0.03591537, -0.1346948, -0.07466877, -0.1294701, 
    -0.06783295, -0.07431078, -0.03405976, 0.0753479, 0.08197212, 0.07954645, 
    0.1138573, 0.2021546, 0.115387, 0.0807513, 0.1232803, 0.09209561,
  0.07791889, -0.1645774, -0.6518499, -0.8638449, -0.5624783, -0.5247177, 
    -0.7671494, -0.5549085, -0.3577743, 0.03512955, 0.5640688, 0.210992, 
    0.01213145, -0.05334693, 0.3244035, 0.2111062, 0.2401586, 0.4552629, 
    0.4392633, 0.3695862, 0.1807512, 0.2641008, 0.3297098, 0.1638241, 
    -0.02706122, -0.003460854, 0.02106714, -0.1138124, -0.2993922, 
    -0.3174262, -0.3797789, -0.3505149, 0.04072952, -0.09247494, -0.4497013, 
    -0.501621, -0.5353453, -0.2613876, -0.08303463, -0.1557398, -0.2378521, 
    -0.2565209, -0.1603134, 0.0874083, 0.2489643, 0.07917273, 0.04549754, 
    0.02238524, -0.0878849, -0.1639104, -0.2089624, -0.1917259, -0.02798915, 
    0.05716705, 0.1599829, 0.2264378, 0.2662497, 0.3495991, 0.3233454, 
    0.2599506, 0.05554008, -0.1236424, -0.236371, -0.1296005, -0.1792102, 
    -0.3882265, -0.1761825, 0.07424068, 0.04170516, -0.008799314, 0.06602144, 
    -0.1849878, 0.264101, 1.106923, 0.7542374, 0.8517964, 0.8435118, 
    0.6423725, 0.4832579, 0.2492898, 0.1713276, 0.01467061, -0.1151471, 
    -0.1750268, -0.0574162, -0.03975666, -0.003265619, 0.04473209, 
    0.02668238, 0.006484032, -0.08025169, 0.2764049, 0.5634661, 0.4271544, 
    0.1764054, 0.1225648,
  -0.3974223, -0.1119895, -0.4917259, -0.7716088, -0.519835, -0.6923931, 
    -1.009077, -0.9597759, -0.8148048, -0.2854104, 0.1980038, 0.105377, 
    0.1416073, -0.1129823, 0.1545793, 0.1314838, 0.2538307, 0.4441791, 
    0.2050513, 0.1570206, 0.1122777, 0.08387613, 0.214817, 0.1450415, 
    -0.08322974, -0.08876383, -0.01602584, -0.2485294, -0.5886496, 
    -0.6278591, -0.3668399, -0.3015246, -0.08126068, -0.2108345, -0.5437288, 
    -0.6466246, -0.5707293, -0.2572529, -0.08864951, -0.1179142, -0.1904891, 
    -0.242605, -0.2839462, -0.1738549, -0.04926181, -0.05284262, -0.08073962, 
    -0.1598086, -0.1721947, -0.2009709, -0.2932723, -0.3413031, -0.2919216, 
    -0.2702744, -0.1280379, 0.03801024, 0.1493223, 0.2585831, 0.1432836, 
    0.04940367, -0.06402421, -0.2356057, -0.3552837, -0.2810326, -0.2023544, 
    -0.3093858, -0.201117, 0.07035112, 0.138808, -0.07092524, -0.08215541, 
    0.05407465, 0.4419492, 0.8260965, 0.6831601, 0.7228575, 0.696653, 
    0.7006081, 0.6337136, 0.3241921, 0.1571511, 0.04946885, -0.05777399, 
    -0.1794862, -0.1852806, -0.125401, -0.05271244, 0.03089762, 0.06875587, 
    -0.0924418, -0.5621355, -0.5455346, 0.01141524, 0.380507, -0.02601957, 
    -0.5559347,
  -0.7307718, -0.3900985, -0.3652935, -0.6861268, -0.5421002, -0.5490826, 
    -0.7944928, -0.9551539, -1.039756, -0.3141708, -0.1292748, -0.2742291, 
    -0.04035866, 0.06209886, -0.01487023, -0.1130801, -0.06506586, 0.1932026, 
    0.250364, 0.3535053, 0.6017308, 0.3636615, -0.01592851, 0.02090438, 
    -0.09791064, -0.2592716, 0.0119524, -0.07950234, -0.3711365, -0.432497, 
    -0.3761497, -0.2269473, -0.2107849, -0.2984486, -0.2896914, -0.2909932, 
    -0.2972269, -0.2535746, -0.2307558, -0.3097925, -0.3132595, -0.1928003, 
    -0.2434675, -0.3337345, -0.3418885, -0.1868105, -0.09888729, -0.2012473, 
    -0.2017356, -0.2527447, -0.2935976, -0.327761, -0.2962994, -0.1296978, 
    0.09733665, 0.2133035, 0.2664936, 0.399013, 0.3467834, 0.07598281, 
    -0.2430935, -0.4375589, -0.5463152, -0.6374779, -0.3790793, -0.1942649, 
    -0.1708928, -0.09159562, -0.06054097, -0.2655702, -0.237136, 0.2931536, 
    0.6566465, 0.5674862, 0.3757545, 0.3923562, 0.3773333, 0.5351784, 
    0.5252826, 0.2403054, -0.03101619, -0.2002219, -0.2746523, -0.3901958, 
    -0.3874941, -0.2470644, -0.09795955, 0.07240188, 0.1686417, 0.1157936, 
    -0.2872176, -0.8533788, -0.6727803, 0.05397701, 0.3135639, -0.2240341,
  -0.05783904, -0.01231509, 0.03566675, -0.2514426, -0.5632915, -0.9218528, 
    -0.7948834, -1.034906, -1.449734, -0.6906354, -0.3740501, -0.4478945, 
    -0.1332784, 0.01548447, -0.06438208, -0.2158795, -0.2459091, -0.09073311, 
    0.09940371, 0.08377874, 0.021734, -0.2090111, -0.8681421, -0.7519639, 
    -0.4268498, -0.4969504, -0.3010356, -0.1639423, -0.03277421, 0.1523334, 
    0.06997633, 0.09491158, 0.004205227, -0.2624292, -0.1816025, -0.0280385, 
    0.0362854, 0.1187401, 0.02759385, -0.2375596, -0.3375108, -0.3107202, 
    -0.3407329, -0.3726504, -0.4050071, -0.3850527, -0.3167095, -0.3379824, 
    -0.2512472, -0.2895448, -0.441856, -0.5267521, -0.4186794, -0.2188747, 
    -0.07722414, 0.134869, 0.2308816, 0.1931049, 0.1206602, 0.01655865, 
    -0.2591414, -0.5263128, -0.721153, -0.7931089, -0.4563737, -0.08532953, 
    -0.1726505, -0.2049908, -0.1570252, -0.1598411, -0.2362896, -0.04460669, 
    0.1445697, 0.1833393, 0.1654845, 0.1918191, 0.1743872, 0.3149799, 
    0.4156961, 0.2684467, -0.06734432, -0.3215109, -0.3714784, -0.4692487, 
    -0.6413516, -0.6733828, -0.3819113, 0.07232037, 0.4207742, 0.4738341, 
    0.1185116, -0.5004503, -1.078135, -1.072195, -0.3194114, 0.03179306,
  -0.08495504, 0.04854108, 0.05900659, -0.0853132, -0.3532818, -0.4364851, 
    -0.1559836, -0.2960554, -0.656944, -0.7391706, -0.5922467, -0.5056746, 
    -0.09107479, 0.01543558, -0.05453509, -0.05492571, -0.08296932, 
    -0.04577857, 0.08166283, -0.04618548, -0.3384708, 0.03993118, 0.1569556, 
    -0.06387752, -0.2506287, -0.2083927, -0.04765022, -0.1469178, -0.2714133, 
    -0.1413189, -0.1697696, -0.04320717, 0.08962202, -0.0009865761, 
    0.1196837, 0.3008692, 0.1754614, 0.1672746, 0.286952, 0.168577, 
    -0.05114985, -0.2036725, -0.2525331, -0.2420351, -0.2283469, -0.1988873, 
    -0.2095808, -0.2984806, -0.2652775, -0.1952416, -0.2910423, -0.4382428, 
    -0.3732364, -0.2265406, -0.1036727, 0.1051977, 0.300494, 0.3144424, 
    0.1729709, 0.01320577, -0.2273541, -0.5271752, -0.7439072, -0.7391541, 
    -0.5073351, -0.2818302, -0.07087624, 0.04924098, 0.07928655, 0.034495, 
    -0.07234097, -0.1183208, 0.004497886, 0.1460669, 0.1880593, 0.1235574, 
    0.04670173, 0.2043189, 0.3884174, 0.2760313, 0.02375251, -0.1266544, 
    -0.286534, -0.4336044, -0.5407658, -0.6357037, -0.5993106, -0.2665471, 
    0.3187885, 0.7361876, 0.5496967, 0.02241808, -0.5053489, -1.033637, 
    -1.028933, -0.4098899,
  -0.3847108, -0.2101341, -0.2145123, -0.2489687, -0.2503684, 0.01248971, 
    0.3893452, 0.573541, 0.2871153, -0.1141542, -0.4639263, -0.4523703, 
    -0.1609969, -0.04566463, -0.1144146, -0.0233339, -0.05072648, 
    -0.09878957, 0.1737847, 0.4183813, 0.09512293, 0.2560443, 0.5503152, 
    0.2922748, 0.1928608, 0.3258848, 0.4047585, 0.1244526, -0.1050234, 
    -0.1228131, -0.2900169, -0.4153914, -0.3120223, -0.2108018, 0.03011632, 
    0.1447158, 0.1093645, 0.09758081, 0.2178768, 0.286546, 0.1471899, 
    -0.06731176, -0.2141379, -0.2683209, -0.2341737, -0.1429793, -0.09157956, 
    -0.1283306, -0.1571071, -0.0565536, -0.03542733, -0.1080999, -0.1298118, 
    -0.1534607, -0.2139425, -0.2075784, -0.16155, -0.06262398, -0.0322535, 
    -0.1405869, -0.3765897, -0.7582948, -0.8445253, -0.4368593, -0.214675, 
    -0.3473573, -0.1467875, 0.1706602, 0.1218972, -0.006992757, 0.04509059, 
    0.07523358, 0.0689187, 0.1704323, 0.2703507, 0.2260308, 0.06777942, 
    0.1352274, 0.4200418, 0.4405333, 0.3796934, 0.3121476, 0.0469296, 
    -0.166726, -0.149994, -0.1734804, -0.3046005, -0.2648382, 0.1491103, 
    0.6545465, 0.714784, 0.3904519, -0.03933316, -0.5045187, -0.6426862, 
    -0.6194766,
  -0.3290631, -0.4804469, -0.3837506, -0.0315533, 0.196523, 0.267698, 
    0.3631896, 0.6374408, 0.8515033, 0.667177, 0.3517962, 0.1366268, 
    0.1706601, 0.142877, 0.03740829, 0.03329045, 0.00430283, -0.1000428, 
    -0.01387787, 0.2004775, 0.2105038, 0.1694558, 0.187929, 0.05498642, 
    0.02342717, 0.169472, 0.2409728, 0.2010964, 0.1339089, 0.06193629, 
    -0.1593853, -0.358832, -0.3528425, -0.1600201, -0.03313208, -0.001068473, 
    0.03718066, 0.1804419, 0.2412983, 0.3041889, 0.2988991, 0.1401915, 
    -0.1480083, -0.3807885, -0.4782817, -0.35587, -0.1236925, 0.04232359, 
    0.1116109, 0.2256083, 0.3803935, 0.514606, 0.5762596, 0.5243881, 
    0.4152567, 0.3115296, 0.1152737, -0.09857774, -0.171201, -0.1462667, 
    -0.3256776, -0.7750921, -0.9807067, -0.4621196, -0.1189067, -0.1739039, 
    -0.1564398, -0.03222084, -0.02701229, -0.1053001, -0.033539, 0.04043543, 
    0.000428915, 0.1067111, 0.364557, 0.4469457, 0.2723688, 0.1724506, 
    0.3183816, 0.4183978, 0.393821, 0.4304421, 0.4061581, 0.2501196, 
    0.1662815, 0.143609, 0.1183813, 0.1518123, 0.3550191, 0.6208231, 
    0.7678607, 0.6326721, 0.2595758, -0.09278417, -0.2520127, -0.2849551,
  0.1094456, 0.1803442, 0.2524799, 0.1599181, 0.2004617, 0.2629127, 
    0.1997128, 0.3955952, 0.7532122, 0.8201556, 0.7336968, 0.6127822, 
    0.3900447, 0.3363826, 0.25899, 0.04777586, -0.01224995, 0.02726832, 
    -0.007529885, 0.02407789, 0.2847387, 0.4043025, 0.3823622, 0.2236876, 
    0.01130152, -0.09107482, -0.1237896, -0.02551508, 0.08503181, 0.04867131, 
    0.03524357, 0.02858651, 0.01444268, 0.1372292, 0.2399148, 0.1929746, 
    0.187571, 0.3428121, 0.397939, 0.3494035, 0.2900125, 0.204547, 
    0.06397086, -0.1733505, -0.4163351, -0.4488876, -0.2635031, -0.07312226, 
    0.07096958, 0.324306, 0.6053934, 0.7862039, 0.9310291, 1.035878, 
    1.017632, 0.8377991, 0.5233459, 0.1914773, 0.0722723, 0.02136087, 
    -0.2173433, -0.6401305, -0.7850201, -0.4609971, -0.2053981, -0.09385777, 
    -0.05595088, 0.004400253, 0.009250736, 0.0650613, 0.1898986, 0.1896054, 
    0.1043841, 0.1705135, 0.2089901, 0.3166721, 0.3527073, 0.2501034, 
    0.1807514, 0.2407448, 0.2140684, 0.2328673, 0.2629126, 0.2909724, 
    0.3546278, 0.3811576, 0.2372777, 0.1129775, 0.2961161, 0.5968812, 
    0.6505105, 0.4741924, 0.3296611, 0.2606833, 0.1378803, 0.0645411,
  0.1188531, 0.5407286, 0.5917382, 0.3666396, 0.2956109, 0.3518125, 
    0.4365453, 0.7096571, 0.9710508, 0.9899634, 0.9970433, 0.8926654, 
    0.667258, 0.5738502, 0.5184138, 0.2799045, 0.0669328, 0.03317642, 
    -0.02144611, -0.1482202, -0.1781193, -0.1448019, -0.1293397, -0.1458273, 
    -0.04774785, -0.1329858, -0.1606063, -0.1376405, -0.06669328, 
    -0.01337296, 0.04129803, 0.007997036, -0.02582455, 0.003748894, 
    0.0389055, -0.01674211, -0.05686254, 0.1454973, 0.3933005, 0.3232322, 
    0.1079972, 0.05101478, 0.1442441, 0.1149148, -0.1608827, -0.3682235, 
    -0.3021427, -0.1056581, 0.0948298, 0.3469458, 0.5987854, 0.8232157, 
    1.074127, 1.36529, 1.472907, 1.262425, 0.8765855, 0.4828675, 0.221426, 
    0.1188865, 0.02500534, -0.03728294, -0.01752305, 0.01260376, 0.1305726, 
    -0.068923, -0.06254292, 0.1061093, 0.2253804, 0.3520405, 0.4160377, 
    0.3584694, 0.2887427, 0.266119, 0.2476783, 0.3685602, 0.4949763, 
    0.4323625, 0.2847553, 0.2074766, 0.2953347, 0.2536355, 0.2366272, 
    0.2569555, 0.3629127, 0.5449599, 0.4482638, 0.1117404, -0.05573988, 
    0.1135798, 0.2167053, -0.0009217262, -0.1882427, -0.1995707, -0.2523704, 
    -0.2266374,
  0.1123922, -0.007089853, 0.184284, 0.4778223, 0.5724671, 0.3527076, 
    0.3592999, 0.7942607, 1.284348, 1.392095, 1.300299, 1.21078, 1.103521, 
    0.9911032, 0.9150777, 0.7465062, 0.441607, 0.3073785, 0.3183005, 
    0.2628312, 0.06746984, -0.1049743, -0.1268988, -0.07572651, -0.009499073, 
    -0.06252646, 0.02056241, -0.0179956, -0.05875057, -0.0114361, 
    -0.01819068, -0.02699649, 0.03371346, 0.06856012, 0.07033467, 
    -0.01980186, -0.107986, 0.03224897, 0.09048414, -0.04859447, -0.1927185, 
    -0.09963584, 0.1336974, 0.3233781, 0.2126846, 0.005978942, -0.06871152, 
    0.05897404, 0.3188862, 0.5782775, 0.7631245, 0.9124082, 1.085716, 
    1.229612, 1.321913, 1.300332, 1.095156, 0.7008038, 0.3236232, 0.1356015, 
    0.1998105, 0.3092508, 0.4463439, 0.5283265, 0.2851787, -0.02291107, 
    -0.119965, 0.01843053, 0.2311258, 0.4283587, 0.5482969, 0.6635475, 
    0.8372781, 0.8754453, 0.7804254, 0.7745987, 0.8805716, 0.8064022, 
    0.7311907, 0.5985247, 0.4050353, 0.4132223, 0.2948954, 0.2594785, 
    0.4283751, 0.79247, 0.9512591, 0.5521538, -0.04325616, -0.2912053, 
    -0.2440209, -0.3334091, -0.475287, -0.3619895, 0.009446144, 0.204206,
  -0.5515568, -0.5364368, -0.261029, 0.1727438, 0.2330623, -0.04896903, 
    -0.1021912, 0.3603413, 0.9187068, 1.226812, 1.342519, 1.4148, 1.305881, 
    1.26275, 1.158909, 1.057379, 0.9146049, 0.800331, 0.7688855, 0.7293509, 
    0.661659, 0.4967997, 0.2882223, 0.09279585, 0.05360317, 0.03700161, 
    0.01094294, -0.01537514, -0.02115309, -0.09350014, -0.05058038, 
    -0.02548236, 0.02653563, 0.09203053, 0.07858664, 0.01551652, 0.1291406, 
    0.1269746, 0.2811093, 0.113287, 0.005131721, 0.03975201, 0.03651333, 
    0.04837847, 0.3416557, 0.297873, 0.184185, 0.08809209, 0.2353899, 
    0.6598042, 1.195204, 1.552089, 1.637718, 1.535764, 1.309918, 1.177529, 
    0.9591204, 0.6140189, 0.3310933, 0.3395569, 0.4793193, 0.7041402, 
    0.5366762, 0.3536189, 0.1670954, 0.1608293, 0.1457739, 0.1331438, 
    0.2139708, 0.3594299, 0.4893939, 0.7171609, 0.8876362, 0.9696674, 
    0.9025776, 0.7514382, 0.7021376, 0.7732476, 0.8597715, 0.8158752, 
    0.7569231, 0.5558487, 0.3454647, 0.3295956, 0.5353085, 0.9114966, 
    1.118186, 0.9338926, 0.4279193, -0.04813886, -0.3526146, -0.7023377, 
    -1.04407, -1.121056, -0.8349719, -0.4984477,
  -1.336291, -0.9957132, -0.5050075, -0.1641707, -0.2457134, -0.4089783, 
    -0.337901, -0.1644149, 0.126243, 0.433697, 0.7416719, 1.036773, 1.086887, 
    0.9227432, 0.9230036, 1.062782, 1.095253, 1.056321, 0.9046767, 0.7882704, 
    0.7676973, 0.6625054, 0.4514539, 0.2760472, 0.1363337, 0.1040257, 
    0.09437418, 0.04735279, 0.01063395, -0.0228132, 0.03397381, -0.02230853, 
    -0.0795188, -0.1174257, -0.1009381, -0.1190207, -0.1431423, -0.0282979, 
    -0.1599708, -0.06309652, -0.1612248, -0.03056002, -0.180284, -0.4426861, 
    -0.3449645, -0.1506786, -0.07717562, 0.1963925, 0.3887758, 0.8533254, 
    1.426585, 1.699159, 1.428603, 1.078912, 0.7443094, 0.5327696, 0.4490945, 
    0.3659565, 0.1994363, 0.0703671, 0.1945695, 0.3049371, 0.2629287, 
    0.01608646, 0.03744096, 0.09487899, 0.05648392, -0.03725004, -0.00440526, 
    0.1531309, 0.4618224, 0.7408748, 0.812685, 0.8856343, 0.9083878, 
    0.9439349, 0.8554748, 0.8682677, 1.028066, 1.07958, 1.059413, 0.7084695, 
    0.2771704, 0.03530848, 0.07817972, 0.3180394, 0.4898982, 0.4762104, 
    0.2102273, -0.1951112, -0.5782004, -0.9601668, -1.356358, -1.658718, 
    -1.763031, -1.63253,
  -1.559515, -1.509565, -1.385298, -1.143972, -0.8595321, -0.6759219, 
    -0.4965763, -0.3253684, -0.1729923, 0.09185135, 0.3724993, 0.666249, 
    0.8573786, 0.9431044, 0.9279841, 0.9207898, 0.8990124, 0.8930721, 
    0.8350482, 0.7296609, 0.6541071, 0.5948296, 0.5171441, 0.3976617, 
    0.2832088, 0.2196506, 0.1786029, 0.1830137, 0.2024148, 0.08600855, 
    0.07671505, 0.08436453, -0.04532278, -0.1264914, -0.08585018, -0.073399, 
    -0.1545513, -0.270274, -0.3487896, -0.2316027, -0.1963644, -0.2052991, 
    -0.4540625, -0.7288837, -0.8119731, -0.7113869, -0.7625589, -0.3565049, 
    0.1919813, 0.7899957, 1.387034, 1.764686, 1.595807, 1.03246, 0.5575581, 
    0.3372944, 0.2520404, 0.2233296, 0.1213274, 0.05298424, -0.001166105, 
    0.1004452, 0.1624732, 0.1141009, -0.01936245, -0.1133893, -0.1935813, 
    -0.2684511, -0.1666771, 0.06297791, 0.2792377, 0.4452045, 0.5124243, 
    0.4158912, 0.2698786, 0.3999733, 0.5538797, 0.4935444, 0.6383196, 
    0.9258199, 1.260634, 1.166136, 0.5440326, 0.1586811, -0.03161848, 
    -0.07131553, 0.03586197, 0.1373587, 0.0363493, -0.1822531, -0.3991313, 
    -0.6333278, -0.8916446, -1.119802, -1.33419, -1.503038,
  -0.9614037, -1.270144, -1.448285, -1.431455, -1.263845, -0.9773052, 
    -0.7347763, -0.5787215, -0.4168724, -0.1673933, 0.1399797, 0.4215879, 
    0.6474828, 0.6913304, 0.6498102, 0.6406956, 0.6488172, 0.6853895, 
    0.6586973, 0.6117083, 0.4883685, 0.3549858, 0.2282612, 0.1838276, 
    0.1609762, 0.06859279, 0.0253638, 0.01340109, -0.03082088, -0.02556372, 
    -0.01716527, -0.08008845, -0.1416444, -0.1431746, -0.1382591, -0.1247661, 
    -0.1033306, 0.0112364, -0.08515021, -0.139024, -0.1844995, -0.1919701, 
    -0.2976993, -0.3782982, -0.3481876, -0.5328395, -0.7864685, -1.026165, 
    -0.9487896, -1.439741, -1.255025, -0.264513, 0.2377665, 0.6231015, 
    0.4906961, 0.3688211, 0.3224181, 0.3086649, 0.3551167, 0.3130268, 
    0.3162494, 0.3099343, 0.2717996, 0.1404683, -0.004844189, -0.18253, 
    -0.3405865, -0.3386008, -0.1942649, -0.01317781, 0.1699441, 0.2977599, 
    0.3796121, 0.4540911, 0.3073788, 0.3954809, 0.2312232, 0.3076392, 
    0.5504777, 0.8775123, 1.157135, 1.050819, 0.4375217, 0.0368222, 
    -0.2999614, -0.4713159, -0.3645279, -0.1111932, 0.07404566, 0.06107283, 
    -0.3405533, -0.2176704, -0.01216841, -0.0651145, -0.2572862, -0.5641868,
  -0.1882433, -0.4747174, -0.7365663, -0.908767, -0.9719503, -0.9064555, 
    -0.7378196, -0.5132591, -0.2330507, 0.1151913, 0.4607806, 0.7061257, 
    0.8033426, 0.8049538, 0.7494362, 0.3532447, 0.5225807, 0.5399473, 
    0.5848203, 0.4781635, 0.475071, 0.3907281, 0.3039119, 0.1741109, 
    0.02985573, -0.07530355, -0.1251897, -0.08591527, -0.007383384, 
    0.09050074, 0.1699441, 0.1251199, -0.04887104, -0.206309, -0.351231, 
    -0.4045188, -0.3095481, -0.2447205, -0.2456809, -0.2301211, -0.3514915, 
    -0.4013776, -0.4017357, -0.3341413, -0.2253522, -0.180642, -0.2199324, 
    -0.3782337, -0.6084573, -0.7562764, -0.7168884, -0.5004821, -0.2775328, 
    -0.1427516, -0.07045329, -0.02030671, 0.02848876, 0.08385992, 0.1521379, 
    0.1982805, 0.1894428, 0.1882872, 0.0821674, -0.1706972, -0.2906353, 
    -0.3779889, -0.4040468, -0.3581321, -0.3174583, -0.03171611, -0.1047304, 
    -0.02750057, 0.2667052, 0.2192117, 0.3111225, 0.3111389, 0.3278865, 
    0.3177794, 0.284202, 0.5483782, 0.9340066, 0.5081111, 0.2396872, 
    0.008990526, -0.06732774, -0.1170025, -0.1176047, 0.0126853, 0.06719303, 
    0.05091619, -0.1890898, -0.6642857, -0.8001084, -0.5252867, 0.1147034, 
    0.08888888,
  -0.09579468, -0.05982518, -0.2826439, -0.4674584, -0.6381289, -0.6850039, 
    -0.5930768, -0.4342226, -0.2325299, -0.07473367, 0.1224994, 0.2382872, 
    0.2586974, 0.1328673, -0.002777256, -0.1889589, -0.2651145, -0.2524843, 
    -0.1549257, -0.01908585, 0.05863225, 0.09930611, 0.1255593, 0.08128846, 
    -0.04058683, 0.005702376, -0.04779673, -0.03492248, -0.01913467, 
    -0.0128033, -0.04328832, -0.1244895, -0.1708925, -0.2381451, -0.2783795, 
    -0.2623476, -0.221983, -0.1780539, -0.1266868, -0.1493918, -0.2459413, 
    -0.3784122, -0.4820254, -0.4978459, -0.4297143, -0.3314885, -0.2251896, 
    -0.1619084, -0.1473738, -0.1586044, -0.1827255, -0.1746038, -0.1510035, 
    -0.1092066, -0.07403409, -0.0260359, 0.03231359, 0.07100189, 0.08932841, 
    0.06768155, 0.005035043, -0.07204831, -0.1443301, -0.1549746, -0.1363872, 
    -0.1215761, -0.09706438, -0.06657931, -0.04024464, -0.05425841, 
    -0.1024355, -0.1623639, -0.1771588, -0.1837668, -0.06675838, -0.09745499, 
    -0.06089902, 0.05877873, 0.2550515, 0.269, 0.1969621, 0.1384823, 
    0.09969687, 0.1197002, 0.1335018, 0.08835208, 0.06818628, 0.1258196, 
    0.1290913, 0.03348637, -0.008929729, -0.07183695, -0.03187799, 
    -0.02569389, -0.08150434, -0.2375591,
  0.2216694, 0.1603898, 0.118121, -0.09727597, -0.3817974, -0.4731549, 
    -0.4932232, -0.4054953, -0.3781679, -0.34197, -0.3230247, -0.3242779, 
    -0.3748801, -0.430593, -0.4875429, -0.5335064, -0.582123, -0.6067812, 
    -0.6053163, -0.5821067, -0.5284609, -0.4576764, -0.3823834, -0.3053489, 
    -0.2150494, -0.1163189, -0.06602597, -0.1109804, -0.07903054, 
    -0.06449601, -0.1024517, -0.1477317, -0.202468, -0.2484804, -0.2594504, 
    -0.2340598, -0.1929628, -0.1457297, -0.09644589, -0.07095759, 
    -0.06244525, -0.07922578, -0.1134868, -0.1341901, -0.1533795, -0.1822532, 
    -0.2063254, -0.2197857, -0.234776, -0.248871, -0.257595, -0.2528099, 
    -0.2334251, -0.1845644, -0.1351015, -0.08124423, -0.04849696, 
    -0.03031635, -0.01609135, 0.006109238, 0.02056229, 0.008794785, 
    0.008827329, 0.007216215, 0.02788675, 0.04486269, 0.05842066, 0.07357365, 
    0.08169538, 0.09557888, 0.06722599, 0.1388406, 0.1295795, 0.07772416, 
    0.127789, 0.1233455, 0.1747779, 0.2141171, 0.2129292, 0.206533, 
    0.1801331, 0.1033425, 0.05796504, 0.01130152, -1.049042e-005, 0.02604723, 
    0.0895079, 0.1744198, 0.2799212, 0.3097386, 0.3120499, 0.3080785, 
    0.3188205, 0.3385472, 0.3285863, 0.2877498,
  0.2810932, 0.2580788, 0.1876525, 0.1227111, 0.06138289, -0.007481039, 
    -0.05536518, -0.09540421, -0.1316347, -0.1609967, -0.1932232, -0.2289491, 
    -0.2699648, -0.3160097, -0.3569276, -0.3945579, -0.4283958, -0.4576438, 
    -0.4867454, -0.5005311, -0.4898052, -0.4737082, -0.4414491, -0.403591, 
    -0.3626242, -0.326524, -0.2754009, -0.2624778, -0.2426535, -0.2357036, 
    -0.249343, -0.2718527, -0.297455, -0.3292583, -0.3536724, -0.3689557, 
    -0.3728944, -0.3575462, -0.3287376, -0.2908795, -0.2493918, -0.2044049, 
    -0.1653098, -0.1319927, -0.09677139, -0.07154354, -0.04511127, 
    -0.01835346, 0.003961086, 0.01348263, 0.02136022, 0.02344352, 0.01939064, 
    0.01867449, 0.01626569, 0.01667255, 0.02803326, 0.03662699, 0.04526967, 
    0.04990828, 0.04504174, 0.04906189, 0.06022722, 0.07528257, 0.1033263, 
    0.1153216, 0.1186745, 0.1067116, 0.07985616, 0.07111597, 0.07256453, 
    0.05093368, 0.0340066, 0.02370381, 0.0448463, 0.08960533, 0.1124408, 
    0.1538471, 0.2400448, 0.2249895, 0.1992081, 0.1796607, 0.1261939, 
    0.1139054, 0.1300352, 0.1564513, 0.183974, 0.2165261, 0.2301818, 
    0.2933491, 0.3343647, 0.3614967, 0.3682186, 0.3522355, 0.3274146, 
    0.3011615,
  0.2667215, 0.2271218, 0.188336, 0.1474832, 0.1036518, 0.05023381, 
    0.00524683, -0.03153702, -0.07471737, -0.1134869, -0.153233, -0.1919211, 
    -0.2275657, -0.264789, -0.302761, -0.3318138, -0.3614198, -0.38808, 
    -0.4126894, -0.4356548, -0.4508241, -0.4600526, -0.4725526, -0.485606, 
    -0.4943462, -0.5030864, -0.5028423, -0.4971132, -0.4893007, -0.4795351, 
    -0.4805442, -0.4858013, -0.4894309, -0.4859315, -0.4802024, -0.4705833, 
    -0.4644634, -0.4523866, -0.4377707, -0.4179302, -0.3946392, -0.3680767, 
    -0.3437278, -0.317914, -0.2866965, -0.2524192, -0.218093, -0.1841738, 
    -0.1498639, -0.1191347, -0.09210017, -0.06526098, -0.03925192, 
    -0.01781631, 0.006076992, 0.02583611, 0.04613233, 0.05630487, 0.0681538, 
    0.07472938, 0.07280874, 0.07074171, 0.07674754, 0.08021438, 0.09079385, 
    0.09492791, 0.09479773, 0.08892202, 0.09310499, 0.1074767, 0.1229877, 
    0.1387104, 0.1579161, 0.1658751, 0.1814024, 0.2018777, 0.2214089, 
    0.237685, 0.2532774, 0.2674702, 0.2836811, 0.2993386, 0.3149962, 
    0.328017, 0.3414773, 0.3542703, 0.3642312, 0.3692442, 0.3739643, 
    0.381435, 0.3877175, 0.3814512, 0.3678608, 0.3483132, 0.3261778, 0.2995014,
  -0.136373, -0.113652, -0.09080005, -0.06770468, -0.04623628, -0.02493095, 
    -0.004960299, 0.009411335, 0.02018619, 0.02822661, 0.03198624, 
    0.03058624, 0.02199221, 0.01011086, -0.005399942, -0.02305949, 
    -0.04174447, -0.06070578, -0.07839793, -0.09312794, -0.1037399, 
    -0.1087692, -0.1095341, -0.1059696, -0.09996378, -0.09210265, -0.0819298, 
    -0.07346654, -0.06711864, -0.06355405, -0.06248045, -0.06357098, 
    -0.06612611, -0.07161117, -0.08087254, -0.09164715, -0.1020799, 
    -0.1150846, -0.1290007, -0.1397591, -0.1466765, -0.1506803, -0.1509082, 
    -0.1462533, -0.1404588, -0.1320772, -0.1224413, -0.1076133, -0.0948205, 
    -0.0770309, -0.06430316, -0.04874313, -0.02955365, -0.01192689, 
    0.0132035, 0.02934945, 0.05171275, 0.07065791, 0.0869177, 0.09471393, 
    0.1073115, 0.1332719, 0.1478877, 0.1571, 0.1635778, 0.1672237, 0.1679561, 
    0.1650427, 0.1567907, 0.1465368, 0.1323441, 0.114001, 0.09228876, 
    0.06168985, 0.04954785, 0.02589887, 0.00322628, -0.02491501, -0.04652959, 
    -0.06980431, -0.09330691, -0.116663, -0.1390426, -0.1609827, -0.1808395, 
    -0.1973434, -0.2111455, -0.2202112, -0.2248497, -0.2250288, -0.2220832, 
    -0.2143843, -0.2040331, -0.1913866, -0.17555, -0.1570437,
  0.1111691, 0.1022825, 0.1107786, 0.1311886, 0.1598184, 0.1893916, 
    0.2162306, 0.2317744, 0.2316769, 0.2161494, 0.1846553, 0.1400916, 
    0.08499718, 0.02666378, -0.0336878, -0.09215131, -0.1444788, -0.1947555, 
    -0.240426, -0.2855921, -0.3223271, -0.3466272, -0.3581995, -0.355872, 
    -0.3443811, -0.3262659, -0.2967086, -0.2621548, -0.2251918, -0.1908655, 
    -0.1597135, -0.1276176, -0.09792948, -0.07712889, -0.07011414, 
    -0.07854509, -0.09709978, -0.1238737, -0.1562304, -0.1979296, -0.2261524, 
    -0.2644005, -0.2930791, -0.3424444, -0.3682259, -0.3567671, -0.3832971, 
    -0.3740848, -0.3430464, -0.2997687, -0.253984, -0.2439091, -0.1946903, 
    -0.1625127, -0.09631799, -0.07362919, -0.0350875, -0.008085579, 
    0.01719117, 0.0554561, 0.09412795, 0.1322302, 0.1667029, 0.1980506, 
    0.2230667, 0.2621619, 0.2820675, 0.2906123, 0.2912471, 0.2718949, 
    0.2608271, 0.2259151, 0.1884153, 0.1560746, 0.1136594, 0.06732142, 
    0.01852584, -0.0201298, -0.0447067, -0.06324506, -0.08022094, 
    -0.08129519, -0.07535444, -0.05925745, -0.04317672, -0.02026007, 
    0.007327855, 0.04193074, 0.07612664, 0.104626, 0.1239295, 0.1399773, 
    0.1489133, 0.1507522, 0.1433468, 0.1271849,
  -0.1187792, -0.2102506, -0.2519329, -0.2402468, -0.1866174, -0.1045049, 
    -0.02278268, 0.02604529, 0.03397173, 0.01424515, -0.007890284, 
    -0.03788698, -0.09024698, -0.1626265, -0.2459274, -0.3204879, -0.3686487, 
    -0.3918095, -0.3878382, -0.3641566, -0.3361942, -0.3040978, -0.2670861, 
    -0.2287723, -0.1903283, -0.1707321, -0.1733851, -0.1928349, -0.2151656, 
    -0.2282192, -0.2268518, -0.2110643, -0.1862755, -0.1574018, -0.126754, 
    -0.09701777, -0.07017851, -0.06213808, -0.07740521, -0.1185184, 
    -0.1752243, -0.2297331, -0.2594203, -0.3030237, -0.3035282, -0.3385706, 
    -0.3215457, -0.2846155, -0.2413538, -0.2121058, -0.1735153, -0.1391402, 
    -0.1084762, -0.0687952, -0.01181275, 0.05273801, 0.09150749, 0.1169471, 
    0.1476111, 0.1795121, 0.2303748, 0.2830763, 0.3324091, 0.3726599, 
    0.4050328, 0.4280472, 0.4275753, 0.4116572, 0.3838904, 0.3440306, 
    0.2898797, 0.2293332, 0.1630242, 0.1038771, 0.05998063, 0.02244806, 
    0.02824259, -0.01147103, -0.0439254, -0.07615197, -0.09576464, 
    -0.09205359, -0.07257123, -0.04348596, 0.006725639, 0.06614944, 
    0.1302772, 0.1989131, 0.2465857, 0.2785844, 0.3050817, 0.2949744, 
    0.2540886, 0.1838088, 0.09476304, -0.0109663,
  -0.127275, -0.1833459, -0.2127568, -0.2083136, -0.1753055, -0.1227177, 
    -0.07400355, -0.04312789, -0.04083288, -0.05541646, -0.08817983, 
    -0.1348759, -0.1845342, -0.2284956, -0.2752405, -0.3081508, -0.3042444, 
    -0.2652636, -0.2256148, -0.2006636, -0.2011682, -0.2129682, -0.1806768, 
    -0.1117311, -0.03640604, -0.001379728, -0.0116663, -0.0246383, 
    -0.003967643, 0.02021861, 0.02705443, 0.006074727, -0.01576787, 
    -0.02193648, -0.02110642, -0.01669538, -0.00769484, -0.008395076, 
    -0.02493143, -0.05730486, -0.09307909, -0.1349738, -0.1328905, 
    -0.1206832, -0.1207809, -0.147083, -0.1421027, -0.190719, -0.2604781, 
    -0.3062788, -0.3410934, -0.3360966, -0.2665329, -0.1488894, -0.03632438, 
    0.08291376, 0.1679724, 0.2538285, 0.3066279, 0.2944047, 0.2844763, 
    0.2754106, 0.2561234, 0.2620153, 0.2804398, 0.3089554, 0.3107134, 
    0.2873734, 0.2155308, 0.1109409, -0.01164997, -0.1361455, -0.2288374, 
    -0.25623, -0.2286423, -0.2034309, -0.1348436, -0.05253553, 0.005016685, 
    0.0580765, 0.02583379, -0.0008425713, -0.0444788, -0.07229456, 
    -0.09133752, -0.08738244, -0.05413049, 0.02130896, 0.09997106, 0.1161169, 
    0.1303421, 0.1394242, 0.1259477, 0.1032752, 0.04004252, -0.04941034,
  -0.03887984, -0.03284143, -0.04521123, -0.05263311, -0.07818648, 
    -0.08595014, -0.1194299, -0.1547818, -0.2516075, -0.2627079, -0.2649217, 
    -0.24054, -0.1986129, -0.1287398, -0.05287725, 0.006562948, 0.06898165, 
    0.05801177, 0.0498898, -0.01427042, -0.07499637, -0.104928, -0.106344, 
    -0.02076435, 0.1244988, 0.2745967, 0.3536984, 0.3497107, 0.2587602, 
    0.1386105, 0.05472374, 0.03042364, 0.0442583, 0.06839573, 0.08828473, 
    0.1041377, 0.1064982, 0.07536173, 0.01789141, -0.02808857, -0.04830337, 
    -0.03433871, 0.02038145, 0.1047564, 0.1387246, 0.1598673, 0.05973673, 
    -0.04195619, -0.2175582, -0.3892216, -0.5065393, -0.5107223, -0.4029749, 
    -0.2220341, -0.04016565, 0.08130245, 0.1834672, 0.2464717, 0.2904822, 
    0.3070837, 0.3098668, 0.2605016, 0.1781449, 0.07886106, 0.00737685, 
    -0.02885365, -0.03816354, -0.03136027, -0.02356398, -0.03695929, 
    -0.04177696, -0.07572865, -0.1026493, -0.1043746, -0.1028447, 
    -0.08598262, -0.02781224, 0.02733105, 0.07474315, 0.09414423, 0.05946004, 
    -0.03767538, -0.1033655, -0.1165003, -0.104928, -0.06002242, 0.01349646, 
    0.05731159, 0.06375688, 0.03262082, 0.01592159, -0.04163048, -0.03406212, 
    -0.04607385, -0.05675095, -0.04635054,
  -0.1282353, -0.0903284, -0.0334762, -0.04093063, -0.02976525, -0.03791946, 
    -0.03700805, -0.03212523, -0.05177057, -0.07927692, -0.07545209, 
    -0.06557254, -0.01988569, 0.06640986, 0.1412797, 0.1483599, 0.1079297, 
    0.04779029, -0.03873324, -0.05341434, -0.03235316, 0.001061566, 
    0.06012732, 0.1385453, 0.2350298, 0.2897173, 0.2343624, 0.0905962, 
    -0.07361317, -0.1627245, -0.1559696, -0.121204, -0.1087854, -0.07727528, 
    -0.04845023, -0.03044868, -0.03135991, -0.06807876, -0.1300421, 
    -0.1559211, -0.1322883, -0.07196927, -0.01173151, 0.03447604, 
    -0.004472256, -0.002112269, 5.233288e-005, -0.0631637, -0.2194951, 
    -0.4134241, -0.6319463, -0.7158003, -0.6578088, -0.4804326, -0.3194463, 
    -0.2278447, -0.1231734, -0.025387, 0.07176469, 0.1533891, 0.176615, 
    0.10168, -0.05304, -0.2358036, -0.3443486, -0.3747686, -0.3353804, 
    -0.2167445, -0.0592249, 0.04477903, 0.07654986, 0.1085485, 0.10946, 
    0.04376991, -0.009078413, -0.08993778, -0.1746871, -0.2061162, 
    -0.2184046, -0.1889612, -0.1486455, -0.2051071, -0.3054327, -0.3306279, 
    -0.3210087, -0.2566696, -0.1467412, -0.0378219, 0.02632198, 0.04865271, 
    0.03888708, 0.02508503, -0.02079713, -0.08793575, -0.1366174, -0.1399703,
  -0.369316, -0.2565068, -0.1757287, -0.08949822, -0.01884389, -0.003268003, 
    -0.001200676, -0.06931603, -0.1854293, -0.2597621, -0.3057255, 
    -0.3523889, -0.3640263, -0.3721155, -0.3917606, -0.4452279, -0.4804163, 
    -0.4302862, -0.3552374, -0.2195604, -0.03593409, 0.07824266, 0.05579787, 
    -0.03051394, -0.1318648, -0.176217, -0.1927536, -0.223857, -0.2646773, 
    -0.213945, -0.1420211, -0.1333296, -0.2145797, -0.2822882, -0.3459599, 
    -0.2893193, -0.1987268, -0.2219689, -0.2255986, -0.2301884, -0.2456507, 
    -0.2254521, -0.1943974, -0.244609, -0.2952275, -0.2477666, -0.2271285, 
    -0.337708, -0.5810998, -0.8985803, -1.198727, -1.275029, -1.097945, 
    -0.8963993, -0.6713343, -0.4949183, -0.3589808, -0.2435999, -0.2071253, 
    -0.2193649, -0.3694137, -0.4199019, -0.4854943, -0.5634403, -0.5969364, 
    -0.5734664, -0.5353642, -0.3758753, -0.1695602, -0.02374312, 0.04691118, 
    0.08919632, 0.1235388, 0.1270218, 0.09806678, -0.05968061, -0.1874801, 
    -0.3172164, -0.4055465, -0.3341598, -0.3448694, -0.3709925, -0.337236, 
    -0.3070927, -0.2961715, -0.31943, -0.3734664, -0.4031214, -0.3849573, 
    -0.2648727, -0.1473434, -0.1148564, -0.1681929, -0.3288375, -0.4547977, 
    -0.4682255,
  -0.3544561, -0.2252731, -0.1149378, -0.07450807, -0.00777638, -0.008069277, 
    -0.2035445, -0.316598, -0.372848, -0.3435347, -0.4075484, -0.5937626, 
    -0.7019168, -0.6709275, -0.5589156, -0.4518032, -0.2796189, -0.1079065, 
    0.06105518, 0.1908891, 0.2367548, 0.1634802, -0.03581995, -0.3183068, 
    -0.4977014, -0.4854781, -0.4162723, -0.4542932, -0.590068, -0.7585087, 
    -0.8840621, -0.9747685, -1.055091, -1.113961, -1.033899, -0.8206508, 
    -0.5866989, -0.4090295, -0.3130335, -0.3223271, -0.3455042, -0.3520146, 
    -0.3206995, -0.2345179, -0.2163701, -0.2778935, -0.4178674, -0.6268842, 
    -0.9474245, -1.210788, -1.357207, -1.332679, -1.14028, -0.9149701, 
    -0.7911258, -0.7240033, -0.6910933, -0.6269333, -0.6796025, -0.8733525, 
    -1.095846, -1.178447, -1.077617, -0.9478154, -0.9120894, -0.8866662, 
    -0.8018518, -0.6700484, -0.447262, -0.2665003, -0.2385869, -0.273792, 
    -0.2644332, -0.2287073, -0.2316858, -0.2628056, -0.377568, -0.4985641, 
    -0.535706, -0.5636357, -0.5885543, -0.6211389, -0.6142054, -0.5880498, 
    -0.6019007, -0.6418095, -0.7495732, -0.7850875, -0.6710087, -0.45304, 
    -0.2425257, -0.1138147, -0.1661097, -0.3363896, -0.4967411, -0.4818323,
  -0.4124964, -0.3790491, -0.4770146, -0.5295862, -0.5864547, -0.7365687, 
    -0.9770308, -1.001884, -0.8198205, -0.7141728, -0.9061649, -1.208102, 
    -1.377047, -1.310543, -1.10011, -0.859355, -0.5900517, -0.352747, 
    -0.1965784, -0.1769495, -0.2448206, -0.4553023, -0.7793259, -1.095504, 
    -1.184518, -1.138034, -1.09915, -1.168535, -1.458623, -1.838245, 
    -2.045178, -1.899247, -1.574687, -1.316842, -1.116028, -0.8999151, 
    -0.688945, -0.494544, -0.4603152, -0.5661257, -0.6941532, -0.6894657, 
    -0.5680302, -0.47109, -0.6255496, -0.9358524, -1.168844, -1.235381, 
    -1.286439, -1.385576, -1.472978, -1.511487, -1.420195, -1.234583, 
    -1.11038, -1.041468, -0.9302534, -0.8194625, -0.8419397, -1.007288, 
    -1.208997, -1.301982, -1.277894, -1.270862, -1.245846, -1.241386, 
    -1.066305, -0.876917, -0.7167608, -0.6021123, -0.6086228, -0.6621058, 
    -0.7217576, -0.7366336, -0.7942996, -0.9114386, -1.078561, -1.146969, 
    -1.053789, -0.936764, -0.9164189, -1.007483, -1.104977, -1.227568, 
    -1.323792, -1.332906, -1.232793, -1.003007, -0.6769333, -0.4099085, 
    -0.2209111, -0.2555302, -0.4365035, -0.5645146, -0.5467411, -0.4740524,
  -0.6309531, -0.8178676, -0.9823694, -1.148239, -1.278496, -1.404196, 
    -1.475338, -1.369674, -1.118307, -0.9709601, -1.145586, -1.442737, 
    -1.577145, -1.48027, -1.287838, -1.074524, -0.8392215, -0.7024704, 
    -0.6554488, -0.6712205, -0.8137009, -1.084665, -1.385381, -1.567526, 
    -1.607353, -1.621464, -1.662008, -1.739807, -1.97109, -2.321416, 
    -2.448369, -2.2207, -1.841516, -1.568567, -1.436015, -1.33372, -1.149166, 
    -0.9328091, -0.8432254, -0.8376917, -0.8976525, -0.9890102, -1.058867, 
    -1.146009, -1.390785, -1.613196, -1.628821, -1.441924, -1.350192, 
    -1.415313, -1.46095, -1.479212, -1.394088, -1.173613, -0.9945441, 
    -0.9690557, -0.9671188, -0.8942833, -0.8659467, -0.9243127, -1.131051, 
    -1.337431, -1.455888, -1.454944, -1.431572, -1.354261, -1.267021, 
    -1.129814, -0.891484, -0.7100226, -0.7179815, -0.8653283, -0.8938767, 
    -0.8046025, -0.8409307, -1.091891, -1.346823, -1.379586, -1.186113, 
    -1.106539, -1.232077, -1.326771, -1.403138, -1.548011, -1.636211, 
    -1.535918, -1.282402, -1.022539, -0.8064903, -0.6051232, -0.4928348, 
    -0.5544885, -0.5737268, -0.4473758, -0.3638635, -0.4751589,
  -1.038505, -1.094576, -1.212415, -1.417965, -1.555432, -1.590914, 
    -1.585511, -1.473629, -1.332971, -1.347408, -1.462057, -1.524004, 
    -1.462806, -1.327698, -1.163587, -1.078626, -1.026168, -0.9658009, 
    -0.8767543, -0.7979295, -0.8366337, -0.9809697, -1.234469, -1.479912, 
    -1.654619, -1.880839, -2.127324, -2.332207, -2.527454, -2.6387, 
    -2.559615, -2.305726, -2.060316, -1.884794, -1.759306, -1.614124, 
    -1.319284, -0.9926398, -0.7847946, -0.6435511, -0.6022749, -0.8145473, 
    -1.036895, -1.140214, -1.237887, -1.292705, -1.175013, -1.084648, 
    -1.179505, -1.26095, -1.255058, -1.196822, -1.129033, -1.039482, 
    -1.037187, -1.127487, -1.052324, -0.830742, -0.6958625, -0.7088995, 
    -0.8397752, -1.07944, -1.286178, -1.345651, -1.371302, -1.380628, 
    -1.238099, -1.003496, -0.7745409, -0.6801071, -0.7204065, -0.7821579, 
    -0.7023077, -0.5877728, -0.721334, -1.052779, -1.148385, -0.8737273, 
    -0.5571088, -0.6512983, -1.04596, -1.258199, -1.307012, -1.39028, 
    -1.383248, -1.218421, -1.070097, -0.9715945, -0.8450157, -0.6667931, 
    -0.5460738, -0.5329553, -0.5024703, -0.483476, -0.599834, -0.849313,
  -0.619544, -0.7582645, -0.8487918, -1.013489, -1.182565, -1.245716, 
    -1.238278, -1.185006, -1.12677, -1.097408, -1.041826, -0.9433395, 
    -0.9035606, -0.911894, -0.9160283, -0.8584931, -0.7568002, -0.618974, 
    -0.5219693, -0.5521126, -0.6872358, -0.847343, -1.08538, -1.374199, 
    -1.641272, -1.853674, -2.07441, -2.249573, -2.296513, -2.187855, 
    -2.034209, -1.917102, -1.789238, -1.563278, -1.297783, -1.045114, 
    -0.6941209, -0.3546023, -0.1820436, -0.1048303, -0.1813114, -0.3272917, 
    -0.3319142, -0.3400848, -0.6787729, -0.9060028, -0.8618288, -0.8942833, 
    -1.084876, -1.084827, -0.9149864, -0.9038537, -1.012024, -1.126201, 
    -1.200045, -1.07931, -0.7093226, -0.3316858, -0.3214157, -0.4442347, 
    -0.5697391, -0.7092249, -0.9047816, -1.024882, -1.057711, -0.9675093, 
    -0.7578576, -0.593909, -0.5629194, -0.553447, -0.4898894, -0.4138315, 
    -0.2817507, -0.213424, -0.2324181, -0.1518521, -0.05432606, -0.06191087, 
    -0.1175095, -0.3699509, -0.7960087, -0.9506801, -0.9686486, -1.032142, 
    -0.9301397, -0.6987759, -0.6202602, -0.6130172, -0.5539514, -0.4931771, 
    -0.4577112, -0.3046515, -0.1650193, -0.276201, -0.4318328, -0.5034955,
  -0.0928514, -0.26069, -0.3036425, -0.4172649, -0.5455203, -0.49067, 
    -0.4064417, -0.3506476, -0.2892543, -0.2832808, -0.4059858, -0.5602504, 
    -0.6387823, -0.6699183, -0.6229944, -0.465312, -0.2954063, -0.1962206, 
    -0.2529752, -0.3998339, -0.4778452, -0.5472455, -0.6782675, -0.8741012, 
    -0.9906702, -1.016614, -1.171464, -1.376119, -1.336765, -1.170765, 
    -0.9742475, -0.7418745, -0.565589, -0.3772588, -0.1465132, 0.09796882, 
    0.3096228, 0.4414427, 0.5867553, 0.7171098, 0.6713253, 0.561625, 
    0.5861688, 0.3372917, -0.3095996, -0.5642059, -0.4055467, -0.5184858, 
    -0.8140261, -0.6570437, -0.4422002, -0.5661261, -0.7979296, -0.8024702, 
    -0.5620244, -0.08287418, 0.3114941, 0.35181, 0.08465552, -0.1631472, 
    -0.3076625, -0.3577764, -0.462431, -0.6203249, -0.6354291, -0.5155885, 
    -0.4435351, -0.3900192, -0.3165815, -0.1806602, 0.006579161, 0.1187701, 
    0.3822465, 0.5889034, 0.7475947, 1.248197, 1.567028, 1.128454, 0.4138381, 
    -0.2306279, -0.586357, -0.5152794, -0.2921352, -0.3064905, -0.3007125, 
    -0.1452274, -0.05133092, -0.07476842, -0.1740685, -0.2223759, -0.137871, 
    0.04030299, 0.1735058, 0.09604836, 0.02379894, 0.02705407,
  0.5451531, 0.4098828, 0.318119, 0.3184283, 0.4010129, 0.4081905, 0.3045285, 
    0.2428747, 0.1314488, -0.2298303, -0.6494269, -0.8424118, -0.6816533, 
    -0.3509567, -0.09737611, 0.0591507, 0.1502316, 0.2083848, 0.2008336, 
    0.1880569, 0.2174678, 0.1492386, -0.0009570122, -0.08507109, -0.07130194, 
    -0.02849627, -0.1467578, -0.2496061, -0.1355104, 0.06427789, 0.3401567, 
    0.510339, 0.4323931, 0.4071815, 0.5479366, 0.7910517, 1.084216, 1.403682, 
    1.592598, 1.363822, 1.084037, 1.100394, 0.9995964, 0.6106153, 0.1502964, 
    0.0917356, 0.1642616, -0.08741474, -0.2541628, -0.1629033, -0.1780236, 
    -0.3587691, -0.3218875, -0.05544889, 0.2854526, 0.6136754, 0.7431347, 
    0.6512406, 0.5093302, 0.3322469, 0.1184282, -0.009680271, -0.09796166, 
    -0.2471478, -0.2452111, -0.1667929, -0.1554487, -0.05455351, 0.1665566, 
    0.3481319, 0.5501013, 0.7970902, 1.198994, 1.4703, 1.610258, 2.265726, 
    2.725459, 1.566263, 0.1607134, -0.633525, -0.5939743, -0.2898401, 
    0.01243836, 0.1413285, 0.15487, 0.1700232, 0.09855509, 0.0017941, 
    -0.1335087, -0.09797835, 0.1698925, 0.2908077, 0.357409, 0.4939322, 
    0.5536819, 0.5991895,
  0.8818722, 0.8170283, 0.8746455, 1.065987, 1.279333, 1.148913, 0.8547885, 
    0.5262891, -0.1414028, -0.8361292, -0.7779749, -0.3014288, 0.186169, 
    0.5311399, 0.5467485, 0.5594437, 0.7293818, 0.9255409, 1.038529, 
    1.017695, 0.8318229, 0.5979199, 0.5234084, 0.5926948, 0.6372917, 
    0.6012895, 0.5290567, 0.564473, 0.6586951, 0.9499059, 1.330684, 1.023148, 
    0.4884802, 0.5368037, 0.716638, 1.000167, 1.2321, 1.521976, 1.723995, 
    1.299011, 0.8932815, 0.9942421, 0.690563, 0.3879921, 0.3803911, 
    0.4021361, 0.3482782, 0.1867224, 0.115417, 0.1233436, 0.09583688, 
    0.1527869, 0.3150916, 0.5619826, 0.8017289, 0.9468949, 0.9128616, 
    0.8270056, 0.7250687, 0.5512081, 0.346016, 0.2137729, 0.1440629, 
    0.09800184, 0.1392449, 0.204154, 0.1342322, 0.2138869, 0.3717319, 
    0.5219109, 0.8743851, 1.124629, 1.204805, 1.416329, 1.763285, 2.378455, 
    2.343135, 0.8818066, -0.6204392, -0.5922328, 0.2505733, 0.4511104, 
    0.3710486, 0.2385453, 0.1472206, 0.0557816, -0.3219852, -0.3954393, 
    -0.1310675, 0.1249709, 0.4816768, 0.6775424, 0.8414583, 1.062422, 
    1.117028, 1.020446,
  0.8373246, 0.971895, 1.175622, 1.433874, 1.478503, 1.169518, 0.5850787, 
    0.1620641, -0.3962693, -0.7560346, -0.2701299, 0.2884151, 0.5302283, 
    0.6975623, 0.598506, 0.7078974, 1.003161, 1.156872, 1.134851, 0.9578001, 
    0.7690629, 0.6270547, 0.6393265, 0.7156938, 0.6784866, 0.6255082, 
    0.6367223, 0.7415401, 0.9241574, 1.574076, 1.885355, 1.055488, 0.3429399, 
    0.5692579, 0.647204, 0.8932978, 1.084688, 1.111934, 1.302754, 0.8159704, 
    0.3679721, 0.7063999, 0.7039909, 0.7363644, 0.8625362, 0.7635127, 
    0.6139359, 0.4916215, 0.484167, 0.4702022, 0.5000362, 0.4684444, 
    0.4368038, 0.5374222, 0.6847529, 0.7443233, 0.6037309, 0.6566443, 
    0.7536007, 0.5857296, 0.4319047, 0.278145, 0.2341182, 0.3028357, 
    0.3178259, 0.2948605, 0.2026076, 0.2508824, 0.4216996, 0.5887569, 
    0.8694047, 1.05168, 1.057067, 1.374222, 1.692338, 1.629723, 0.7043982, 
    -0.1481087, -0.3372686, 0.2868689, 0.764538, 0.4194697, 0.3097531, 
    0.2697465, -0.3129197, -0.5847459, -0.729977, -0.5054653, 0.01175523, 
    0.3984413, 0.7106969, 0.9355342, 1.044991, 1.043786, 1.026403, 0.9683141,
  0.7446163, 0.8342154, 0.8858438, 0.9965529, 0.7280474, 0.02938151, 
    -0.7627242, -0.6960901, -0.2400517, -0.11165, 0.2238482, 0.5863806, 
    0.3671257, 0.08050501, 0.08636439, 0.4457556, 0.6459347, 0.6567094, 
    0.6057817, 0.4063839, 0.3892614, 0.3498409, 0.331628, 0.4251013, 
    0.5018592, 0.489473, 0.4930699, 0.6281931, 0.9373899, 1.309183, 
    0.6248407, -0.2586718, -0.3218387, 0.2321491, 0.2967973, 0.4442421, 
    0.7478714, 0.9829788, 1.052152, 0.1769404, 0.04298902, 1.166133, 
    1.564229, 1.507897, 1.287862, 1.052087, 0.8673702, 0.5895545, 0.4072301, 
    0.2961787, 0.2934933, 0.1633337, 0.1060095, 0.1671748, 0.1641638, 
    0.3278193, 0.4314489, 0.6653356, 0.7339554, 0.4973994, 0.4170121, 
    0.419307, 0.485697, 0.5462114, 0.4838741, 0.3646358, 0.2776403, 
    0.3225134, 0.4744015, 0.6545935, 0.8947792, 1.089327, 1.077982, 1.101452, 
    1.092875, 0.7143764, -0.1856732, -0.347034, -0.1679814, 0.1676143, 
    0.1955928, -0.1845016, -0.1149052, -0.09359989, -0.6200159, -1.216142, 
    -0.8579714, -0.0185349, 0.3533564, 0.6741085, 0.9181027, 0.9629107, 
    1.011381, 0.9327186, 0.8927283, 0.8277544,
  0.6317742, 0.5717487, 0.2534552, 0.1535349, 0.0259161, -0.3818487, 
    -0.4754521, -0.1481084, 0.1536983, 0.2668657, 0.464229, 0.5506225, 
    0.06824875, -0.388538, -0.1540816, 0.3314327, 0.291589, 0.20238, 
    0.2198116, 0.1114131, 0.2229365, 0.285404, 0.2242711, 0.2737504, 
    0.3230338, 0.3199251, 0.4140823, 0.506319, 0.5085487, 0.1607943, 
    -0.702405, -0.747246, -0.5503218, -0.3049443, -0.1376591, 0.2614943, 
    0.6843138, 0.6418984, 0.119356, -0.3628221, 0.5918007, 1.782133, 
    1.607816, 1.301973, 1.055733, 0.7763708, 0.462878, 0.1284218, 
    -0.08331347, -0.03515291, -0.0261848, -0.3092899, -0.3985965, -0.2734338, 
    -0.04954052, 0.5163774, 0.7720253, 0.7841021, 0.7698277, 0.7107459, 
    0.8031611, 0.8562536, 0.7697139, 0.5880895, 0.4277217, 0.393721, 
    0.3724484, 0.38822, 0.4609737, 0.6747104, 0.8398311, 0.8025918, 
    0.9281125, 0.8855186, 0.7342, 0.5304718, -0.1155066, -0.06109655, 
    -0.04586226, -0.06396121, -0.2015426, -0.3714322, -0.2126753, 
    -0.08681279, -0.2475223, -0.9819462, -0.8464642, 0.4538119, 0.7149124, 
    0.8421749, 0.843249, 0.8137732, 0.8449416, 0.7126503, 0.6732621, 0.6017454,
  0.2947793, -0.01645088, -0.3460083, -0.3760695, -0.1846806, -0.187415, 
    -0.07691687, -0.01570275, 0.01974647, 0.2163123, 0.3929237, 0.2962111, 
    -0.04670861, -0.03126252, 0.1727089, 0.1958532, 0.1291866, 0.1820837, 
    0.2456744, 0.2666054, 0.2771195, 0.1757684, 0.1531122, 0.1604519, 
    0.1921582, 0.1555042, 0.1505899, 0.09611416, -0.1050577, -0.4668255, 
    -0.5924268, -0.4997525, -0.5835737, -0.2804652, 0.07147157, 0.3880246, 
    0.611413, 0.06315464, -0.1690392, 0.2039099, 1.139392, 1.471586, 
    1.090157, 0.7992716, 0.5091667, 0.1808138, -0.08647132, -0.179847, 
    -0.1860323, -0.1173301, -0.3537073, -0.5889124, -0.317672, 0.2120153, 
    0.6758336, 0.9843622, 0.9310419, 0.8984414, 0.9449905, 0.9809282, 
    0.9800656, 0.7624875, 0.5497106, 0.4866737, 0.4488808, 0.4860876, 
    0.3849971, 0.4537144, 0.5367875, 0.7024615, 0.7808137, 0.6416371, 
    0.8318396, 0.5838261, 0.4813843, 0.4565625, 0.1948276, 0.2687213, 
    -0.06360315, -0.1712693, -0.3403611, -0.1498659, 0.2057654, 0.1629105, 
    0.1517126, -0.4401008, -0.1582308, 0.9206903, 0.9057977, 0.8582882, 
    0.7982133, 0.8127154, 0.7319373, 0.5747595, 0.5525751, 0.3708529,
  0.05112696, -0.1440229, -0.1551394, -0.1342087, 0.1258501, 0.01014364, 
    -0.2644983, -0.1862106, 0.03076534, 0.2105668, 0.1675329, 0.08955455, 
    -0.0837692, -0.2129521, -0.03342748, 0.1786983, 0.1783892, 0.1035031, 
    0.01380551, 0.1440465, 0.1547563, 0.05322599, 0.05617189, -0.01295257, 
    0.006042004, 0.01437616, -0.07006454, -0.225256, -0.4211874, -0.7084265, 
    -0.7303829, -0.6573048, -0.6643683, -0.302096, -0.170797, 0.07194372, 
    -0.02100875, -0.4885218, -0.04145145, 0.4064652, 0.6311562, 0.6484413, 
    0.4198606, 0.07830715, -0.1035612, -0.05738592, -0.1626437, -0.08499002, 
    -0.10776, -0.2288048, -0.4864383, -0.3718063, 0.0867551, 0.5411821, 
    0.8875037, 0.8842973, 0.8717972, 0.9506872, 0.980619, 0.9101763, 
    0.7728064, 0.5903032, 0.4284216, 0.4298702, 0.3652381, 0.4275914, 
    0.3878782, 0.4858925, 0.5385942, 0.5487499, 0.5957878, 0.6241739, 
    0.6334672, 0.329659, 0.639473, 0.50142, 0.4243038, 0.1978878, -0.4136844, 
    -0.308688, 0.01663756, 0.219763, 0.2400427, 0.112878, 0.01458704, 
    -0.06609321, 0.5883169, 1.014115, 0.752852, 0.7606155, 0.6269403, 
    0.5521358, 0.4256222, 0.3880246, 0.29333, 0.1104202,
  -0.1625295, -0.246839, -0.1547492, -0.1755335, 0.009769253, -0.08761031, 
    -0.2904749, -0.3349897, -0.2414026, -0.1150029, -0.2846643, -0.1742148, 
    -0.1027633, -0.3490362, -0.2328088, 0.1746457, 0.1472857, -0.0409143, 
    -0.08499002, -0.06690741, -0.04455996, -0.08481097, -0.189873, 
    -0.1418097, -0.1554005, -0.1991827, -0.2613082, -0.4716272, -0.618258, 
    -0.6536751, -0.5612922, -0.3709763, -0.1307581, -0.06999946, -0.2901658, 
    -0.1398076, -0.4350877, -0.7071578, -0.2470666, 0.06183612, 0.5550494, 
    0.3659217, 0.1155963, 0.02137423, 0.01893258, -0.03479445, -0.5178348, 
    -0.3643193, -0.3147752, -0.5339157, -0.5639775, -0.2247522, 0.06183632, 
    0.2089717, 0.4741735, 0.5393591, 0.5914261, 0.6236526, 0.6449907, 
    0.6368851, 0.4595741, 0.3808467, 0.3098832, 0.335713, 0.2895873, 
    0.3417356, 0.3757362, 0.4190464, 0.4640007, 0.5394402, 0.533011, 
    0.532181, 0.4332399, 0.3845906, 0.4388871, 0.1330602, -0.163538, 
    0.008141756, -0.001184702, 0.2884802, 0.2126665, 0.09847379, 0.07684281, 
    0.097839, 0.01234087, 0.2773799, 0.9258987, 0.8763382, 0.608679, 
    0.5132846, 0.4036982, 0.3298216, 0.2229199, 0.1780469, 0.03602219, 
    -0.03381824,
  -0.1308718, -0.05666947, -0.04031205, -0.03280887, 0.01512408, -0.1292931, 
    -0.1247199, 0.01435912, 0.03532273, 0.01847696, -0.03787088, 0.2424679, 
    0.1439164, 0.005130649, 0.1613156, 0.2051796, 0.1897008, -0.1345341, 
    -0.3182906, -0.3090947, -0.233232, -0.1672325, -0.2158978, -0.2272098, 
    -0.2748008, -0.1303184, -0.2048953, -0.4151981, -0.5653284, -0.5173304, 
    -0.3126104, -0.1562301, -0.01788375, 0.02280635, -0.07717735, -0.1426067, 
    -0.3978152, -0.3143193, -0.03627563, 0.003519297, 0.2741898, -0.1877568, 
    -0.07050383, 0.04461622, -0.2567998, -0.2673305, -0.4497034, -0.05167282, 
    -0.08157189, -0.3042281, -0.003772378, 0.1324256, 0.09409541, 0.3505245, 
    0.6613969, 0.6952835, 0.6537797, 0.615303, 0.4867224, 0.4141314, 
    0.3892287, 0.4778683, 0.4559118, 0.3963416, 0.4032264, 0.3903847, 
    0.4027214, 0.4810586, 0.458483, 0.4663117, 0.3732944, 0.3942742, 
    0.3065789, 0.2720571, 0.1161661, -0.07595666, 0.1296749, 0.07816118, 
    0.1821976, 0.205212, 0.07104856, 0.1168493, 0.09531613, 0.03260455, 
    -0.1060348, 0.154919, 0.5156939, 0.5034705, 0.3799839, 0.1838738, 
    0.1867063, 0.09015679, 0.05739307, 0.04302144, -0.03961205, -0.0730114,
  -0.1988569, -0.1638637, -0.1368941, 0.02243209, 0.03128618, -0.1127892, 
    -0.01038039, 0.08494818, 0.07016963, 0.05703497, 0.2385453, 0.7725295, 
    0.2995153, -0.09934533, -0.1161911, -0.2617313, 0.07259479, -0.06518191, 
    -0.3098271, -0.09464157, -0.03666627, -0.04229772, 0.0002638102, 
    -0.2170048, -0.2530077, 0.05775082, -0.1843551, -0.3173628, -0.2423791, 
    -0.349264, -0.2565393, -0.04871053, -0.163538, -0.4773889, -0.4396774, 
    -0.1155889, 0.0344764, 0.1534542, 0.1369665, -0.05930627, -0.3985317, 
    -0.4388311, -0.1984176, -0.1901006, -0.3319137, 0.03473672, 0.2746294, 
    0.5499873, 0.2675493, 0.02148807, 0.3053582, 0.2204139, 0.2205275, 
    0.679512, 0.8591506, 0.823913, 0.7500688, 0.7052445, 0.636462, 0.5585974, 
    0.4771846, 0.3921585, 0.3870969, 0.375264, 0.3744988, 0.4380245, 
    0.4598017, 0.4723182, 0.359916, 0.309623, 0.2640982, 0.199271, 
    0.07221937, -0.04845047, -0.1301396, 0.01997432, 0.01894894, 0.1270381, 
    0.09020545, 0.05975297, 0.182279, 0.09458372, -0.0168258, 0.004219115, 
    -0.05756474, -0.2385867, -0.05845982, 0.2548864, 0.1816932, 0.06743532, 
    0.04655313, -0.1172327, -0.1077278, -0.1155239, -0.1706021, -0.1662235,
  -0.3178675, -0.2987431, -0.2258428, -0.02084601, 0.01554725, -0.04623661, 
    -0.08637334, -0.09695275, -0.07602177, 0.00402379, 0.1509477, 0.7727087, 
    1.036674, 0.8781281, 0.5154495, 0.1510941, 0.07106477, -0.07720992, 
    -0.2457321, -0.111178, -0.06524703, -0.08982387, -0.1112431, -0.1847783, 
    -0.04989871, 0.003844768, -0.1614059, -0.07802372, -0.1127567, 
    -0.2235481, -0.1220993, -0.1154423, -0.1144658, -0.6161909, -0.580823, 
    -0.02382451, 0.01953489, -0.08246708, -0.1355106, -0.5135868, -0.7115197, 
    -0.4651006, -0.6176398, -0.7691694, -0.6336713, -0.3710251, -0.3191047, 
    -0.2906866, -0.3780077, -0.4648564, -0.4163537, -0.4415491, -0.4461552, 
    -0.2601688, -0.1537724, -0.02567983, 0.07990271, 0.06906301, 0.06123406, 
    -0.01345667, -0.08671513, -0.1859176, -0.2257614, -0.1848921, -0.1833135, 
    -0.1748337, -0.190719, -0.1814417, -0.1188604, -0.08196247, -0.0930953, 
    -0.1631639, -0.1142864, -0.1370084, -0.3201298, -0.1671188, 0.08621782, 
    0.2523962, 0.1279984, 0.1291052, 0.08437863, -0.1347457, -0.2230432, 
    -0.2981408, -0.1722455, -0.4903774, -0.3796514, -0.103691, -0.1111129, 
    -0.06817675, -0.148564, -0.1795211, -0.1759403, -0.2973759, -0.3551723, 
    -0.3153934,
  -0.006246567, -0.03655231, -0.1120243, -0.005953401, 0.002575237, 
    0.04025428, 0.01956743, 0.1037634, 0.2816442, 0.1077836, 0.1093949, 
    0.3320512, 0.7266798, 1.293348, 1.272351, 1.050443, 0.5309607, 0.1622106, 
    0.03906614, 0.06364298, 0.2080604, 0.203796, 0.02125996, -0.1057909, 
    -0.02161092, 0.07622433, 0.2147499, 0.06849319, -0.143404, -0.3463836, 
    -0.03324819, -0.001754194, -0.0251103, -0.2803836, -0.5890589, 
    -0.4229295, -0.1254685, -0.1455692, -0.2897748, -0.3841599, -0.4989058, 
    -0.5186163, -0.7579715, -0.9710249, -1.087838, -1.015784, -1.137854, 
    -1.3554, -1.245113, -1.086666, -1.068925, -1.111797, -1.190247, -1.12402, 
    -0.97887, -1.049134, -1.133151, -1.139205, -1.110071, -1.10055, 
    -1.025973, -0.8918422, -0.8701625, -0.8498662, -0.7284307, -0.618665, 
    -0.4585576, -0.3335252, -0.2449508, -0.1835575, -0.1471155, -0.1387008, 
    -0.1062952, 0.1041378, 0.2547076, 0.126615, 0.4076209, 0.6394731, 
    0.346374, 0.2708044, 0.03081441, -0.1124966, -0.2048794, -0.161356, 
    -0.2315722, -0.388522, -0.3284632, -0.3033004, -0.3075647, -0.2489059, 
    -0.284111, -0.2279098, -0.2554163, -0.17804, -0.08870125, -0.01464462,
  0.06265011, -0.04298141, 0.01740271, -0.0109176, 0.02313161, 0.2549353, 
    0.3423537, 0.3429561, 0.2215204, 0.0523311, 0.1965043, 0.4554887, 
    0.7542353, 1.312, 1.164734, 1.297335, 1.283093, 0.8791864, 0.7108923, 
    0.9652706, 1.029398, 0.7681677, 0.5777705, 0.3110874, 0.1360059, 
    0.1854362, 0.1526079, 0.3164099, 0.9809446, 0.02336025, -0.08407784, 
    -0.1645962, -0.1138475, -0.1086551, -0.7617151, -0.7619594, -0.1686815, 
    0.01364279, -0.2812302, -0.2698693, -0.1109014, -0.07815385, -0.2195275, 
    -0.3292935, -0.5206993, -0.5165007, -0.6516564, -0.9760215, -1.151477, 
    -1.231181, -1.302893, -1.357402, -1.354961, -1.412529, -1.436308, 
    -1.548059, -1.642509, -1.72096, -1.832597, -1.774296, -1.681344, 
    -1.492281, -1.187366, -0.90693, -0.6956344, -0.6060836, -0.5433069, 
    -0.4609013, -0.2670374, -0.1368291, -0.08069283, 0.0594275, -0.06060791, 
    -0.01493776, 0.5738482, 0.1083695, -0.01026654, 0.345674, 0.3643916, 
    -0.1054327, -0.1404099, -0.06265926, 0.3107944, 0.1649446, -0.03162098, 
    -0.1271782, -0.07729125, -0.01845336, 0.00570035, -0.03853822, 
    -0.03046513, -0.05188429, -0.1161097, 0.07501991, 0.07960975, 0.08612016,
  0.2324417, -0.01083636, -0.2426558, -0.2598269, -0.3667443, -0.2388312, 
    0.0515337, 0.0823276, 0.2181349, 0.2838904, 0.2024613, 0.4282426, 
    0.6172073, 0.8835645, 0.8074589, 0.9666877, 1.255945, 0.9543819, 
    0.6877639, 0.9122432, 0.9397497, 0.7459669, 0.699271, 0.5756218, 
    0.2433953, 0.01431036, 0.1474485, 0.6007524, 1.587667, 0.6738, 0.2975297, 
    0.1006069, -0.06262589, 0.009866953, -0.6008101, -0.6796999, -0.4230924, 
    -0.1614549, -0.1246872, -0.2178347, 0.003795624, 0.152575, -0.0876267, 
    -0.1614063, -0.1894987, -0.1874151, -0.0861783, -0.1194139, -0.1749482, 
    -0.1795378, -0.2137175, -0.25138, -0.1282353, -0.1282024, -0.1555142, 
    -0.127861, -0.2271938, -0.2865849, -0.393291, -0.4792285, -0.4732227, 
    -0.4792936, -0.5761361, -0.557337, -0.5287564, -0.4460739, -0.4821578, 
    -0.4412235, -0.2580369, -0.1851529, -0.04636693, 0.4133828, 0.7528844, 
    0.1397343, -0.04399049, -0.1347296, -0.4002408, -0.3737917, -0.3617318, 
    -0.1866498, 0.1092644, 0.2265332, 0.1711457, 0.1241405, 0.003225803, 
    -0.03233719, -0.02026033, 0.08076501, 0.2254591, 0.306823, 0.3314974, 
    0.3411984, 0.3338578, 0.3370155, 0.325036, 0.284476,
  0.1659539, 0.09477901, -0.1076133, -0.2334929, -0.3223109, -0.5346808, 
    -0.463099, -0.3634562, -0.3034468, -0.3159623, -0.1811163, 0.06037146, 
    0.1205928, 0.2635125, 0.6218629, 0.4714403, 0.6048222, 0.7316775, 
    0.6272981, 0.4679563, 0.4429885, 0.8002317, 1.076323, 0.9743197, 
    0.5591183, 0.1853218, 0.3411167, 0.3490925, 0.7242382, 0.6462603, 
    0.7797737, 0.6085982, 0.2471557, 0.1423697, -0.03492522, -0.127666, 
    -0.2095344, 0.03496408, 0.0561235, -0.06113005, 0.09539771, 0.2587268, 
    0.2035184, 0.1293001, 0.1103873, -0.07509446, -0.1500945, -0.1726041, 
    -0.1057093, 0.02801442, 0.07485676, 0.02733064, 0.08449221, 0.1744823, 
    0.1733761, 0.2657583, 0.3341508, 0.4515171, 0.4073286, 0.157393, 
    -0.06052637, -0.195569, -0.3391886, -0.3758588, -0.4151335, -0.411113, 
    -0.5224082, -0.6005663, -0.4430791, -0.1690722, 0.1564653, 0.2882845, 
    0.548522, 0.04863644, -0.3310351, -0.1416302, -0.06568646, 0.05063856, 
    0.2809768, 0.7681842, 0.8352895, 0.5049679, 0.2591994, 0.1498568, 
    0.06146169, -0.02992845, -0.05847645, 0.01461935, 0.05902052, 0.1582718, 
    0.2713909, 0.3988485, 0.2586788, 0.2519729, 0.2628943, 0.2059443,
  0.2599807, 0.05793047, -0.03795195, -0.01015234, -0.01848578, -0.3056445, 
    -0.5383425, -0.3261685, -0.2392049, -0.3048625, -0.4532351, -0.1211552, 
    0.003974978, -0.05019164, 0.2578321, 0.3351927, 0.354301, 0.4003301, 
    0.3907104, 0.1864128, 0.05832082, 0.3779008, 0.7543492, 0.8863964, 
    0.5469276, -0.009566694, 0.105749, 0.1288774, 0.456579, 1.148654, 
    1.073442, 0.7984586, 0.7984576, 0.6053753, 0.2844934, 0.06247067, 
    -0.1654751, 0.07353783, 0.1993527, 0.03859425, 0.09388399, 0.2667356, 
    0.2869987, 0.1268101, 0.1597846, -0.01231766, -0.1836555, -0.2554984, 
    -0.2885382, -0.1597948, 0.05111003, 0.1806998, 0.2634306, 0.344502, 
    0.2685575, 0.3593941, 0.5685253, 0.6131706, 0.4478223, 0.382165, 
    0.2641635, 0.1743855, 0.0549202, -0.1582799, -0.2381139, -0.2917442, 
    -0.5236945, -0.7180465, -0.4627566, -0.1396611, -0.08975863, -0.1441698, 
    -0.1709763, -0.3887501, -0.0410769, 0.434818, 0.5539261, 0.7192745, 
    0.8315954, 0.7460648, 0.4218134, 0.3039098, 0.2117875, -0.02195263, 
    -0.1858523, -0.2998495, -0.3263965, -0.197067, -0.02465487, 0.09552765, 
    0.1038451, 0.2515988, 0.2271197, 0.3156123, 0.4779491, 0.4760287,
  0.8490922, 0.4046749, -0.2168581, -0.3485644, -0.1847785, -0.3354455, 
    -0.6375778, -0.4716437, -0.2242308, -0.1473269, -0.2323041, -0.0940721, 
    -0.06088504, -0.3110151, -0.08186507, 0.215287, 0.1213744, 0.08304358, 
    0.4090207, 0.3493204, -0.1066859, -0.1927046, -0.09566694, 0.2293494, 
    0.3744664, -0.06345665, 0.04287472, 0.1927933, 0.1928258, 0.6140509, 
    0.8727422, 0.8245487, 0.8262572, 0.7779016, 0.4185424, 0.2765985, 
    0.00543952, -0.07585931, 0.2112014, 0.08516002, -0.08010697, 0.1324742, 
    0.206286, 0.1456091, 0.2098017, 0.09559298, -0.03415942, -0.2239871, 
    -0.3526328, -0.2902145, -0.1219852, 0.02604532, 0.1366081, 0.3852575, 
    0.5665562, 0.6637896, 0.7074255, 0.8248897, 0.785615, 0.6857128, 
    0.5338907, 0.4184604, 0.2956262, 0.06234169, -0.006326675, -0.0538373, 
    -0.1416945, -0.3088021, -0.09993136, -0.03113246, 0.008483291, 0.2080929, 
    -0.2154751, -0.5848759, -0.1168259, 0.3226599, 0.5926142, 0.8600134, 
    0.935176, 0.8563023, 0.6933954, 0.4602575, 0.1169796, -0.1166632, 
    -0.3085738, -0.3679324, -0.4009895, -0.3548141, -0.1066692, 0.05884123, 
    0.1364129, 0.3004103, 0.4101111, 0.4684608, 0.5155146, 0.7737663,
  0.5392449, 0.6779332, 0.2067094, -0.1886034, -0.2448372, -0.4626429, 
    -0.7260541, -0.7594361, -0.5199511, -0.2755823, -0.2268353, -0.1801395, 
    -0.2545374, -0.3457483, -0.07655907, 0.1064975, 0.03965187, 0.04136109, 
    0.08862686, 0.1140983, -0.0202601, -0.07712877, 0.1346879, 0.1397336, 
    -0.0465133, -0.1630172, -0.06267554, 0.06577516, 0.1748573, 0.2308137, 
    0.3946981, 0.4543333, 0.2976766, 0.5175824, 0.3166385, 0.3334508, 
    0.3428907, 0.1121941, 0.2579629, 0.2761918, 0.03408563, -0.008150697, 
    -0.04148424, -0.04877591, -0.04163063, -0.09233046, -0.09412098, 
    -0.2559211, -0.3586714, -0.4608849, -0.3253056, -0.05745077, -0.0349735, 
    0.05010128, 0.3509476, 0.7458043, 0.8875035, 0.8841507, 0.7709669, 
    0.632686, 0.5462925, 0.4555211, 0.4009151, 0.2731977, 0.0443244, 
    -0.08881426, 0.03314209, 0.08200216, 0.07405961, 0.1429399, 0.2455276, 
    0.136755, -0.4369105, -0.385055, -0.1387824, 0.03963578, 0.4365922, 
    0.7395707, 0.9595252, 0.8558956, 0.5734572, 0.2757848, -0.06874657, 
    -0.3227175, -0.763473, -1.026559, -0.9318973, -0.5708947, -0.1928023, 
    -0.02319002, 0.2109413, 0.3104851, 0.3364948, 0.4252477, 0.2269894, 
    0.2031116,
  0.2090044, 0.3770057, 0.3340695, 0.08924517, -0.02323854, -0.2558557, 
    -0.6421025, -0.877991, -0.6984988, -0.2846805, -0.1663212, -0.07999311, 
    -0.1571251, -0.214775, 0.04137731, 0.04279333, -0.04161441, -0.1337694, 
    -0.1026819, 0.3647008, 0.4594595, -0.04084945, -0.07953739, -0.2949183, 
    -0.4159472, -0.1506149, 0.1874224, -0.270895, -0.3182092, 0.08854485, 
    0.277705, 0.3985877, 0.4157758, 0.5532598, 0.5849652, 0.5293658, 
    0.5786166, 0.4922559, 0.3755568, 0.3640174, 0.3293816, 0.2124711, 
    0.1305539, 0.1087277, 0.06362671, 0.05176145, 0.009948194, -0.06506807, 
    -0.1504684, -0.4663701, -0.5861617, -0.4353805, -0.2631311, 0.02342492, 
    0.3199254, 0.7586786, 1.037146, 0.9921424, 0.9701045, 0.889652, 
    0.6649938, 0.3705442, 0.1684761, 0.02409267, -0.07414913, -0.09275246, 
    -0.08267856, -0.0423629, -0.0278284, 0.04305375, 0.2253129, -0.08455086, 
    -0.5515914, -0.29845, -0.03210896, 0.1787797, 0.4712439, 0.5114294, 
    0.8180537, 0.8696001, 0.6890011, 0.4616573, -0.09189092, -0.5990524, 
    -1.10553, -1.527812, -1.580937, -1.075322, -0.4068322, 0.003502972, 
    0.3362342, 0.3781772, 0.4523309, 0.5348831, 0.3921098, 0.2356644,
  0.7749873, 0.6078324, 0.2403846, -0.08625939, -0.2717575, -0.5472132, 
    -0.7274216, -1.03372, -1.064303, -0.3731083, -0.1553674, -0.1274378, 
    -0.1002731, 0.004088912, 0.1990434, 0.1266312, 0.08376023, 0.01331744, 
    -0.2196253, -0.1217899, -0.006246328, -0.5270149, -1.023287, -0.976624, 
    -0.9882946, -1.045602, -0.5784473, -0.4743781, -0.3185349, 0.06103873, 
    0.1555049, 0.09458351, 0.3041053, 0.4185748, 0.6940956, 0.7769899, 
    0.6683304, 0.767956, 0.6561556, 0.4294468, 0.2808143, 0.128975, 
    0.01266638, -0.07073206, -0.07322228, 0.06929082, 0.1331579, 0.1806026, 
    0.2906123, 0.1654497, -0.09656203, -0.3024377, -0.3276007, -0.1641402, 
    0.05355191, 0.5664427, 0.964587, 0.9996943, 1.03018, 0.942777, 0.6921911, 
    0.4253778, 0.08304429, -0.1181288, -0.0683887, -0.01324522, -0.1345015, 
    -0.1618291, -0.1859502, 0.0105505, 0.2722693, 0.1758826, 0.02788448, 
    0.1343135, 0.09993853, 0.3486039, 0.6415564, 0.6134641, 0.6360716, 
    0.533337, 0.3524937, 0.1494828, -0.237301, -0.6249963, -1.231881, 
    -1.902812, -2.13595, -1.735511, -0.96943, -0.2730597, 0.3779823, 
    0.6181352, 0.5813675, 0.5684443, 0.3823115, 0.5463253,
  0.5530472, 0.7512569, 0.4387568, 0.05299842, -0.2194137, -0.493372, 
    -0.7945602, -1.034941, -1.042103, -0.7352666, -0.3753544, -0.2265752, 
    0.02622432, 0.1335646, 0.09847343, 0.09412777, 0.3131711, 0.5131872, 
    0.1957231, -0.2592249, -0.2527144, -0.02540302, -0.2081342, -0.1475549, 
    -0.1469039, -0.5929167, -0.4825974, -0.09897098, -0.1003056, 0.01751667, 
    0.05771852, -0.1324673, 0.07750964, -0.005497456, 0.2440629, 0.2774284, 
    0.02990282, 0.02347368, 0.3496289, 0.3501987, 0.186169, 0.01471722, 
    -0.1504033, -0.3608363, -0.4928839, -0.4114224, -0.2648889, -0.14609, 
    0.02440155, 0.1388545, 0.1381874, 0.1018753, 0.06784248, -0.03512096, 
    0.02026701, 0.4846389, 0.9699578, 1.094079, 1.044698, 0.9755247, 
    0.8149937, 0.4494502, -0.09005165, -0.3713508, -0.3443973, -0.3120733, 
    -0.368144, -0.2817346, -0.4080531, -0.5085414, -0.3253381, -0.01721638, 
    0.1967158, 0.252396, 0.1535031, 0.2882523, 0.7703486, 1.228129, 1.253357, 
    0.9574091, 0.6344601, 0.1484249, -0.3771447, -0.7606897, -1.302128, 
    -1.964596, -2.342689, -2.196122, -1.65872, -0.885576, 0.03115511, 0.5821, 
    0.7083371, 0.5943558, 0.3949418, 0.2961137,
  0.3126989, 0.8850784, 0.5901241, 0.1090531, -0.02608681, -0.2403446, 
    -0.5979457, -0.519544, -0.5242802, -0.6696091, -0.7995895, -0.3887169, 
    -0.01010406, 0.04046589, -0.06418908, -0.04431593, 0.03229541, 0.4113806, 
    0.6810911, 0.5097532, -0.01482368, -0.01773727, 0.0745967, -0.128691, 
    -0.1902306, -0.3419885, -0.3139775, -0.05828089, 0.007734746, 0.09188187, 
    0.1728387, 0.1765012, 0.2349315, -0.01796532, -0.03593421, 0.1752644, 
    0.001386642, -0.2109827, -0.3104455, -0.1442351, -0.02374339, 
    -0.09039342, -0.2809533, -0.4852015, -0.6491174, -0.7392868, -0.7658491, 
    -0.7526002, -0.6651657, -0.4837697, -0.2818489, -0.07348299, 0.05470657, 
    0.02947927, -0.06685877, 0.02134275, 0.3359904, 0.7219119, 0.9456904, 
    0.8016317, 0.4602089, 0.2531611, -0.01744449, -0.309827, -0.4437302, 
    -0.6767542, -0.6223922, -0.4484175, -0.5052859, -0.7470993, -0.8024704, 
    -0.4860153, -0.1500614, 0.2082231, 0.4622273, 0.4449253, 0.5020218, 
    0.8493363, 1.135469, 1.140254, 1.032539, 0.6670769, 0.04642296, 
    -0.5527469, -1.10444, -1.595944, -2.052161, -2.218828, -1.92223, 
    -1.342395, -0.567493, 0.1916864, 0.7185423, 0.7161496, 0.2493688, 
    -0.01648402,
  0.4544633, 0.7511432, 0.419958, -0.1570276, -0.3683882, -0.3241988, 
    -0.6692672, -0.6765426, -0.3794397, -0.3113736, -0.247197, -0.1501267, 
    -0.3402959, -0.3378219, -0.3593063, -0.01786757, 0.24071, 0.3235062, 
    0.4719924, 0.3476274, -0.2362597, -0.189661, 0.01689816, -0.08591759, 
    -0.253154, -0.2087692, -0.1221155, -0.02647749, -0.04276982, -0.05362593, 
    0.0276078, 0.2567908, 0.3295609, 0.1379917, -0.1176071, 0.05963826, 
    0.3308153, 0.1457391, -0.2678024, -0.5971968, -0.5959276, -0.497734, 
    -0.4834598, -0.5462854, -0.5958948, -0.6431768, -0.7333624, -0.8126426, 
    -0.7975554, -0.7316372, -0.6890762, -0.5023079, -0.2188282, 0.001045227, 
    0.1312704, 0.2033405, 0.1290565, 0.2320514, 0.5377645, 0.6268759, 
    0.3546259, 0.1835971, 0.01167321, -0.2580371, -0.2585416, -0.2176883, 
    -0.4573369, -0.6384078, -0.568909, -0.7153937, -0.7793745, -0.7045049, 
    -0.444495, 0.002705574, 0.5926144, 0.7307004, 0.7060745, 0.8123246, 
    1.001517, 0.9605831, 0.8583207, 0.7159703, 0.4411495, -0.07248974, 
    -0.6867639, -1.133199, -1.426022, -1.557255, -1.437366, -1.14513, 
    -0.7077923, -0.1017213, 0.4222374, 0.5615597, 0.3854201, 0.2215858,
  0.4110715, 0.3755243, 0.2383988, -0.02571252, -0.1032353, -0.1127243, 
    -0.4106084, -0.6956995, -0.6933558, -0.4616499, -0.2062302, -0.1006801, 
    -0.3076786, -0.5859014, -0.657353, -0.2361621, 0.3041377, 0.4823442, 
    0.4923866, 0.3915724, 0.1520219, 0.02480841, 0.0622108, 0.009183049, 
    -0.08798466, -0.04506475, 0.03532263, 0.1368526, 0.04103565, -0.1602503, 
    -0.1729782, -0.03206038, 0.06855834, -0.04250944, -0.1957483, -0.2508265, 
    -0.1375453, 0.1079144, -0.009370804, -0.3826947, -0.7100551, -0.7247683, 
    -0.5770633, -0.5606898, -0.5921676, -0.5827925, -0.6150193, -0.5956508, 
    -0.3356895, -0.1838667, -0.3217409, -0.4003386, -0.2169564, -0.01567078, 
    0.2207394, 0.5538454, 0.6360726, 0.4583702, 0.3982453, 0.3918333, 
    0.2185097, 0.03008318, -0.09451151, -0.1815233, 0.0635612, 0.05703425, 
    -0.2828093, -0.5110804, -0.481458, -0.5548467, -0.5929489, -0.5393682, 
    -0.4946904, -0.3623824, 0.041475, 0.3420935, 0.563285, 0.6932818, 
    0.7485225, 1.003959, 1.178275, 0.9306189, 0.5144733, 0.1994828, 
    -0.1229779, -0.5642867, -1.075078, -1.390638, -1.298174, -0.9253864, 
    -0.5149698, -0.05110264, 0.3354697, 0.441915, 0.5341668, 0.4857616,
  0.6677284, 0.461072, 0.2996941, 0.02187848, -0.06793249, -0.06750965, 
    -0.1575649, -0.4523889, -0.6339808, -0.655449, -0.4393842, -0.1693323, 
    -0.1748827, -0.3673146, -0.4087369, -0.1506634, 0.04901099, 0.1295123, 
    0.2266963, 0.3856968, 0.3534702, 0.1843626, 0.04359198, -0.2543914, 
    0.01011086, -0.1912723, -0.1768521, -0.05627893, -0.009940982, 
    0.02838907, 0.1137407, 0.09040046, 0.04215837, -0.05779278, -0.1128383, 
    -0.1539677, -0.1292119, -0.01472628, 0.2625537, 0.1254926, -0.2111456, 
    -0.3658328, -0.2615523, -0.204082, -0.2661583, -0.398027, -0.5929815, 
    -0.5727503, -0.1044398, 0.3653357, 0.3740597, 0.1598343, 0.1084023, 
    0.116703, 0.1962278, 0.5483427, 0.9391632, 0.9865441, 0.7045774, 
    0.3201699, 0.008419037, -0.1132774, -0.124362, -0.0910449, -0.2084601, 
    -0.1974573, -0.2494432, -0.2417769, -0.3289514, -0.4856409, -0.5034469, 
    -0.430807, -0.4108363, -0.2870894, -0.06970668, 0.2709184, 0.5296425, 
    0.6044958, 0.6459835, 0.8608924, 1.414733, 1.049499, 0.8284216, 
    0.4901728, 0.3043005, 0.05239618, -0.3266401, -0.622148, -0.7052534, 
    -0.7070277, -0.5906706, -0.1923461, 0.2349, 0.4253621, 0.5780957, 
    0.7480989,
  0.7211137, 0.6418169, 0.3890011, 0.2644899, 0.1509316, 0.01772797, 
    -0.2118777, -0.5115685, -0.6467899, -0.730579, -0.7166306, -0.4283003, 
    -0.2633426, -0.370944, -0.316761, -0.1241663, -0.02144837, 0.0004920959, 
    0.0008985996, 0.05482149, 0.1080117, 0.08257174, 0.07446671, 0.2145543, 
    0.2318234, 0.06642628, -0.06330991, -0.07076454, -0.06373322, 
    -0.01951134, 0.07562214, 0.1600456, 0.1149452, 0.07300162, -0.01352215, 
    -0.007353306, 0.02436876, -0.04700184, -0.2711058, -0.3490515, 
    -0.4320929, -0.1808071, 0.01712584, 0.3308301, 0.1823275, -0.09788036, 
    -0.316191, -0.2257936, 0.2411981, 0.7583043, 0.8413284, 0.6168493, 
    0.5331254, 0.5690139, 0.6056191, 0.5906444, 0.6147656, 0.6614451, 
    0.6202512, 0.4541869, 0.2675986, 0.1169467, 0.15308, -0.1223433, 
    -0.1781538, -0.1108692, -0.1924932, -0.2845016, -0.3284306, -0.2154261, 
    -0.1590784, -0.1982711, -0.2786585, -0.1413863, 0.08286482, 0.3762406, 
    0.3349322, 0.4565953, 0.510941, 0.6918982, 0.9684607, 1.499124, 1.498376, 
    1.231351, 0.8936071, 0.5809281, 0.3600949, 0.2230017, 0.2150593, 
    0.1259966, 0.02737999, 0.07723331, 0.2501836, 0.3262897, 0.4032097, 
    0.6104856,
  0.6676309, 0.5775266, 0.5198278, 0.4299186, 0.4623408, 0.3355669, 
    0.05626965, -0.07209897, -0.1055304, -0.241012, -0.4030727, -0.3920046, 
    -0.2949178, -0.1734502, -0.1230435, -0.06599545, -0.06519818, -0.1297653, 
    -0.1536422, -0.1461711, -0.09540629, -0.01155233, 0.03952169, 0.04876614, 
    0.04253316, -0.06562114, -0.06659818, -0.1152632, -0.07068312, 
    -0.0716598, -0.04359972, -0.03074181, -0.009468913, 0.003014803, 
    -0.04926395, -0.0329392, 0.02366877, -0.102356, -0.4217091, -0.3414025, 
    -0.4898877, -0.3467417, -0.09862995, -0.1175747, 0.2376838, 0.1979051, 
    0.2178593, 0.4090853, 0.7598667, 1.185501, 1.344746, 1.180016, 0.9801468, 
    0.9884962, 1.017761, 1.130684, 0.9192584, 0.632865, 0.4255402, 0.3954456, 
    0.5348177, 0.3864126, 0.1902382, 0.08325577, 0.07656598, 0.1297238, 
    0.07345748, -0.01303339, -0.05414677, 0.004691124, -0.1014938, 
    -0.5853968, -0.9330369, -0.79596, -0.2971481, 0.1634476, 0.2003779, 
    0.3293331, 0.4403682, 0.6494013, 1.1022, 1.710778, 1.888479, 1.808907, 
    1.621211, 1.393379, 1.001648, 0.6391639, 0.5262895, 0.5680702, 0.5655799, 
    0.5365922, 0.5421913, 0.5734899, 0.640352, 0.6506062,
  0.945853, 0.9016154, 0.6849322, 0.5401728, 0.3906939, 0.2247595, 0.1016476, 
    0.1632361, 0.1165727, -0.01793253, -0.1849082, -0.2677044, -0.2100712, 
    -0.1631473, -0.1110803, -0.05118454, -0.07893538, -0.1065557, -0.1492476, 
    -0.09438086, 0.04370499, 0.07181382, 0.008418322, -0.04623699, 
    -0.01682615, -0.02349925, 0.03198612, 0.01920927, -0.02079713, 
    -0.06978798, -0.1227016, -0.1133915, -0.106344, -0.1612594, -0.2464156, 
    -0.2265752, -0.1998173, -0.1527309, -0.4115853, -0.5140581, -0.6941528, 
    -0.4631467, -0.4324179, -0.5160613, -0.5797648, -0.3505163, -0.3344035, 
    0.05563545, 0.3508182, 0.9116583, 1.357524, 1.36379, 0.8461947, 
    0.3595086, 0.2216506, 0.3530309, 0.4179561, 0.4158404, 0.2006711, 
    0.2135128, 0.2253451, 0.207116, 0.1957879, 0.1114947, 0.1350622, 
    0.2799515, 0.2904496, 0.1453162, -0.07602167, -0.3097945, -0.6772749, 
    -1.22708, -1.561341, -1.519121, -1.146041, -0.7127891, -0.6002893, 
    -0.6637496, -0.6961229, -0.30527, 0.7619011, 1.684834, 1.579186, 
    0.8966182, 0.8869828, 1.176436, 1.231563, 1.22751, 1.165238, 1.072399, 
    0.8810256, 0.6754267, 0.5549679, 0.5948931, 0.7788939, 0.9233437,
  0.9589717, 0.8712273, 0.7789094, 0.6614459, 0.5825558, 0.413106, 0.3851924, 
    0.3168166, 0.2581416, 0.1430048, 0.06426144, -0.03349221, -0.08572257, 
    -0.07297826, -0.04963827, -0.0491662, -0.07999301, -0.0908004, 
    -0.02966785, 0.09575558, 0.2354693, 0.2650917, 0.1518919, 0.03603888, 
    0.01546597, -0.06469381, -0.001965761, 0.01955104, -0.009110957, 
    -0.05515588, -0.09875941, -0.1353155, -0.2576136, -0.3547815, -0.3101201, 
    -0.2780074, -0.3490198, -0.3731084, -0.5395632, -0.6083626, -0.5945437, 
    -0.6766243, -0.7877243, -0.8575485, -0.8732874, -0.7940071, -0.7842083, 
    -0.5548134, -0.2240033, 0.09469843, 0.5249233, 0.2103076, 0.6723666, 
    0.3388058, 0.0755083, 0.009655297, 0.03154659, 0.07174841, 0.0890826, 
    0.1466997, 0.1265336, 0.1767941, 0.1805051, 0.1571162, 0.1471065, 
    0.2061885, 0.2185095, 0.05661166, -0.1690718, -0.3710901, -0.5407516, 
    -0.6556118, -0.7910281, -0.8888149, -0.9634567, -1.078723, -1.156653, 
    -1.306507, -1.034827, -0.4943972, 0.2529655, 0.8801138, 0.790482, 
    0.3829626, -0.08941686, -0.1553998, 0.2687535, 1.159802, 1.814474, 
    2.222513, 2.344306, 1.90264, 1.874694, 1.605603, 1.3446, 1.084867,
  1.577185, 1.126273, 0.7282099, 0.4183304, 0.2067742, 0.1571164, 0.1397338, 
    0.1643265, 0.1757849, 0.1823604, 0.2018431, 0.08359754, 0.08639693, 
    0.2378457, 0.1254916, 0.2669466, 0.2819374, 0.287699, 0.3134966, 
    0.3527707, 0.3598181, 0.3408403, 0.2703321, 0.2039258, 0.1289258, 
    0.04767632, 0.07921898, 0.1001014, 0.05778357, -0.0115198, -0.1110641, 
    -0.274329, -0.4042119, -0.3882937, -0.3236128, -0.204749, -0.1303512, 
    -0.1392705, -0.21554, -0.3224083, -0.369674, -0.3596158, -0.3263309, 
    -0.3061976, -0.2704554, -0.2487917, -0.2927048, -0.4042773, -0.5299277, 
    -0.5801063, -0.9154096, -0.8922977, -0.3516736, 0.2138546, 0.3046098, 
    0.3201696, 0.2942092, 0.2378291, 0.2599483, 0.1840694, 0.1898311, 
    0.202445, 0.1820186, 0.1100785, 0.03817099, 0.00729531, -0.07667285, 
    -0.2589482, -0.4154098, -0.5761031, -0.6280237, -0.6806115, -0.6076624, 
    -0.5646611, -0.4167607, -0.4664191, -0.5766401, -0.6923143, -0.5851853, 
    -0.5790656, -0.3005171, 0.2308142, 0.2530961, 0.07944679, -0.1129194, 
    -0.1876591, -0.1690071, 0.2986374, 0.9264531, 0.8839073, 0.4471722, 
    0.9394412, 1.847449, 2.316914, 2.348766, 2.039782,
  2.311689, 2.070414, 1.676192, 1.230586, 0.8615434, 0.6424679, 0.5686886, 
    0.6255406, 0.7465204, 0.8492223, 0.8722204, 0.7934443, 0.7904494, 
    0.7561883, 0.722074, 0.2837603, 0.3996619, 0.5402218, 0.6191118, 
    0.6102739, 0.5816441, 0.4943235, 0.4185905, 0.30181, 0.2119663, 
    0.1225786, 0.08166027, 0.04713917, 0.006090857, -0.06482385, -0.1245406, 
    -0.1547977, -0.1548954, -0.1190066, -0.07719362, -0.04063761, 0.01125038, 
    -0.02515914, -0.09480432, -0.1402145, -0.1437138, -0.1750453, -0.1758265, 
    -0.1488571, -0.07006472, 0.02126014, 0.1014198, 0.1525425, 0.1429563, 
    0.08724284, 0.06094074, 0.05867839, 0.1160684, 0.254463, 0.3422726, 
    0.3883338, 0.4167354, 0.3850785, 0.3470577, 0.3113806, 0.3010616, 
    0.3331254, 0.3028519, 0.1428746, 0.02043009, -0.1374313, -0.3140752, 
    -0.5215621, -0.7023727, -0.7693974, -0.9032028, -0.9061975, -0.9023075, 
    -0.7363409, -0.6689906, -0.528105, -0.5650194, -0.7970014, -0.8622525, 
    -0.829342, -0.479456, -0.02870727, 0.08576179, 0.3499055, 0.5451205, 
    0.4932981, 0.3711137, 0.2767129, 0.1116734, 0.03921366, 0.08304501, 
    0.2766156, 0.7540073, 0.9333041, 1.432767, 2.161234,
  1.333694, 1.652705, 1.874385, 1.811511, 1.624548, 1.332718, 1.188627, 
    1.066459, 1.120576, 1.13529, 1.184997, 1.129691, 0.9699093, 0.7384639, 
    0.5246944, 0.4017452, 0.3939326, 0.4436071, 0.4998734, 0.5437861, 
    0.5689977, 0.534867, 0.46641, 0.3224809, 0.1681514, 0.09212601, 
    -0.04862916, -0.1689255, -0.2647588, -0.3132776, -0.3830041, -0.3519983, 
    -0.3314091, -0.273564, -0.2202437, -0.2078252, -0.1968388, -0.1794723, 
    -0.1645309, -0.1659469, -0.1863408, -0.2239222, -0.2671351, -0.3000126, 
    -0.2796513, -0.2038864, -0.09582949, 0.03699923, 0.1597854, 0.2570835, 
    0.3041376, 0.3134311, 0.313952, 0.3300653, 0.3549514, 0.382881, 
    0.4049677, 0.4202509, 0.4183465, 0.4017614, 0.3498409, 0.2912797, 
    0.2425492, 0.2128129, 0.1500687, -0.009989865, -0.1318486, -0.2588994, 
    -0.3955531, -0.511943, -0.6011031, -0.6327438, -0.6395797, -0.4922002, 
    -0.4303512, -0.4922491, -0.4118454, -0.5584275, -0.2040166, -0.09259078, 
    -0.07042277, 0.05320954, 0.2451048, 0.4050977, 0.4960163, 0.526631, 
    0.5054235, 0.3918983, 0.2439492, 0.1427441, 0.1410518, 0.2879276, 
    0.4900913, 0.7011263, 0.9766145, 1.235924,
  0.7223018, 0.8676795, 1.02808, 1.013171, 0.9922887, 0.9793167, 0.9869664, 
    0.8398799, 0.8528683, 0.8501014, 0.8154985, 0.7751502, 0.7559932, 
    0.7372921, 0.7179072, 0.6912308, 0.6693395, 0.6671423, 0.6676793, 
    0.6534541, 0.635404, 0.6205928, 0.5626175, 0.467663, 0.3793004, 0.283272, 
    0.1557817, 0.0924027, -0.02891886, -0.1428186, -0.2538701, -0.3240849, 
    -0.3711389, -0.4025353, -0.4192671, -0.4130009, -0.4001265, -0.3891728, 
    -0.3699671, -0.3458134, -0.3346643, -0.3266891, -0.323499, -0.3272262, 
    -0.3328577, -0.3323858, -0.3110479, -0.2801234, -0.2363083, -0.1757288, 
    -0.1156377, -0.03889608, 0.04316771, 0.117712, 0.1940303, 0.2467158, 
    0.286755, 0.2920771, 0.2732946, 0.2496293, 0.2228552, 0.1901566, 
    0.155212, 0.1200719, 0.08315778, 0.02967489, -0.05040336, -0.1392704, 
    -0.2469365, -0.3341272, -0.4102503, -0.4037724, -0.4661259, -0.507174, 
    -0.4782028, -0.4931442, -0.4435513, -0.3342575, -0.2382774, -0.1049936, 
    0.05788088, 0.1305859, 0.2093132, 0.2317586, 0.2870151, 0.3442254, 
    0.3669145, 0.3152216, 0.2093297, 0.09183335, 0.03994536, 0.1190794, 
    0.1328487, 0.3080931, 0.4540079, 0.5966182,
  0.2599481, 0.3568557, 0.4674026, 0.5604364, 0.63376, 0.7047073, 0.7566116, 
    0.784167, 0.792712, 0.7748735, 0.7454627, 0.7175655, 0.687113, 0.6645056, 
    0.6385942, 0.6143103, 0.6045283, 0.6119665, 0.611706, 0.6035192, 
    0.6033238, 0.5987829, 0.5787796, 0.5620804, 0.5451859, 0.5169306, 
    0.4710322, 0.4184443, 0.3195023, 0.2309607, 0.1466833, 0.05799514, 
    -0.03241825, -0.1118941, -0.1835413, -0.2492315, -0.3127242, -0.3530725, 
    -0.3814742, -0.3972294, -0.4010217, -0.3887333, -0.3616826, -0.338652, 
    -0.3189254, -0.3031865, -0.2862431, -0.2793746, -0.2746546, -0.268665, 
    -0.2449672, -0.2120082, -0.1806767, -0.1575159, -0.1328089, -0.1071579, 
    -0.0817672, -0.04872686, -0.01568645, 0.008320689, 0.03465533, 
    0.05674189, 0.0741573, 0.08515978, 0.08255571, 0.0767777, 0.06317097, 
    0.03776407, -0.003918886, -0.06741175, -0.1282516, -0.1759892, 
    -0.2224898, -0.2339156, -0.1695765, -0.1871548, -0.1631477, -0.1212043, 
    -0.08988917, -0.05043602, 0.01899779, 0.008499861, 0.02778697, 
    0.02663136, 0.01645875, -0.03975874, -0.08415979, -0.1161259, -0.1727178, 
    -0.199785, -0.1851525, -0.1414514, -0.09394169, -0.01954389, 0.0739944, 
    0.1670933,
  0.2479204, 0.2850786, 0.3254918, 0.3639684, 0.394307, 0.4253128, 0.4567907, 
    0.4799516, 0.4913936, 0.5076859, 0.5146846, 0.5128617, 0.5154984, 
    0.527445, 0.53057, 0.5256058, 0.5226111, 0.5245479, 0.5133826, 0.4991247, 
    0.4925492, 0.479805, 0.4710647, 0.4526403, 0.4344925, 0.4124385, 
    0.3840368, 0.3542678, 0.3189651, 0.2819372, 0.24696, 0.2038773, 
    0.1659704, 0.1214718, 0.08216512, 0.03765011, -0.005904555, -0.0510543, 
    -0.08510381, -0.1171675, -0.1466435, -0.1743127, -0.1952437, -0.2234989, 
    -0.2514775, -0.2738896, -0.2883753, -0.3027308, -0.3130172, -0.3226852, 
    -0.3319463, -0.3351038, -0.3393356, -0.342428, -0.3351201, -0.328333, 
    -0.3206344, -0.3117477, -0.299443, -0.2824671, -0.2703252, -0.2610316, 
    -0.2506312, -0.2439906, -0.2425258, -0.2356897, -0.2218877, -0.2112106, 
    -0.2166142, -0.2179163, -0.2233688, -0.22415, -0.2375289, -0.2418095, 
    -0.2491989, -0.2560185, -0.2564905, -0.2548304, -0.2513473, -0.2468714, 
    -0.2387171, -0.2284143, -0.2174443, -0.201331, -0.1833948, -0.1629359, 
    -0.1367965, -0.1136845, -0.08552697, -0.05474898, -0.01454714, 
    0.02985385, 0.07412463, 0.1117223, 0.1517452, 0.1936723 ;
}
