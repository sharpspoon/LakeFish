netcdf CGMR_SRA1B_1_pr-change_2070-2099 {
dimensions:
	time = 12 ;
	latitude = 48 ;
	longitude = 96 ;
	bounds = 2 ;
data:
 precipitation_flux_anomaly =
  1.153742e-007, 1.342489e-007, 1.585875e-007, 1.826777e-007, 1.980756e-007, 
    1.995658e-007, 1.936052e-007, 1.829261e-007, 1.657897e-007, 
    1.461699e-007, 1.312687e-007, 1.228248e-007, 1.233211e-007, 
    1.310201e-007, 1.49895e-007, 1.796973e-007, 2.117348e-007, 2.360732e-007, 
    2.544514e-007, 2.666206e-007, 2.76058e-007, 2.842536e-007, 2.961744e-007, 
    3.075988e-007, 3.197681e-007, 3.346695e-007, 3.483285e-007, 
    3.627331e-007, 3.753989e-007, 3.88065e-007, 4.024694e-007, 4.171222e-007, 
    4.282979e-007, 4.350036e-007, 4.379838e-007, 4.347551e-007, 
    4.315266e-007, 4.327685e-007, 4.431993e-007, 4.531337e-007, 
    4.610808e-007, 4.667929e-007, 4.702695e-007, 4.742433e-007, 
    4.804519e-007, 4.975882e-007, 5.278876e-007, 5.63402e-007, 6.03387e-007, 
    6.508226e-007, 7.039703e-007, 7.541375e-007, 7.911417e-007, 
    8.132452e-007, 8.189577e-007, 8.102652e-007, 7.975991e-007, 
    7.812077e-007, 7.665553e-007, 7.523986e-007, 7.372487e-007, 
    7.064532e-007, 6.632401e-007, 6.093478e-007, 5.427889e-007, 
    4.814458e-007, 4.325204e-007, 3.994894e-007, 3.853334e-007, 
    3.957641e-007, 4.300366e-007, 4.799556e-007, 5.388151e-007, 
    6.053738e-007, 6.711871e-007, 7.223477e-007, 7.514047e-007, 
    7.521498e-007, 7.297981e-007, 6.908067e-007, 6.43123e-007, 5.939494e-007, 
    5.450238e-007, 5.010655e-007, 4.481664e-007, 3.903001e-007, 
    3.341725e-007, 2.864887e-007, 2.470008e-007, 2.117346e-007, 
    1.774619e-007, 1.496463e-007, 1.258046e-007, 1.123936e-007, 
    1.044463e-007, 1.041982e-007,
  9.242585e-007, 8.172183e-007, 7.044666e-007, 6.110857e-007, 5.20437e-007, 
    4.136455e-007, 2.949333e-007, 1.724953e-007, 9.178063e-008, 
    8.184634e-008, 1.146287e-007, 1.665348e-007, 2.251459e-007, 
    2.683593e-007, 3.155465e-007, 3.537926e-007, 3.999863e-007, 
    4.523887e-007, 5.040461e-007, 5.368287e-007, 5.47011e-007, 5.278879e-007, 
    4.804524e-007, 4.451865e-007, 4.355007e-007, 4.129007e-007, 
    3.433619e-007, 2.425307e-007, 1.31517e-007, 5.601748e-008, 4.459321e-008, 
    6.073617e-008, 1.032045e-007, 1.692665e-007, 2.149634e-007, 
    2.395504e-007, 2.343351e-007, 2.08258e-007, 1.888865e-007, 2.102444e-007, 
    2.696007e-007, 3.339239e-007, 4.056982e-007, 4.77472e-007, 5.251557e-007, 
    5.542131e-007, 5.874924e-007, 5.949435e-007, 5.827737e-007, 
    6.297123e-007, 6.768992e-007, 7.216026e-007, 8.683792e-007, 
    9.945425e-007, 1.008202e-006, 1.011679e-006, 1.030306e-006, 
    1.002987e-006, 9.205337e-007, 7.69287e-007, 6.421301e-007, 5.668794e-007, 
    5.711013e-007, 6.590185e-007, 6.64234e-007, 5.532202e-007, 3.816081e-007, 
    2.589218e-007, 2.882275e-007, 3.975026e-007, 4.037115e-007, 
    2.735749e-007, 1.178576e-007, 5.651441e-008, 9.798941e-008, 
    1.469145e-007, 1.5362e-007, 1.24066e-007, 8.507459e-008, 2.671163e-008, 
    -2.295883e-008, -5.524475e-008, -7.436756e-008, -8.827533e-008, 
    -1.461415e-007, -2.410122e-007, -2.991267e-007, -2.459797e-007, 
    -8.256347e-008, 8.358438e-008, 2.231588e-007, 3.53544e-007, 5.1547e-007, 
    7.121657e-007, 8.87751e-007, 9.632504e-007,
  4.769754e-007, 3.880652e-007, 3.575178e-007, 3.622366e-007, 3.816082e-007, 
    3.446037e-007, 3.284607e-007, 3.316892e-007, 2.989068e-007, 
    2.432758e-007, 2.047808e-007, 2.561897e-007, 3.694385e-007, 
    4.071881e-007, 3.783795e-007, 3.026319e-007, 2.20427e-007, 1.556069e-007, 
    1.585872e-007, 2.455107e-007, 2.770516e-007, 3.041222e-007, 
    4.111622e-007, 4.851712e-007, 4.869098e-007, 4.903867e-007, 
    4.883999e-007, 4.496566e-007, 4.541271e-007, 4.690282e-007, 
    4.186127e-007, 3.339245e-007, 2.944364e-007, 2.869856e-007, 
    3.443554e-007, 4.523883e-007, 5.981715e-007, 6.530576e-007, 
    6.244967e-007, 4.75237e-007, 2.936911e-007, 8.358461e-008, 
    -1.898518e-007, -3.458172e-007, -3.428368e-007, -1.853812e-007, 
    1.595804e-007, 5.929569e-007, 7.968538e-007, 6.316995e-007, 
    5.199408e-007, 5.589322e-007, 1.051912e-006, 1.820067e-006, 
    2.240527e-006, 2.38631e-006, 2.468019e-006, 2.448151e-006, 2.2748e-006, 
    2.062707e-006, 1.89507e-006, 1.592575e-006, 1.414755e-006, 1.427421e-006, 
    1.161933e-006, 6.778928e-007, 5.778065e-007, 6.177916e-007, 
    5.507359e-007, 2.681104e-007, -5.573838e-009, -1.292533e-007, 
    -2.407637e-007, -2.725533e-007, -4.553413e-007, -8.161971e-007, 
    -1.098823e-006, -1.301727e-006, -1.271179e-006, -7.382143e-007, 
    1.106537e-008, 4.675376e-007, 6.801279e-007, 8.293878e-007, 
    9.210303e-007, 1.119961e-006, 1.297284e-006, 1.395135e-006, 
    1.450518e-006, 1.506397e-006, 1.562028e-006, 1.460949e-006, 
    1.175343e-006, 1.0159e-006, 8.942079e-007, 6.654752e-007,
  4.225863e-007, 2.897175e-007, 9.82368e-009, -2.586453e-007, -3.87789e-007, 
    -1.851331e-007, -1.004446e-008, 2.484906e-007, 4.225858e-007, 
    5.77558e-007, 4.730014e-007, 2.820184e-007, 2.974164e-007, 2.810253e-007, 
    3.085921e-007, 3.356624e-007, 2.221654e-007, 1.638025e-007, 
    1.558552e-007, 2.48739e-007, 3.955157e-007, 4.861646e-007, 2.753129e-007, 
    3.160426e-007, 3.781308e-007, 5.353381e-007, 5.293778e-007, 
    3.284608e-007, 2.566868e-007, 2.484911e-007, 3.570211e-007, 
    4.228348e-007, 3.681971e-007, 2.986584e-007, 2.792868e-007, 
    3.192716e-007, 4.191094e-007, 6.389012e-007, 1.115738e-006, 
    1.316904e-006, 7.27315e-007, -1.766884e-007, -6.714072e-007, 
    -8.422744e-007, -1.01761e-006, -7.772051e-007, 2.869956e-008, 
    9.741775e-007, 1.404821e-006, 1.355647e-006, 1.450022e-006, 
    1.877933e-006, 2.079099e-006, 1.439093e-006, -4.334861e-007, 
    -1.637748e-006, -1.167617e-006, 1.245617e-007, 1.395879e-006, 
    2.421079e-006, 2.160309e-006, 1.627344e-006, 1.978764e-006, 
    2.229101e-006, 1.826274e-006, 1.276173e-006, 7.990875e-007, 
    3.036239e-007, 1.456729e-007, 2.554452e-007, 3.170371e-007, 
    7.980957e-007, 7.625813e-007, 1.625622e-007, -4.52857e-007, 
    -8.442607e-007, -1.073987e-006, -5.325783e-007, 3.118207e-007, 
    5.89976e-007, 1.036514e-006, 1.688937e-006, 2.182661e-006, 2.244005e-006, 
    2.166767e-006, 1.939276e-006, 1.820812e-006, 1.685708e-006, 
    1.557558e-006, 1.387188e-006, 1.148024e-006, 1.128901e-006, 
    1.677264e-006, 1.676519e-006, 1.058617e-006, 5.293778e-007,
  -8.653706e-008, 1.546134e-007, 1.533715e-007, -2.25366e-007, 
    -3.917626e-007, 6.222649e-008, 7.22348e-007, 1.104563e-006, 8.50001e-007, 
    5.00072e-007, 2.48491e-007, 2.301128e-007, 5.805384e-007, 7.94867e-007, 
    1.208377e-007, 3.615241e-009, 4.47918e-007, 4.566106e-007, 3.786276e-007, 
    3.45845e-007, 3.883133e-007, 2.502295e-007, -3.326545e-007, 
    -1.068275e-006, -7.543572e-007, -4.481399e-008, 7.538847e-008, 
    -2.89938e-007, -6.788582e-007, -5.589038e-007, 2.070155e-007, 
    8.373349e-007, 1.143802e-006, 1.367071e-006, 8.912275e-007, 
    -8.802544e-009, -1.404296e-007, -4.754565e-008, 2.005586e-007, 
    6.893169e-007, 8.514912e-007, 1.205146e-006, 1.293064e-006, 
    1.403331e-006, 1.737862e-006, 1.560787e-006, 1.591085e-006, 
    7.285553e-007, -1.0442e-007, -1.190962e-006, -1.760435e-006, 
    -1.852822e-006, -4.148606e-007, -2.074867e-007, -1.173826e-006, 
    -1.603476e-006, -6.242226e-007, 6.175414e-007, 7.866702e-007, 
    1.164663e-006, 1.107045e-006, 1.171111e-007, 7.886501e-008, 
    5.383172e-007, 1.400846e-006, 1.777845e-006, 8.989255e-007, 
    5.087641e-007, 1.51138e-007, -4.384528e-007, -5.586553e-007, 
    2.335905e-007, 6.086025e-007, 3.344221e-007, 6.560376e-007, 1.13933e-006, 
    7.941198e-007, 7.702783e-007, 1.230725e-006, 1.294057e-006, 
    7.936264e-007, -4.804133e-008, -3.848081e-007, -2.76526e-007, 
    -2.37535e-007, 3.448522e-007, 1.017143e-006, 1.78033e-006, 1.785795e-006, 
    1.303493e-006, 1.269469e-006, 1.219054e-006, 1.823047e-006, 
    2.736985e-006, 2.182662e-006, 7.432095e-007,
  6.451105e-007, 7.531437e-007, 7.407255e-007, 9.838632e-007, 1.86626e-006, 
    2.110391e-006, 2.843777e-006, 2.976397e-006, 1.151253e-006, 8.96443e-007, 
    1.007705e-006, 1.285363e-006, 1.730908e-006, 2.095242e-006, 
    1.679002e-006, 8.512434e-007, -6.93999e-008, -1.050642e-006, 
    -6.224823e-007, -2.226343e-007, -4.943322e-007, -6.460759e-007, 
    -1.489233e-006, -2.004316e-006, -1.328548e-006, 2.949337e-007, 
    2.663728e-007, -8.76546e-007, -1.034002e-006, -6.808446e-007, 
    3.793725e-007, 3.103314e-007, 5.301235e-007, 1.718987e-006, 
    1.623102e-007, -1.629802e-006, -2.344561e-006, -1.976005e-006, 
    -9.902924e-007, -1.575909e-006, -1.733363e-006, -1.367542e-006, 
    -4.568328e-007, 1.595058e-006, 2.409405e-006, 3.767896e-006, 
    2.748408e-006, 7.136541e-007, 3.450987e-007, -1.155448e-006, 
    -1.784028e-006, -3.584846e-007, 7.971003e-007, 1.545884e-006, 
    1.191236e-006, 8.706047e-008, 8.802981e-007, 1.6415e-006, 1.217313e-006, 
    1.704581e-006, 1.196949e-006, 2.845009e-007, 1.906246e-007, 
    2.273737e-008, -8.579082e-008, 1.311191e-006, 1.421708e-006, 
    6.480905e-007, 5.03549e-007, -8.803909e-009, -2.248707e-007, 
    9.202722e-008, 3.664445e-008, 8.035477e-008, 6.023856e-008, 
    6.078553e-007, 5.557013e-007, -1.035246e-006, -5.025295e-007, 
    -4.853973e-008, -1.572184e-006, -1.148742e-006, -4.839003e-007, 
    -4.071603e-007, 3.138075e-007, 5.447764e-007, 6.500768e-007, 
    6.257378e-007, 8.611769e-007, 1.143554e-006, 1.437355e-006, 
    1.774618e-006, 1.363595e-006, 1.132378e-006, 1.672049e-006, 1.000751e-006,
  1.848378e-006, 1.695392e-006, 2.335895e-006, 4.227846e-006, 3.482041e-006, 
    2.584743e-006, 3.407039e-006, 3.237664e-006, 3.550836e-006, 3.99166e-006, 
    5.359091e-006, 6.293642e-006, 4.758325e-006, 3.701337e-006, 
    3.693886e-006, 3.463168e-006, 2.146649e-006, 2.141433e-006, 2.06817e-006, 
    -2.104653e-007, -1.294524e-006, -1.120429e-006, 6.967639e-008, 
    9.634996e-007, 1.398364e-006, 1.824039e-006, 1.706568e-006, 
    1.031297e-006, 1.349437e-006, 2.511976e-006, 3.050405e-006, 3.05736e-006, 
    3.146269e-006, 2.860414e-006, 3.678489e-006, 3.24114e-006, 
    -3.217292e-007, -1.341215e-006, -1.848866e-007, 1.310943e-006, 
    1.162924e-006, -2.42504e-007, -2.025181e-007, 1.893579e-006, 
    3.769884e-006, 4.675872e-006, 3.267217e-006, 2.066929e-006, 
    4.995745e-007, -1.030279e-006, 1.313178e-006, 3.371028e-006, 
    3.299006e-006, 3.098833e-006, 2.190856e-006, 1.428662e-006, 
    2.629697e-006, 3.565239e-006, 3.64993e-006, 2.216188e-006, 3.157938e-007, 
    9.6449e-007, 1.516082e-006, 2.018251e-006, 2.224384e-006, 7.106737e-007, 
    1.14379e-007, 2.243987e-007, 1.392899e-006, 1.929838e-006, 2.364951e-006, 
    2.658504e-006, 2.846755e-006, 1.880911e-006, 1.41227e-006, 1.714267e-006, 
    2.527126e-006, 1.824039e-006, 3.406285e-007, 7.737435e-008, 
    4.737458e-007, -4.324929e-007, -1.182269e-006, 8.115057e-007, 
    9.615114e-007, 1.454489e-006, 5.17939e-008, -4.464009e-007, 
    6.123355e-008, 8.028137e-007, 2.917031e-007, 3.585101e-007, 
    8.142388e-007, 1.383462e-006, 2.171238e-006, 2.168754e-006,
  2.394008e-006, 1.324602e-006, 2.430019e-006, 3.565488e-006, 3.853329e-006, 
    4.722812e-006, 3.064561e-006, 2.439953e-006, 3.169365e-006, 3.52898e-006, 
    4.428513e-006, 5.050389e-006, 5.259252e-006, 5.98345e-006, 6.410121e-006, 
    4.971414e-006, 4.648059e-006, 4.637877e-006, 3.751755e-006, 
    3.996629e-006, 3.63602e-006, 2.524145e-006, 3.077475e-006, 2.610572e-006, 
    4.702198e-006, 5.439062e-006, 3.772861e-006, 4.44416e-006, 4.565604e-006, 
    4.146881e-006, 1.425682e-006, -1.444041e-007, 6.090977e-007, 
    1.917419e-006, 4.286209e-006, 2.129015e-006, -5.007905e-007, 
    -4.414342e-007, 1.7545e-006, 2.259651e-006, 9.972737e-007, 1.444558e-006, 
    2.646833e-006, 2.732764e-006, 5.000472e-006, 6.629669e-006, 
    6.934397e-006, 4.990292e-006, 3.479806e-006, 4.184882e-006, 5.6221e-006, 
    4.614285e-006, 4.062196e-006, 2.489378e-006, 2.148392e-006, 
    1.001994e-006, 1.948714e-006, 4.763295e-006, 4.395483e-006, 
    4.137444e-006, 3.984956e-006, 4.335135e-006, 4.619747e-006, 
    2.250709e-006, 2.080338e-006, 2.237795e-006, 1.16069e-006, 3.970054e-007, 
    2.193838e-006, 1.872717e-006, -8.050229e-007, -4.737212e-007, 
    1.613191e-006, 7.317849e-007, 5.335987e-007, 2.282746e-006, 
    2.854207e-006, 1.9204e-006, 1.870732e-006, 4.886469e-007, 4.469239e-007, 
    7.397311e-007, 3.249816e-007, 1.365332e-006, 2.983101e-006, 
    3.443547e-006, 3.250328e-006, 2.484906e-006, 3.29975e-006, 3.775595e-006, 
    1.981991e-006, 1.75301e-006, 2.35005e-006, 3.82899e-006, 4.120059e-006, 
    3.062077e-006,
  3.348677e-006, 4.458067e-006, 5.607198e-006, 3.728906e-006, 3.169615e-006, 
    4.17147e-006, 4.294901e-006, 4.184137e-006, 4.863879e-006, 5.937506e-006, 
    6.923963e-006, 6.770234e-006, 7.732106e-006, 7.928054e-006, 
    7.580857e-006, 7.064284e-006, 7.238628e-006, 8.869807e-006, 
    8.436185e-006, 7.015109e-006, 5.992641e-006, 6.340088e-006, 
    7.308665e-006, 6.798298e-006, 5.971533e-006, 7.310649e-006, 
    7.508834e-006, 7.342686e-006, 7.213543e-006, 4.664698e-006, 
    3.745545e-006, 4.369407e-006, 2.993036e-006, 3.47658e-006, 3.422933e-006, 
    3.002475e-006, 3.330795e-006, 3.784038e-006, 2.928961e-006, 
    3.560027e-006, 5.426398e-006, 7.592282e-006, 7.309405e-006, 
    7.250052e-006, 4.434478e-006, 5.589565e-006, 6.150349e-006, 
    6.059203e-006, 7.082414e-006, 4.429014e-006, 5.257023e-006, 
    7.080676e-006, 6.047281e-006, 6.048271e-006, 5.133094e-006, 
    3.563258e-006, 4.160047e-006, 5.038224e-006, 4.662466e-006, 
    5.422424e-006, 5.465143e-006, 4.493584e-006, 1.593573e-006, 
    2.477209e-006, 4.113606e-006, 3.37699e-006, 3.236422e-006, 5.068274e-006, 
    6.49804e-006, 4.279505e-006, 3.379228e-006, 1.80045e-006, 2.330931e-006, 
    2.809009e-006, 8.259303e-008, 3.282148e-007, 3.227506e-007, 
    -2.102151e-007, -1.220487e-007, 1.057197e-008, 2.14715e-006, 
    2.385566e-006, 5.09759e-007, 3.305464e-006, 4.099697e-006, 2.117842e-006, 
    2.391029e-006, 3.81732e-006, 7.318598e-006, 6.304074e-006, 4.946332e-006, 
    3.848115e-006, 4.11311e-006, 5.037975e-006, 4.131731e-006, 4.577031e-006,
  1.778842e-006, 3.674022e-006, 6.738941e-006, 6.739687e-006, 6.358714e-006, 
    6.091734e-006, 3.213328e-006, 5.128373e-006, 7.607432e-006, 8.19553e-006, 
    7.512557e-006, 9.059053e-006, 1.158331e-005, 1.025661e-005, 
    9.116422e-006, 6.900866e-006, 6.425522e-006, 8.221357e-006, 
    7.629034e-006, 6.806744e-006, 4.94658e-006, 7.233413e-006, 7.671009e-006, 
    5.821774e-006, 6.057215e-006, 7.454444e-006, 7.601222e-006, 
    8.806726e-006, 8.908797e-006, 7.432838e-006, 6.778926e-006, 
    7.682436e-006, 8.359197e-006, 4.705182e-006, 3.395868e-006, 
    2.839557e-006, 4.924972e-006, 4.431e-006, 2.719107e-006, 5.073738e-006, 
    8.983801e-006, 7.849078e-006, 6.402177e-006, 7.699817e-006, 
    8.295612e-006, 6.971153e-006, 7.501631e-006, 6.423039e-006, 4.73374e-006, 
    8.099663e-006, 1.044958e-005, 7.01188e-006, 5.722186e-006, 6.379329e-006, 
    5.023818e-006, 6.123275e-006, 9.043657e-006, 7.79171e-006, 4.16253e-006, 
    3.290565e-006, 6.786875e-006, 4.894675e-006, 2.057786e-007, 1.10084e-006, 
    1.948716e-006, 1.786293e-006, 1.845896e-006, 1.557806e-006, 
    2.584004e-006, 3.447278e-006, 3.177071e-006, 2.243016e-006, 
    -2.983779e-007, -1.762668e-006, -1.378712e-006, 2.358265e-007, 
    2.313793e-006, 2.58872e-006, 1.20167e-006, 1.425686e-006, 1.532479e-006, 
    2.844028e-006, 3.178562e-006, 2.097977e-006, 3.64894e-006, 4.596155e-006, 
    4.734487e-006, 5.337241e-006, 7.923583e-006, 7.134322e-006, 
    5.220516e-006, 5.580128e-006, 6.590677e-006, 6.194057e-006, 
    4.866364e-006, 2.251954e-006,
  3.849604e-006, 5.843136e-006, 8.361925e-006, 7.60122e-006, 4.980851e-006, 
    4.687299e-006, 5.690645e-006, 4.997988e-006, 5.154947e-006, 
    6.709637e-006, 5.59279e-006, 6.06168e-006, 8.29214e-006, 9.231904e-006, 
    8.662928e-006, 7.937244e-006, 8.161504e-006, 7.097809e-006, 
    6.655493e-006, 5.505372e-006, 2.049543e-006, 4.347305e-006, 
    5.216538e-006, 4.547972e-006, 4.429759e-006, 4.718844e-006, 
    4.559155e-006, 3.668803e-006, 4.81073e-006, 8.38378e-006, 6.682811e-006, 
    4.281741e-006, 3.189982e-006, 4.326444e-006, 3.464413e-006, 
    3.130875e-006, 3.009432e-006, 2.96398e-006, 8.187126e-007, 3.309691e-006, 
    7.321327e-006, 7.771843e-006, 7.059316e-006, 5.763659e-006, 
    5.648675e-006, 7.788727e-006, 7.900984e-006, 4.061449e-006, 
    4.789621e-006, 5.067277e-006, 3.090638e-006, 2.148889e-006, 
    2.169256e-006, 4.834326e-006, 6.791097e-006, 8.202236e-006, 
    7.683922e-006, 5.355372e-006, 3.9713e-006, 4.37959e-006, 6.631406e-006, 
    4.09349e-006, 1.352671e-006, 2.509993e-006, 2.283743e-006, 
    -5.569746e-009, -8.137085e-007, 1.774373e-006, 7.859289e-007, 
    -4.116264e-007, -1.318364e-006, -3.870189e-006, -6.774424e-006, 
    -4.11556e-006, 7.591043e-007, 8.206989e-007, -7.518793e-007, 
    -2.895413e-006, -1.168359e-006, 2.472516e-007, 3.207642e-007, 
    1.024844e-006, 1.422208e-006, 1.782817e-006, 2.624978e-006, 
    1.424693e-006, 1.636787e-006, 4.093496e-006, 4.775464e-006, 
    2.716875e-006, 3.3909e-006, 7.742537e-006, 7.219011e-006, 2.493853e-006, 
    -2.370143e-008, 2.672165e-006,
  2.847446e-007, 1.826771e-006, 2.445671e-006, 3.299254e-006, 3.775851e-006, 
    3.997626e-006, 1.807897e-006, -8.11724e-007, -4.33236e-007, 
    -2.988781e-007, 3.263001e-006, 5.908445e-006, 4.225112e-006, 
    3.071509e-006, 5.289799e-006, 7.235642e-006, 3.814333e-006, 
    2.933924e-006, 2.639626e-006, 2.983343e-006, 4.074358e-006, 
    1.972301e-006, 3.545319e-007, -5.253823e-007, -1.009466e-007, 
    7.860945e-008, -3.264358e-008, 1.144792e-006, 2.81422e-006, 
    -1.285338e-006, -3.488723e-006, -6.569971e-007, -7.228155e-007, 
    -3.160112e-007, -1.419936e-006, -3.067507e-006, -2.339089e-006, 
    -1.126391e-006, 2.558914e-006, 2.32298e-006, 3.562513e-006, 
    3.798195e-006, 2.768029e-006, 2.191853e-006, 1.493474e-006, 
    5.293732e-007, 2.837813e-006, 2.31653e-006, 3.120193e-006, 
    -8.132156e-007, 1.42194e-007, -7.821727e-007, 1.630822e-006, 
    5.004695e-006, 3.842157e-006, 2.447656e-006, 1.275432e-006, 
    3.475583e-006, 6.230563e-006, 4.41585e-006, -7.804338e-007, 
    -1.484761e-006, 9.351897e-007, -7.141207e-007, -3.186968e-006, 
    -3.997589e-006, -2.731735e-006, -3.992127e-006, -6.248909e-006, 
    -5.744258e-006, -7.588525e-006, -7.690847e-006, -6.504464e-006, 
    -6.269025e-006, -6.147833e-006, -4.990012e-006, -6.635106e-006, 
    -6.677823e-006, -4.218628e-006, -1.478556e-006, -3.269175e-006, 
    -2.759803e-006, -1.007425e-006, -9.036194e-007, 3.51054e-007, 
    4.218156e-006, 7.643193e-006, 8.432206e-006, 7.740797e-006, 
    6.495058e-006, 8.326657e-006, 5.948426e-006, 1.703334e-006, 
    -1.726665e-006, 1.132372e-006, 1.886292e-007,
  1.069311e-007, -1.647677e-007, -1.60596e-006, -2.175429e-006, 
    -1.267452e-006, -3.051118e-006, -3.900488e-006, -2.935634e-006, 
    -2.53703e-006, -1.748758e-006, 5.693619e-007, 8.581919e-007, 
    -2.345809e-006, -3.804384e-006, -3.22075e-006, -2.222867e-006, 
    -5.77038e-007, -1.311902e-006, -2.358462e-006, -3.351623e-006, 
    -2.756085e-006, -4.522371e-006, -4.300586e-006, -3.986675e-006, 
    -5.278849e-006, -7.416667e-006, -6.885935e-006, -8.417526e-006, 
    -1.00877e-005, -9.088822e-006, -8.986251e-006, -7.748711e-006, 
    -5.58978e-006, -5.571652e-006, -6.755798e-006, -6.33633e-006, 
    -6.117281e-006, -4.116553e-006, -4.823367e-006, -8.253115e-006, 
    -8.252624e-006, -7.973227e-006, -5.320564e-006, -4.162004e-006, 
    -1.618631e-006, -6.999937e-006, -1.151846e-005, -4.901602e-006, 
    -6.399663e-006, -3.181263e-006, -1.019602e-006, -7.126364e-007, 
    2.606648e-007, 5.986731e-007, -2.786379e-006, -1.075729e-006, 
    3.383946e-006, 4.648558e-006, 3.963351e-006, -1.531202e-006, 
    -5.025029e-006, -5.067495e-006, -2.164252e-006, -4.582711e-006, 
    -5.246275e-007, -3.558256e-006, -5.997575e-006, -3.217765e-006, 
    -3.148225e-006, -3.476302e-006, -4.902589e-006, -5.786478e-006, 
    -3.303694e-006, -2.508719e-006, -4.383784e-006, -3.698331e-006, 
    -4.633126e-006, -6.525326e-006, -5.100528e-006, -1.612913e-006, 
    -2.317985e-006, -2.106637e-006, 3.139809e-006, 6.544473e-006, 
    6.271785e-006, 8.430965e-006, 9.312615e-006, 8.24569e-006, 4.985068e-006, 
    1.742264e-007, -1.809367e-006, -1.029912e-008, 3.915375e-007, 
    8.621646e-007, -9.058567e-009, -1.245106e-006,
  -3.71894e-006, -2.754587e-006, -1.95117e-006, -2.500278e-006, 
    -4.806231e-006, -4.74936e-006, -5.086126e-006, -5.62207e-006, 
    -3.384661e-006, -3.202369e-006, -3.458914e-006, -4.868816e-006, 
    -7.991854e-006, -7.00192e-006, -3.809102e-006, -4.833058e-006, 
    -6.926421e-006, -8.465217e-006, -8.967883e-006, -1.032935e-005, 
    -9.951107e-006, -8.286144e-006, -6.997196e-006, -7.937211e-006, 
    -8.838237e-006, -9.315572e-006, -9.452167e-006, -1.1211e-005, 
    -1.133989e-005, -1.010012e-005, -1.00949e-005, -8.278947e-006, 
    -8.119752e-006, -1.014631e-005, -9.97296e-006, -8.477629e-006, 
    -6.746362e-006, -7.146458e-006, -1.238297e-005, -1.177526e-005, 
    -1.148195e-005, -1.004473e-005, -7.95435e-006, -7.994086e-006, 
    -9.162834e-006, -1.15736e-005, -1.43693e-005, -1.542281e-005, 
    -1.105454e-005, -6.773938e-006, -6.602077e-006, -3.740799e-006, 
    -1.577893e-006, -4.028385e-006, 8.49257e-007, 1.216318e-006, 
    3.284622e-007, -1.048655e-006, -2.390243e-007, -3.921099e-006, 
    -3.616375e-006, -2.458797e-006, -4.526584e-006, -1.738825e-006, 
    -7.409435e-007, -1.65339e-006, 1.150509e-006, 9.314626e-007, 
    -1.689878e-007, -1.752485e-006, -2.746394e-006, -3.279607e-006, 
    -2.678845e-006, -1.876913e-006, -2.35375e-006, -3.226211e-006, 
    -4.825355e-006, -6.007515e-006, -5.082898e-006, -3.181754e-006, 
    -3.02107e-006, -2.243723e-007, 4.809737e-006, 5.372258e-006, 
    6.138423e-006, 7.653132e-006, 6.837283e-006, 7.806102e-006, 
    1.447279e-006, -3.814817e-006, -1.896293e-006, -2.348785e-006, 
    -4.092966e-006, -4.125006e-006, -4.473439e-006, -4.64778e-006,
  -1.399329e-006, -1.636506e-006, -1.099816e-006, -3.853052e-007, 
    -2.802522e-007, -1.241625e-006, -2.512694e-006, -9.666992e-007, 
    3.473342e-007, -3.893534e-006, -7.546056e-006, -7.918337e-006, 
    -7.941436e-006, -5.081904e-006, -2.216908e-006, -3.895768e-006, 
    -4.532792e-006, -7.946401e-006, -1.029582e-005, -7.680415e-006, 
    -6.804725e-006, -6.342789e-006, -7.17651e-006, -7.26393e-006, 
    -6.221097e-006, -6.273251e-006, -5.938471e-006, -4.870058e-006, 
    -4.864097e-006, -5.27686e-006, -4.322937e-006, -4.404645e-006, 
    -4.685532e-006, -4.144869e-006, -1.443537e-006, -2.155068e-006, 
    -4.25166e-006, -5.303185e-006, -5.447727e-006, -6.175153e-006, 
    -8.993957e-007, -3.254499e-007, -1.448501e-006, -3.35709e-006, 
    -3.974001e-006, -1.150082e-005, -9.580064e-006, -1.332722e-005, 
    -1.058291e-005, -8.71406e-006, -6.791808e-006, -2.423532e-006, 
    -4.453566e-006, -5.424954e-008, 1.311193e-006, -6.045993e-007, 
    2.025481e-007, 2.78492e-006, 3.884872e-006, -4.511185e-007, 
    1.375765e-006, -1.312155e-006, -6.69168e-007, 1.447292e-006, 
    2.249362e-008, 1.025837e-006, -3.699322e-006, -4.32964e-006, 
    -4.967909e-006, -3.622583e-006, -4.108857e-006, -3.238629e-006, 
    -3.005177e-006, -1.213561e-006, -1.124402e-006, -1.153957e-006, 
    -1.239887e-006, -1.834691e-006, -4.308532e-006, -3.307432e-006, 
    7.659335e-006, 8.467476e-006, 6.729009e-006, 2.819441e-006, 
    -2.14186e-007, -1.163638e-006, 2.50055e-006, -1.470118e-006, 
    -6.653238e-006, -9.317566e-006, -1.061744e-005, -5.695079e-006, 
    -4.11829e-006, -3.150713e-006, -7.031977e-007, -1.353328e-009,
  -6.865571e-007, -4.826593e-007, -2.785134e-007, -6.254625e-007, 
    -7.488936e-007, -2.25366e-007, 1.582642e-006, 8.403402e-006, 
    9.266923e-006, -4.234775e-006, -2.285447e-006, -2.021702e-006, 
    -1.454713e-006, 3.424675e-006, -2.159286e-007, -7.966521e-006, 
    -1.167442e-005, -7.367489e-006, -3.544597e-006, -3.520236e-007, 
    -1.187982e-006, -1.583112e-006, -2.639603e-006, -2.214671e-006, 
    -1.382938e-006, -1.317621e-006, -1.672765e-006, -1.449248e-006, 
    -2.313515e-006, -3.770102e-006, -9.324258e-007, 5.554548e-007, 
    1.536199e-006, 2.313046e-006, -1.965591e-007, -3.809841e-006, 
    -4.187833e-006, -4.104635e-006, -2.653263e-006, -1.466137e-006, 
    1.853596e-006, -2.161769e-006, -8.755285e-006, -4.018453e-006, 
    9.578798e-009, -5.702037e-006, -7.162103e-006, -7.092318e-006, 
    -6.27002e-006, -1.371511e-006, 5.163145e-006, 3.750267e-006, 
    4.063189e-006, 4.797321e-006, 5.191954e-006, 7.020824e-006, 
    4.581005e-006, 1.543902e-006, 4.59293e-006, 3.69091e-006, 1.055891e-006, 
    -2.171673e-007, 1.236691e-006, -3.52001e-006, -4.599598e-006, 
    -7.292738e-006, -7.740271e-006, -8.485576e-006, -5.897246e-006, 
    -3.462396e-006, -2.928188e-006, -2.125512e-006, -5.5493e-007, 
    -2.643569e-007, -5.760401e-007, 5.75078e-008, 1.844155e-007, 
    -1.071502e-007, -2.033621e-006, 7.908184e-006, 1.336822e-005, 
    1.678157e-005, 1.309677e-005, 9.627565e-007, 3.870962e-006, 
    2.001609e-006, -9.352083e-006, -1.980102e-005, -1.499242e-005, 
    -7.858482e-006, -3.097561e-006, -9.145424e-007, 8.855022e-008, 
    -2.539282e-007, -2.061686e-006, -1.294524e-006,
  6.900627e-007, 2.293677e-007, 1.82672e-008, 9.451196e-008, -1.627814e-007, 
    1.934558e-006, 4.730512e-006, 1.355125e-005, 1.532548e-005, 
    -1.679222e-006, 1.478586e-006, 1.821558e-006, 8.020192e-006, 
    3.325578e-006, -4.131463e-006, -7.010367e-006, -9.936206e-006, 
    -5.398553e-006, -1.304943e-007, 4.820167e-006, 2.869604e-006, 
    1.616664e-006, 9.826199e-007, 1.250097e-006, 1.075009e-006, 
    4.196063e-007, -2.70069e-007, -5.785232e-007, -2.870322e-006, 
    -1.950174e-006, 2.189119e-006, 2.300381e-006, 4.12602e-006, 
    5.370757e-007, -2.481899e-006, -2.384793e-006, -5.484978e-006, 
    -2.68828e-006, 2.527622e-006, 6.729005e-006, 5.642964e-006, 
    -3.074962e-006, -7.021041e-006, 4.691026e-006, 6.027911e-006, 
    -2.002575e-006, -5.206566e-007, 6.990525e-006, 5.015623e-006, 
    6.626937e-006, 1.049428e-005, 8.280966e-006, 1.194094e-005, 
    1.089562e-005, 7.905455e-006, 6.315007e-006, 1.769655e-006, 
    -2.055021e-007, 1.225817e-007, -3.851568e-006, -2.160526e-006, 
    -6.348753e-006, -8.065112e-006, -9.283778e-006, -1.313325e-005, 
    -1.187286e-005, -9.704492e-006, -6.117534e-006, -1.454464e-006, 
    -8.820107e-007, -9.870473e-008, -4.41185e-007, -4.036829e-007, 
    -2.516913e-007, -3.649407e-007, 4.677863e-007, -1.675016e-008, 
    -1.709769e-007, -4.53677e-006, 1.860347e-005, 9.257234e-006, 
    1.496165e-005, 1.056083e-005, 7.933268e-006, 1.111615e-005, 
    -9.936713e-006, -1.97521e-005, -1.033059e-005, -2.355493e-006, 
    7.851831e-007, 1.805414e-006, 3.750264e-006, 1.008945e-006, 
    -1.196673e-006, -6.706618e-007, -4.228059e-007,
  -6.120508e-007, -6.97733e-007, 6.44618e-008, 5.403064e-008, 3.812846e-006, 
    1.328055e-005, 8.224588e-006, 1.026977e-005, 3.518795e-006, 
    -3.001947e-006, -1.90597e-006, 4.878773e-006, 5.131351e-006, 
    6.746137e-006, -2.087269e-006, -5.341684e-006, -1.132698e-005, 
    -7.179493e-006, -2.261606e-006, 1.332301e-006, 5.339722e-006, 
    2.554196e-006, 3.335514e-006, 1.272448e-006, 1.325844e-006, 
    -6.344035e-007, -1.501898e-006, -6.478131e-007, -4.332126e-006, 
    -2.502512e-006, 1.586366e-006, 4.527111e-006, 4.208473e-006, 
    -9.560208e-007, -2.494068e-006, -3.057083e-006, -8.646248e-007, 
    3.687679e-006, 7.15046e-006, 8.653244e-006, 5.476319e-006, 
    -5.448966e-006, -3.910176e-006, -5.226411e-007, 8.563346e-006, 
    7.066024e-006, 6.730494e-006, -9.957621e-007, 5.601731e-006, 
    1.968407e-005, 1.752142e-005, 2.144241e-005, 1.757109e-005, 
    7.112216e-006, 5.558028e-006, 1.771143e-006, 3.683948e-006, 
    5.813075e-006, 1.141809e-006, -3.957619e-006, -9.757889e-006, 
    -1.355545e-005, -1.736667e-005, -1.635041e-005, -1.212692e-005, 
    -6.359183e-006, -2.612781e-006, -8.089964e-007, 9.60008e-008, 
    1.272938e-007, 2.837551e-007, -5.951633e-007, -7.481485e-007, 
    -7.615599e-007, -5.60394e-007, -9.778746e-007, -1.113227e-006, 
    -5.395324e-007, -1.176011e-005, 6.445371e-006, 8.051731e-006, 
    6.723276e-006, 6.966427e-006, 1.254418e-005, 3.8707e-006, -1.903659e-005, 
    -2.236749e-005, -1.144818e-005, -2.093722e-006, -5.447455e-007, 
    1.981496e-006, 2.14216e-007, -1.452229e-006, -1.298002e-006, 
    -8.738152e-007, -9.17029e-007,
  -8.137131e-007, -5.266179e-007, 1.152494e-006, 4.667927e-007, 
    7.708511e-006, 1.086508e-005, 1.635938e-005, 1.168687e-005, 
    4.165009e-006, -5.368747e-006, -1.345696e-006, 1.201045e-005, 
    4.363683e-006, -4.152076e-006, -5.161386e-006, -2.096133e-005, 
    -1.740045e-005, -1.022008e-005, -1.81929e-006, 1.275181e-006, 
    1.830747e-006, 3.681718e-006, 6.093469e-006, 1.527505e-006, 
    2.951064e-006, 3.587575e-007, -1.998355e-006, -3.420424e-006, 
    -2.977114e-006, -2.966226e-008, 6.696962e-006, 6.556147e-006, 
    -2.692497e-006, 2.4775e-007, -3.278614e-006, 3.236915e-006, 
    2.356506e-006, 2.516446e-006, 6.997227e-006, 9.2478e-006, 7.855286e-006, 
    9.141502e-006, 9.045889e-006, 9.138283e-006, 1.812566e-005, 1.65352e-005, 
    1.931502e-005, 1.101508e-005, 3.121584e-005, 3.576093e-005, 
    1.722364e-005, 3.16666e-005, 2.88607e-005, 2.105646e-005, 1.454318e-005, 
    6.245456e-006, 1.068253e-005, 7.442271e-006, 1.572465e-006, 
    3.962559e-007, -1.012446e-005, -1.419918e-005, -1.310593e-005, 
    -1.020318e-005, -4.833551e-006, -2.182384e-006, 3.652149e-007, 
    3.095847e-007, 7.953622e-007, -4.250423e-007, -9.40624e-007, 
    -8.815159e-007, -1.084916e-006, -1.16091e-006, -1.744788e-006, 
    -9.93522e-007, -1.089384e-006, -1.166126e-006, -1.842341e-005, 
    1.335578e-005, 1.688836e-005, 6.261085e-006, 9.460637e-006, 
    7.998315e-006, -9.160882e-006, -2.41812e-005, -2.353872e-005, 
    4.757385e-008, 4.717622e-007, 3.572677e-007, 1.100587e-006, 
    -6.950022e-007, -6.527825e-007, -5.906941e-007, -7.692588e-007, 
    -6.224827e-007,
  -2.234291e-006, -7.628014e-007, 1.923636e-007, 2.565868e-006, 
    1.358131e-005, 1.125995e-005, 1.193076e-005, -6.575137e-007, 
    -2.162025e-006, -1.003216e-006, -5.387872e-006, 1.148022e-005, 
    1.007258e-005, -3.940972e-006, -8.561576e-006, -2.499384e-005, 
    -2.457958e-005, -6.922201e-006, -1.193221e-007, 4.999714e-006, 
    3.097346e-006, 2.857689e-006, 4.988304e-006, 7.64096e-006, 2.884506e-006, 
    -5.02032e-007, 1.034277e-006, -2.839774e-006, 2.296163e-006, 
    7.359817e-006, 9.346637e-006, 1.785941e-005, 2.68357e-006, 1.738106e-006, 
    -2.962959e-006, 4.854939e-006, 2.681358e-006, -2.8512e-006, 
    1.017018e-005, 1.099049e-005, 7.452451e-006, 1.877038e-005, 
    1.866979e-005, 2.54759e-005, 2.888006e-005, 2.339469e-005, 3.674713e-005, 
    5.382289e-005, 3.993772e-005, 2.350969e-005, 2.891633e-005, 3.39457e-005, 
    3.390398e-005, 1.666259e-005, 2.199051e-005, 1.511635e-005, 
    1.076199e-005, 1.191757e-005, 7.095063e-006, -8.44957e-006, 
    -1.219796e-005, -1.477114e-005, -1.166623e-005, -7.542581e-006, 
    -2.62967e-006, -9.681899e-007, 6.81368e-007, -4.43918e-007, 
    -5.584088e-007, -5.467355e-007, -1.39362e-006, -2.3612e-006, 
    -1.56374e-006, -2.549948e-006, -1.644949e-006, -2.263592e-007, 
    -9.239822e-007, -1.359717e-005, -3.927484e-005, 1.729913e-005, 
    1.747347e-005, 9.856245e-006, 1.05479e-005, -1.518303e-006, 
    -1.804892e-005, -1.586066e-005, -8.910014e-006, -1.923359e-006, 
    4.116628e-007, -1.749756e-006, -4.871308e-007, -6.286928e-007, 
    -1.348667e-006, -1.617135e-006, -1.583609e-006, -1.964332e-006,
  -1.531949e-006, -3.182504e-007, 3.330299e-006, 1.510743e-005, 
    3.028003e-005, 2.052101e-005, 8.351228e-006, -1.978013e-006, 
    1.483539e-006, 6.777162e-006, -9.761359e-006, -1.080953e-006, 
    7.479044e-006, 6.918985e-006, 6.143018e-007, 5.650138e-006, 
    -7.668517e-006, -5.524489e-006, -4.865113e-006, 8.172137e-007, 
    2.974404e-006, -5.844959e-007, -9.962605e-007, 8.332372e-006, 
    5.114471e-006, 2.980629e-006, 1.123388e-005, 1.573925e-005, 
    1.705873e-005, 1.71618e-005, 2.089751e-005, 1.960136e-005, 
    -2.420275e-007, -3.865236e-006, -6.978582e-006, 8.921466e-006, 
    1.223473e-005, 1.062614e-005, 1.596251e-005, 2.302168e-005, 
    1.594088e-005, 3.179288e-006, 1.142758e-005, 2.00777e-005, 3.715392e-005, 
    4.967638e-005, 6.172e-005, 5.577345e-005, 3.120142e-005, 2.276861e-005, 
    2.808982e-005, 6.119517e-006, 2.726603e-005, 6.498522e-006, 
    1.081912e-005, 8.802977e-006, 1.175266e-005, 1.591953e-005, 
    5.173075e-006, -7.66282e-007, -6.459766e-006, -9.552254e-006, 
    -8.376795e-006, -5.485972e-006, -2.77272e-006, -1.588328e-006, 
    -1.806638e-007, -1.970294e-006, -1.794957e-006, -2.124272e-006, 
    -2.009285e-006, -1.88461e-006, -2.641341e-006, -1.238644e-006, 
    -1.796693e-007, 9.312125e-007, 1.100116e-005, 1.45621e-006, 
    2.090994e-006, 6.167735e-006, 5.639464e-006, 3.045177e-006, 
    8.872303e-007, -2.336912e-005, -2.090522e-005, -2.273533e-006, 
    -2.199013e-007, -4.233043e-006, -2.929182e-006, -3.365039e-006, 
    -2.536537e-006, -2.044054e-006, -1.357607e-006, -7.002182e-007, 
    -1.846861e-006, -1.475822e-006,
  3.6467e-006, 1.963863e-006, 9.175528e-006, 1.052408e-005, 9.429092e-006, 
    9.732081e-006, 1.110523e-005, 1.197717e-005, 1.040686e-005, 
    1.356988e-005, 6.632399e-006, 6.621696e-006, 1.762433e-006, 
    -2.397232e-006, 9.23741e-007, 2.419341e-005, 9.10028e-006, 
    -9.970492e-006, -7.384646e-006, -5.939721e-006, 3.550071e-006, 
    1.563028e-006, 5.74837e-007, 4.537287e-006, 6.651269e-006, 8.820381e-006, 
    1.739699e-005, 2.323352e-005, 2.557376e-005, 2.933604e-005, 
    3.670889e-005, 2.227512e-005, 9.064745e-006, 6.705392e-006, 
    -2.102679e-006, 3.871195e-006, 9.162344e-006, 6.794071e-006, 
    1.221884e-005, 3.38573e-005, 2.570513e-005, 3.197281e-005, 2.326979e-005, 
    2.53731e-005, 6.608007e-005, 7.490108e-005, 8.341213e-005, 7.321501e-005, 
    6.358812e-005, 5.817004e-005, 4.710544e-005, 4.245725e-006, 
    9.337935e-006, 5.060065e-006, 1.54052e-005, 7.338451e-006, 7.684401e-006, 
    1.240856e-005, 1.412916e-005, 1.20733e-005, 7.632509e-006, 2.882225e-007, 
    -8.299317e-006, -8.083991e-006, -6.366879e-006, -2.893667e-006, 
    -6.40116e-007, -8.700918e-007, -1.731129e-006, -1.939993e-006, 
    -2.515178e-006, -2.065659e-006, -8.477377e-007, 3.378977e-007, 
    1.164912e-006, 1.650962e-005, 3.089619e-005, -1.04319e-006, 
    3.118948e-006, -1.009612e-007, 2.558394e-006, -2.031898e-006, 
    -8.511917e-006, -1.235469e-005, -1.225087e-005, 5.039714e-006, 
    3.366064e-006, 3.128636e-006, -7.789458e-007, 5.328511e-007, 
    -1.048153e-006, -1.829474e-006, -1.700582e-006, 3.664572e-007, 
    5.055426e-008, 4.278008e-007,
  1.203804e-005, 1.168116e-005, 1.233508e-005, 5.793214e-006, -8.067564e-007, 
    -2.688281e-006, 3.697103e-006, 1.031793e-005, 2.738622e-005, 
    2.906186e-005, 1.524154e-005, 1.051016e-005, 5.836155e-006, 9.29099e-006, 
    -1.226504e-005, 2.201283e-006, -2.463275e-006, -1.224144e-005, 
    6.4286e-007, -3.185989e-006, 4.008783e-006, 9.421128e-007, 7.198119e-006, 
    1.844354e-005, 6.92271e-006, 7.022063e-006, 1.632608e-005, 6.716313e-006, 
    5.529444e-006, 2.657958e-005, 1.961354e-005, 1.337168e-005, 4.63333e-008, 
    -6.892646e-006, -2.435657e-005, -1.312356e-005, 7.409981e-006, 
    1.853815e-005, 1.811149e-005, 4.494378e-005, 4.376037e-005, 
    4.020073e-005, 3.114603e-005, 1.472249e-005, 3.818884e-005, 
    3.547881e-005, 4.625632e-005, 4.645353e-005, 4.430948e-005, 
    3.684151e-005, 3.358984e-005, 1.616888e-005, 2.558617e-005, 
    2.872312e-005, 2.761844e-005, 2.619935e-005, 2.904696e-005, 
    2.797904e-005, 2.971726e-005, 2.978332e-005, 2.736363e-005, 
    2.311184e-005, 2.236851e-005, 1.558625e-005, 1.224865e-005, 
    1.250767e-005, 9.916113e-006, 8.375338e-006, 6.851197e-006, 
    6.795315e-006, 5.494444e-006, 5.806374e-006, 5.153207e-006, 
    4.502523e-006, 6.697962e-006, 1.065744e-005, 4.065923e-006, 
    6.346541e-006, -3.781541e-006, 8.612507e-006, 6.026905e-006, 
    -3.864239e-006, -9.294221e-006, -1.56287e-005, -4.052235e-006, 
    2.531342e-006, 5.610666e-006, 1.182371e-005, 5.874921e-006, 
    5.508355e-006, 4.554433e-006, 4.515183e-006, 8.224342e-007, 
    4.772983e-006, 5.221258e-006, 7.019335e-006,
  3.963352e-006, 3.668305e-006, 2.305344e-006, 3.314344e-007, -4.565882e-007, 
    1.523804e-007, 4.622227e-006, 1.019749e-005, 3.93114e-005, 2.75211e-005, 
    8.945806e-006, -5.817528e-007, 5.871196e-006, 1.214631e-005, 
    -3.98171e-006, -1.108856e-007, 5.54038e-006, 1.650763e-005, 
    -4.724287e-006, 2.018873e-005, 1.267182e-005, 6.491071e-006, 
    1.560611e-005, 5.960093e-006, 6.288421e-006, 7.704519e-006, 
    7.120136e-006, 4.008052e-006, 9.716823e-007, -3.75323e-006, 
    3.231435e-006, 2.057639e-005, 2.357252e-005, 3.190231e-006, 
    -1.152193e-005, 1.432338e-005, 1.44304e-005, 1.509425e-005, 
    1.101034e-005, 6.650036e-006, 4.813715e-006, 6.294125e-006, 
    2.500179e-005, 1.929293e-005, 9.072974e-006, 1.528997e-005, 
    1.124106e-005, 4.03585e-006, 7.068738e-006, -7.543094e-006, 
    -1.434621e-005, -7.347131e-006, 4.265341e-006, 1.24811e-005, 
    1.379614e-005, 1.217216e-005, 1.385152e-005, 1.170575e-005, 
    1.181552e-005, 8.936613e-006, 9.56246e-006, 7.444509e-006, 7.711736e-006, 
    9.014844e-006, 8.953501e-006, 9.405504e-006, 8.412093e-006, 
    9.093076e-006, 1.268252e-005, 9.950887e-006, 1.341988e-005, 
    1.133968e-005, 1.066838e-005, 1.287475e-005, 5.626065e-006, 
    1.145341e-005, 1.640235e-005, 1.845299e-005, 1.283749e-005, 
    5.456201e-006, 2.316025e-006, -3.998091e-006, -4.958223e-006, 
    -1.285336e-005, -2.695483e-006, -4.894155e-006, -4.884212e-006, 
    3.023335e-006, 4.815451e-006, 1.301258e-006, 1.719727e-006, 
    4.327936e-006, 2.863144e-006, 1.775117e-006, 1.859311e-006, 3.991914e-006,
  -2.116078e-006, 4.416837e-006, 1.348442e-006, -7.581824e-006, 
    -2.487857e-006, 6.451082e-007, 3.15621e-006, 5.191456e-006, 
    1.333718e-005, 7.327288e-006, 3.353396e-006, 1.728673e-006, 4.95825e-006, 
    1.154457e-005, 2.037076e-005, 2.993879e-005, 1.09706e-005, 9.679919e-006, 
    3.219793e-006, 4.32568e-006, 7.283554e-006, 3.475579e-006, 1.015005e-005, 
    1.1365e-005, 1.210907e-005, 1.167072e-005, -1.500831e-005, 
    -1.573244e-007, -3.08812e-006, -2.891558e-005, 9.587748e-007, 
    2.740014e-005, 4.682312e-006, 3.662077e-006, -1.508777e-005, 
    -1.633799e-005, -1.20723e-005, -2.008639e-005, -1.53426e-005, 
    -1.489806e-005, -7.260722e-006, -1.452329e-005, -7.56693e-006, 
    1.321103e-006, -4.020207e-006, -1.675071e-007, 8.939583e-006, 
    6.898619e-006, 1.497529e-005, 5.589558e-006, -4.225589e-006, 
    -7.694078e-006, -6.859616e-006, -3.972018e-006, -2.525117e-006, 
    2.109398e-006, 7.190944e-006, 1.048336e-005, 9.349873e-006, 
    9.119402e-006, 8.10513e-006, 6.077575e-006, 5.315381e-006, 5.662827e-006, 
    4.707166e-006, 3.089397e-006, 1.438098e-006, 2.020237e-006, 
    2.091515e-006, 2.305595e-006, 4.645826e-006, 5.940489e-006, 
    6.190579e-006, 1.227e-005, 1.550678e-005, 2.701568e-005, 1.408745e-005, 
    3.691901e-006, 8.699684e-006, 5.819289e-006, -1.714729e-007, 
    -1.986684e-006, -6.233018e-006, -1.303589e-005, -1.263778e-005, 
    -1.499689e-005, -1.427294e-005, -9.912115e-006, -9.564672e-006, 
    -6.723016e-006, -4.16498e-006, -4.147352e-006, -3.889561e-006, 
    -3.579869e-006, 2.660741e-006, -7.588242e-007,
  -1.436829e-006, -1.000473e-006, -1.964083e-006, -2.242735e-006, 
    -9.416153e-007, 1.70508e-007, -6.59486e-007, -6.627147e-007, 
    1.033285e-006, 8.991744e-007, 7.63897e-006, 3.807882e-006, 9.237619e-007, 
    6.808714e-007, 4.484149e-006, 1.437429e-005, 1.983258e-005, 
    2.553128e-005, 8.651754e-006, -2.26366e-007, -2.185116e-006, 
    -1.190783e-007, 5.77802e-007, -4.357171e-007, 1.151166e-007, 
    1.110026e-005, 2.959514e-006, -3.526466e-006, -1.150978e-005, 
    -5.866954e-006, -2.793833e-006, 2.655022e-006, -4.220637e-006, 
    -9.552969e-007, -5.108981e-006, -1.033528e-006, 5.926064e-006, 
    3.72839e-006, 4.355992e-006, 6.449856e-006, 3.843394e-006, 2.910092e-006, 
    2.869274e-008, -2.76478e-006, -2.435205e-006, 3.712765e-006, 
    2.798086e-006, -1.863256e-006, 2.247725e-006, 6.787621e-006, 
    4.161782e-006, 3.962105e-006, 2.587978e-006, -1.283846e-006, 
    -6.481871e-006, -8.361407e-006, -7.967017e-006, -3.129109e-006, 
    -1.579381e-006, -2.060442e-006, -3.026285e-006, -2.797795e-006, 
    1.232711e-006, 7.504023e-007, 2.308072e-006, 2.78715e-006, 5.12664e-006, 
    8.362178e-006, 8.234276e-006, 8.071109e-006, 4.671656e-006, 
    4.527859e-006, 9.812806e-006, 1.13953e-005, 1.991927e-005, 1.005867e-005, 
    3.288079e-006, 1.269717e-006, 2.036879e-006, -1.059831e-006, 
    -1.478305e-006, -4.577499e-006, -4.413586e-006, -3.371996e-006, 
    -7.390341e-006, -4.45084e-006, -4.773201e-006, -6.575744e-006, 
    -5.742519e-006, -6.649256e-006, -6.216875e-006, -7.062019e-006, 
    -3.624071e-006, 1.131635e-006, -2.981585e-006, -1.217783e-006,
  8.830057e-010, -1.426645e-008, -8.703375e-008, -7.809308e-008, 
    -5.59896e-008, 2.00062e-007, -2.673378e-007, -1.324823e-007, 
    4.074364e-007, 1.737365e-007, 5.735594e-006, 4.679599e-006, 1.491e-006, 
    2.018252e-006, 1.258789e-006, 2.3334e-007, 4.059711e-006, 5.877902e-006, 
    4.559151e-006, 1.246373e-006, 1.424414e-007, -1.348171e-006, 
    -2.436449e-006, -2.432225e-006, -1.394612e-006, -9.791174e-007, 
    -2.950043e-006, -1.779804e-006, -5.222222e-006, -4.736444e-006, 
    -2.374611e-006, -3.797923e-006, -6.267295e-006, -1.433855e-006, 
    1.210105e-006, 5.795446e-007, 1.763685e-006, 2.656525e-006, 
    1.511116e-006, -8.338266e-007, 4.312806e-007, -1.881877e-006, 
    -5.586803e-006, -6.910524e-006, -7.364015e-006, -6.49975e-006, 
    -4.607549e-006, -4.578991e-006, -4.07409e-006, -2.841513e-006, 
    -2.488605e-006, -2.581735e-006, -9.748928e-007, -1.203627e-006, 
    -7.157632e-006, -6.323417e-006, -8.716797e-006, -1.157559e-005, 
    -2.142153e-005, -2.519277e-005, -2.762637e-005, -2.767852e-005, 
    -2.674695e-005, -2.041023e-005, -2.057638e-005, -1.524249e-005, 
    -1.273986e-005, -2.77596e-006, 4.737954e-006, 8.598108e-006, 
    9.628031e-006, 1.129125e-005, 5.436577e-006, 1.709798e-006, 
    3.762928e-006, 1.682231e-006, -8.596589e-007, -9.597397e-008, 
    -8.012956e-007, -1.466632e-006, -2.342574e-006, -1.436086e-006, 
    -1.630547e-006, -2.245468e-006, -7.11394e-007, -1.078707e-006, 
    -1.417212e-006, -2.225349e-006, -2.520394e-006, -3.972263e-006, 
    -3.253778e-006, -2.731989e-006, -1.286329e-006, -1.248082e-006, 
    -8.926884e-008, -3.065747e-008,
  -3.162634e-007, -1.896034e-007, -3.289284e-008, -1.496186e-007, 
    -1.148492e-007, 1.270464e-007, 1.975801e-008, 1.238177e-007, 
    2.400468e-007, 4.071881e-007, 7.809588e-007, 7.337721e-007, 
    1.267979e-006, 2.653783e-007, -2.410125e-007, -1.563988e-006, 
    2.035376e-007, 8.974366e-007, 2.20079e-006, -3.833184e-007, 
    -3.410983e-007, 1.638018e-007, -1.992903e-007, -1.300486e-006, 
    -1.004447e-006, -2.089252e-006, -1.055609e-006, 1.345962e-006, 
    -5.300944e-008, -8.139623e-007, 1.999628e-006, 2.474977e-006, 
    1.952934e-006, 4.075606e-006, 3.484525e-006, -1.341214e-006, 
    1.65046e-007, 1.486034e-006, 1.812121e-006, 1.322367e-006, 
    -2.100182e-006, -7.096551e-007, -1.078459e-006, -1.918885e-006, 
    -1.551571e-006, -3.713481e-006, -3.217271e-006, -3.229939e-006, 
    -1.786761e-006, -1.835934e-006, -2.223861e-006, -3.076952e-006, 
    -4.991006e-006, -3.406263e-006, -5.155911e-006, -2.854924e-006, 
    -5.934251e-006, -9.966998e-006, -1.853542e-005, -1.716576e-005, 
    -1.779682e-005, -2.040775e-005, -2.133957e-005, -1.7581e-005, 
    -2.393212e-005, -2.807142e-005, -2.813648e-005, -1.883767e-005, 
    -3.475561e-006, 5.409262e-006, 6.442903e-006, 3.390898e-006, 
    7.871683e-007, -2.304574e-006, -7.409481e-007, 2.730776e-007, 
    3.341711e-008, -1.228462e-006, -1.976749e-006, -1.236162e-006, 
    -6.36639e-007, -6.840755e-007, -2.510459e-006, -3.512812e-006, 
    -1.334511e-006, -1.678231e-006, -7.6777e-007, -2.026669e-006, 
    -2.312522e-006, -1.832208e-006, -2.043308e-006, -1.426151e-006, 
    -9.659536e-007, -8.797754e-007, -7.128826e-007, -4.548441e-007,
  -7.630497e-007, -7.829179e-007, -7.528674e-007, -3.505359e-007, 
    -2.924213e-007, -4.481376e-008, 1.123934e-007, 9.128357e-008, 
    3.912953e-008, 2.293676e-007, 1.032043e-007, 3.458449e-007, 
    2.787897e-007, 7.638209e-008, -2.032627e-007, 7.563767e-008, 
    -1.036237e-006, 5.114966e-007, 1.082211e-006, 1.761704e-006, 
    -1.673759e-006, 1.695641e-006, 1.999874e-006, 2.398065e-008, 
    -1.285335e-006, -5.045149e-007, 1.578451e-008, 7.310398e-007, 
    3.06607e-007, 9.585328e-007, 2.607347e-006, -8.462466e-007, 
    -1.068984e-007, 7.83989e-006, 8.093211e-006, 5.969323e-007, 
    -1.525992e-006, 4.677859e-007, 2.415119e-006, 2.465286e-006, 6.4511e-007, 
    6.895634e-007, -3.51034e-007, -9.359046e-007, -1.212569e-006, 
    -1.736842e-006, -1.633527e-006, -7.374711e-007, -1.219027e-006, 
    1.019607e-007, -5.052616e-007, -1.688909e-006, -3.369016e-006, 
    -3.234405e-006, -8.360621e-007, -6.522805e-007, -1.428134e-006, 
    -5.620082e-006, -1.349212e-005, -1.774938e-005, -1.938131e-005, 
    -1.239838e-005, -1.354577e-005, -1.282629e-005, -1.787033e-005, 
    -1.729614e-005, -2.30075e-005, -2.996386e-005, -9.399759e-006, 
    7.831914e-007, 1.634795e-006, -8.427724e-007, -3.469842e-006, 
    -3.363049e-006, 1.203658e-006, 2.787883e-007, 4.680332e-007, 
    -1.027546e-006, -1.564236e-006, -7.185963e-007, 9.451105e-008, 
    -1.409515e-006, -1.887095e-006, -2.539022e-006, -4.35125e-006, 
    -2.409381e-006, -4.122518e-006, -2.617749e-006, -3.104518e-006, 
    -2.410373e-006, -7.786962e-007, -2.160779e-006, -1.743298e-006, 
    -1.041204e-006, -1.061818e-006, -9.003885e-007,
  -1.162649e-006, -5.050111e-007, -5.271145e-007, -1.057844e-006, 
    -1.050642e-006, -1.099816e-006, -3.207335e-007, 1.561036e-007, 
    2.1695e-007, -7.312536e-009, -5.320817e-007, 6.865849e-007, 
    9.977711e-007, 4.022215e-007, -9.945131e-008, 6.694472e-008, 
    -7.921067e-007, -1.061818e-006, -3.972262e-007, 3.595044e-007, 
    7.134068e-007, 1.238177e-006, 2.433996e-006, 1.328329e-006, 
    -2.936622e-007, -9.654564e-007, -1.08566e-006, 3.649666e-007, 
    2.523649e-006, 1.812366e-006, -6.502987e-007, -2.65674e-006, 
    -6.175123e-007, 4.9138e-006, 6.937376e-006, 1.930835e-006, 3.610445e-006, 
    2.212217e-006, 1.717746e-006, 9.632486e-007, 8.067855e-007, 
    8.542211e-007, 9.62491e-008, -2.938869e-006, -1.79893e-006, 
    -3.28085e-006, -2.802772e-006, -2.147121e-006, -2.081059e-006, 
    -1.0571e-006, -1.330785e-006, -4.109603e-006, -2.076338e-006, 
    -1.268447e-006, -8.127208e-007, 2.891215e-006, 5.574169e-006, 
    3.094367e-006, -2.731738e-006, -1.166399e-005, -1.551396e-005, 
    -1.065618e-005, -7.333221e-006, -6.750586e-006, -8.306266e-006, 
    -8.273484e-006, -1.493058e-005, -1.707685e-005, -8.770188e-006, 
    -2.332883e-006, -1.474576e-006, -4.991256e-006, -2.004315e-006, 
    -1.592545e-006, -2.36244e-006, 1.128938e-007, 4.140429e-006, 
    3.27045e-006, 7.134058e-007, 6.542978e-007, 1.65218e-006, 6.097252e-009, 
    -1.65265e-006, -2.615512e-006, -4.329641e-006, -3.762904e-006, 
    -4.70292e-006, -3.27489e-006, -3.442031e-006, -3.135066e-006, 
    -1.36456e-006, -8.405354e-007, -1.271676e-006, -4.796796e-007, 
    -4.329891e-007, -1.135827e-006,
  -4.789341e-007, -8.753052e-007, -1.011651e-006, -8.04773e-007, 
    -9.408702e-007, -1.367788e-006, -1.431864e-006, -7.302669e-007, 
    -2.405157e-007, 2.102445e-007, 8.209463e-008, 4.956041e-008, 
    1.442074e-006, 2.210726e-006, 1.33255e-006, 7.563722e-008, 
    -3.191939e-006, -5.868933e-006, -2.030642e-006, -5.047629e-007, 
    9.55057e-008, 1.118471e-006, 3.572692e-006, 3.270448e-006, 1.338758e-006, 
    6.53306e-007, 2.730781e-007, 1.615423e-006, 5.619368e-006, 2.354027e-006, 
    -8.209136e-007, -1.413484e-006, -3.305682e-006, -7.044364e-007, 
    8.018178e-007, -1.011644e-006, 1.223774e-006, -1.136568e-006, 
    -1.679715e-006, -1.121152e-007, 5.616675e-007, -3.17752e-007, 
    -4.883696e-007, 3.190216e-007, 2.482411e-007, -1.618379e-006, 
    -2.028408e-006, -3.697584e-006, -5.324047e-006, -3.975491e-006, 
    -2.895655e-006, -1.789738e-006, -1.120425e-006, -1.657614e-006, 
    4.701707e-006, 6.690761e-006, 4.733991e-006, 3.307949e-006, 
    1.863527e-006, -1.237653e-006, -5.516273e-006, -9.598198e-006, 
    -9.916834e-006, -7.22469e-006, -2.308798e-006, -3.209326e-006, 
    -5.667767e-006, -6.067118e-006, -7.897481e-006, -7.272372e-006, 
    -2.079778e-007, 8.663974e-007, -2.011515e-006, -2.566834e-006, 
    3.883179e-007, 5.033035e-007, 3.831727e-006, 5.436583e-006, 
    3.082447e-006, 4.167747e-006, 3.212084e-006, 1.474111e-006, 
    5.949441e-007, -3.167615e-007, -1.722191e-006, -4.163991e-006, 
    -5.06725e-006, -4.030132e-006, -4.357212e-006, -3.791214e-006, 
    -1.240135e-006, -4.675101e-007, -3.959846e-007, -4.526087e-007, 
    3.023836e-007, 1.131411e-008,
  2.621503e-007, 4.844256e-007, -3.361313e-007, -1.131854e-006, 
    -1.456947e-006, -1.608939e-006, -1.505624e-006, -9.659534e-007, 
    -4.011999e-007, -2.35797e-007, -4.06167e-007, 1.906247e-007, 
    1.953431e-007, 2.192099e-006, 1.640508e-006, 1.409292e-006, 
    -2.232554e-006, -6.592137e-006, -6.910523e-006, -3.992131e-006, 
    -2.82239e-006, -2.955009e-006, 1.754502e-006, 1.201668e-006, 
    1.565008e-006, 8.747124e-006, -2.894412e-007, 2.18142e-006, 
    5.368036e-006, 9.428601e-006, 4.514441e-006, 7.027302e-007, 
    -3.435824e-006, -4.604815e-006, -4.648035e-006, -3.25379e-006, 
    -3.841884e-006, -5.631016e-006, -7.991606e-006, -7.847068e-006, 
    -8.607514e-006, -6.460503e-006, -5.802867e-006, -4.707632e-006, 
    -4.347274e-006, -2.925206e-006, -3.006415e-006, -5.879856e-006, 
    -5.588294e-006, -6.194767e-006, -5.897988e-006, -3.197347e-007, 
    1.384209e-006, 3.125409e-006, 1.011952e-005, 7.347902e-006, 
    5.778809e-006, 7.320585e-006, 2.742949e-006, -8.728166e-007, 
    -3.502879e-006, -4.901848e-006, -5.213034e-006, -4.637602e-006, 
    -3.961832e-006, -2.385786e-006, -4.039814e-006, -4.649522e-006, 
    -2.500278e-006, -2.585957e-006, 2.044579e-006, 2.578778e-006, 
    3.347432e-006, 3.521283e-006, 3.993906e-006, 2.928457e-006, 
    3.580139e-006, 4.738711e-006, 6.418568e-006, 3.98024e-006, 5.119187e-006, 
    3.503405e-006, 3.292551e-006, 8.775696e-007, -2.407882e-006, 
    -5.045131e-007, -4.929663e-006, -6.783614e-006, -6.705384e-006, 
    -4.933886e-006, -2.01897e-006, -1.365553e-006, -3.145249e-007, 
    -5.467346e-007, -6.788582e-007, -4.128726e-007,
  -6.709101e-007, -7.709968e-007, -2.102167e-007, -6.296846e-007, 
    -6.371342e-007, -3.160149e-006, -3.837904e-006, -3.083409e-006, 
    -3.049633e-006, -1.448503e-006, -6.664404e-007, 1.029564e-007, 
    -1.496185e-007, 1.652428e-006, 3.296771e-006, 4.55741e-006, 
    4.767019e-006, 2.514465e-006, -3.72664e-006, -4.755319e-006, 
    -3.711989e-006, -4.599602e-006, -2.167734e-006, 1.859057e-007, 
    3.80863e-007, -1.041949e-006, 5.743295e-007, 2.891211e-006, 
    3.324337e-006, 3.144783e-006, 3.534944e-006, 3.785281e-006, 
    2.124299e-006, 3.15173e-006, -5.201582e-008, 2.415363e-007, 
    -1.126893e-006, -2.005327e-007, -4.483882e-007, -1.600241e-006, 
    -4.124762e-006, -8.801988e-006, -8.669114e-006, -5.446986e-006, 
    -7.28331e-006, -7.999799e-006, -8.034567e-006, -3.559748e-006, 
    -6.035581e-006, -7.755178e-006, -6.523846e-006, -3.273897e-006, 
    -1.277142e-006, 2.895929e-006, 7.519509e-006, 7.785249e-006, 
    6.710623e-006, 6.394224e-006, 7.720182e-006, 4.245479e-006, 
    1.398119e-006, -2.418072e-006, -1.611919e-006, -1.199158e-006, 
    -2.818667e-006, -4.009267e-006, -5.134305e-006, -3.371251e-006, 
    -1.254788e-006, -3.425894e-007, 9.709511e-007, 1.802073e-008, 
    1.886368e-006, 6.986302e-006, 1.038848e-005, 8.59363e-006, 6.337359e-006, 
    4.317986e-006, 7.248302e-006, 4.607326e-006, -5.947004e-008, 
    -1.244363e-006, 2.616471e-007, -3.416459e-006, -1.72864e-006, 
    2.018023e-007, -6.601822e-006, -7.498124e-006, -4.287915e-006, 
    1.916196e-007, -8.452553e-007, -2.402428e-006, -1.559767e-006, 
    9.501036e-008, -1.4038e-006, -8.661154e-007,
  -1.758695e-006, -2.903106e-006, -3.894034e-006, -5.539618e-006, 
    -3.880374e-006, -5.905935e-006, -5.282571e-006, -3.672502e-006, 
    -6.544202e-006, -5.06427e-006, -2.573791e-006, -1.20785e-006, 
    -2.812476e-007, 2.619761e-006, 3.073998e-006, 2.736239e-006, 
    3.517059e-006, 3.409026e-006, 3.130128e-006, 2.137462e-006, 
    -3.656869e-007, -1.599801e-009, -5.772745e-008, 9.662303e-007, 
    6.28967e-007, 7.315366e-007, 3.818565e-007, 1.179814e-006, 2.042094e-006, 
    2.462803e-006, 2.367437e-006, 1.541662e-006, 1.186269e-006, 
    3.341725e-006, 3.649186e-006, 4.054993e-006, 6.419312e-006, 
    3.871701e-006, -1.467881e-006, -4.036854e-006, -7.484196e-007, 
    -1.329056e-006, -1.160923e-006, -6.701739e-007, 2.638844e-007, 
    2.616507e-007, -6.234695e-007, 2.1171e-006, 5.275157e-006, 1.428663e-006, 
    4.067166e-006, 1.575689e-006, 2.082328e-006, 3.960115e-006, 
    7.686893e-006, 1.424862e-005, 1.844032e-005, 1.257672e-005, 
    1.319238e-005, 1.173679e-005, 9.160631e-006, 8.116309e-006, 
    4.879277e-006, 3.905237e-006, 1.840435e-006, -1.131608e-006, 
    -3.226956e-006, -2.53306e-006, -1.44875e-006, 3.818559e-007, 
    1.656897e-006, 2.852965e-006, -1.763914e-006, 1.227741e-006, 
    1.096838e-005, 1.26624e-005, 9.660067e-006, 5.126887e-006, 8.491566e-006, 
    8.347517e-006, 6.429735e-006, 2.725305e-006, -3.168345e-006, 
    -3.112222e-006, -2.113593e-006, -6.354021e-007, -1.505879e-006, 
    -3.63823e-006, 9.848009e-008, 6.252671e-006, 3.709536e-006, 
    3.498686e-006, 1.501434e-006, -1.285336e-006, 7.946201e-007, 
    -5.459915e-007,
  -1.055362e-006, -3.772339e-006, -7.280569e-006, -5.962807e-006, 
    -3.390867e-006, -5.160879e-006, -2.750367e-006, 3.860787e-007, 
    -3.719935e-006, -6.602073e-006, 1.438601e-006, 1.077246e-006, 
    1.414257e-006, 2.24897e-006, 1.473366e-006, 4.265585e-007, 5.740812e-007, 
    8.701186e-007, 2.076117e-006, 2.187878e-006, 2.156584e-006, 
    1.331308e-006, 9.39408e-007, 1.146286e-006, 9.220237e-007, 1.195211e-006, 
    1.3025e-006, 5.378217e-007, 4.849226e-007, 4.322717e-007, 6.66965e-007, 
    8.206953e-007, 1.388926e-006, 2.383827e-006, 3.274916e-006, 
    3.914921e-006, 2.366196e-006, 4.926711e-006, 4.66346e-006, 2.039866e-006, 
    3.741443e-007, 7.68523e-007, 3.904221e-006, 7.905677e-006, 7.839379e-006, 
    9.252246e-006, 8.08698e-006, 7.584815e-006, 7.512295e-006, 4.806752e-006, 
    7.118666e-006, 9.381416e-006, 6.993512e-006, 7.144998e-006, 
    8.907555e-006, 1.762e-005, 2.075719e-005, 1.997167e-005, 1.708581e-005, 
    1.434026e-005, 1.164341e-005, 9.748223e-006, 9.541589e-006, 
    3.749021e-006, 5.821275e-006, 2.856443e-006, 2.976649e-007, 
    1.327571e-007, 1.846392e-006, 1.423448e-006, 2.782929e-006, 6.30333e-006, 
    6.288434e-006, 2.722829e-006, 4.867845e-006, 8.584691e-006, 
    1.039022e-005, 8.280967e-006, 4.62e-006, 5.626571e-006, 8.351475e-006, 
    4.873305e-006, 1.982495e-006, 1.975786e-006, 5.576294e-008, 
    -1.469372e-006, -2.022716e-008, -3.362056e-006, -2.312285e-006, 
    5.482274e-006, 8.068375e-006, 8.192546e-006, 6.558392e-006, 
    6.778928e-006, 6.29414e-006, 3.89158e-006,
  6.618988e-006, 1.398114e-006, 1.587856e-006, 3.327321e-006, 2.524896e-006, 
    2.134979e-006, 1.606983e-006, 2.555189e-006, 1.185773e-006, 
    1.430653e-006, 4.966447e-006, 5.409262e-006, 1.374026e-006, 
    9.004161e-007, 1.316655e-006, 1.539181e-006, 1.319636e-006, 
    2.233823e-006, 2.913813e-006, 3.165889e-006, 3.115722e-006, 
    1.489261e-006, 1.034279e-006, 8.333616e-007, 4.975885e-007, 
    4.066915e-007, 5.32855e-007, 5.363316e-007, 2.966711e-007, 1.829256e-007, 
    3.493222e-007, 4.789624e-007, 6.818663e-007, 1.11996e-006, 1.946727e-006, 
    3.176073e-006, 2.848246e-006, 4.524125e-006, 5.169593e-006, 
    4.649799e-006, 7.20832e-006, 6.13743e-006, 5.409504e-006, 4.86214e-006, 
    8.172188e-006, 1.032912e-005, 1.081888e-005, 1.086706e-005, 
    1.041034e-005, 1.025238e-005, 8.312505e-006, 8.339332e-006, 
    8.864838e-006, 9.905685e-006, 1.425434e-005, 1.252829e-005, 
    9.789212e-006, 9.547799e-006, 1.243813e-005, 1.343626e-005, 
    1.416642e-005, 1.359918e-005, 1.296191e-005, 9.453441e-006, 
    4.914291e-006, 3.076231e-006, 1.979761e-006, 1.064576e-006, 
    2.595671e-006, 1.657892e-006, 1.626599e-006, 3.605723e-006, 
    3.959128e-006, 3.551088e-006, 6.178159e-006, 5.969045e-006, 
    7.059563e-006, 6.246952e-006, 3.792975e-006, 4.981099e-006, 
    5.194186e-006, 3.640744e-006, 3.926845e-006, 4.880763e-006, 
    2.169003e-006, 3.277892e-006, 3.508103e-007, -2.444722e-008, 
    2.496745e-008, 3.629557e-006, 1.241405e-005, 1.257746e-005, 
    1.184955e-005, 1.429333e-005, 1.915012e-005, 1.227919e-005,
  8.763764e-006, 7.373237e-006, 1.140151e-005, 9.914129e-006, 4.940868e-006, 
    3.550096e-006, 2.961247e-006, 1.536694e-006, 1.45896e-006, 3.642726e-006, 
    5.413728e-006, 4.941609e-006, 5.163388e-006, 3.546862e-006, 
    1.924124e-006, 1.610458e-006, 1.993417e-006, 2.314538e-006, 
    1.879672e-006, 1.821308e-006, 2.597659e-006, 2.48441e-006, 1.055141e-006, 
    8.355964e-007, 9.533155e-007, 1.140574e-006, 1.11251e-006, 3.649682e-007, 
    3.244867e-007, 7.476798e-007, 9.063773e-007, 6.503257e-007, 
    4.702698e-007, 7.769852e-007, 1.372287e-006, 1.025089e-006, 
    8.447864e-007, 9.426367e-007, 4.595415e-006, 7.903718e-006, 
    7.109978e-006, 8.493549e-006, 7.612645e-006, 3.766159e-006, 
    5.269929e-006, 9.436546e-006, 1.042275e-005, 9.547308e-006, 
    8.213407e-006, 8.392966e-006, 6.855909e-006, 1.315737e-005, 
    1.444955e-005, 1.095571e-005, 1.02889e-005, 1.338287e-005, 1.16598e-005, 
    1.053376e-005, 1.227199e-005, 1.358577e-005, 8.75456e-006, 8.570787e-006, 
    6.749364e-006, 4.623718e-006, 5.842132e-006, 5.270678e-006, 
    2.621005e-006, 1.560289e-006, 1.605737e-006, 1.557061e-006, 
    1.639763e-006, 2.294667e-006, 1.356639e-006, 2.384328e-006, 
    3.424677e-006, 5.520029e-006, 5.288068e-006, 1.041705e-005, 
    9.721654e-006, 8.816412e-006, 8.186085e-006, 5.222006e-006, 6.60359e-006, 
    1.976285e-006, 2.298395e-006, 2.538796e-006, 1.541659e-006, 
    -1.240634e-006, -2.127501e-006, 1.105553e-006, 7.18547e-006, 
    1.001445e-005, 9.719166e-006, 1.206412e-005, 1.34842e-005, 1.10558e-005,
  4.779688e-006, 6.265083e-006, 8.773446e-006, 7.197648e-006, 3.577163e-006, 
    3.7674e-006, 3.752996e-006, 2.304105e-006, 2.605356e-006, 2.908595e-006, 
    3.288575e-006, 4.942852e-006, 4.32346e-006, 3.515073e-006, 4.137692e-006, 
    3.824272e-006, 2.175956e-006, 2.045075e-006, 2.245495e-006, 
    1.756985e-006, 1.205146e-006, 1.311937e-006, 2.59915e-006, 1.883398e-006, 
    1.225759e-006, 1.32808e-006, 1.390416e-006, 1.450269e-006, 1.289834e-006, 
    9.729355e-007, 7.551304e-007, 8.778163e-007, 1.051664e-006, 
    7.419677e-007, 7.278113e-007, 3.470866e-007, 2.19185e-007, 4.499061e-007, 
    2.877304e-006, 4.703445e-006, 3.453486e-006, 2.554447e-006, 
    5.401807e-006, 7.320832e-006, 3.981979e-006, 4.043319e-006, 
    6.051501e-006, 7.141516e-006, 5.340469e-006, 8.678824e-006, 
    9.308395e-006, 1.006115e-005, 1.143703e-005, 9.60493e-006, 9.336705e-006, 
    8.964918e-006, 1.084097e-005, 8.584444e-006, 7.339946e-006, 
    5.629543e-006, 3.91938e-006, 2.93069e-006, 1.716005e-006, -7.441849e-007, 
    1.154476e-006, 1.697133e-006, 4.563608e-007, 9.652349e-007, 
    6.336868e-007, 1.390169e-006, 3.000486e-006, 2.5912e-006, 2.579776e-006, 
    2.682345e-006, 2.031414e-006, 3.742813e-006, 5.981467e-006, 
    7.219258e-006, 7.198149e-006, 6.304575e-006, 6.953269e-006, 
    5.658607e-006, 2.583747e-006, 2.8701e-006, 3.060337e-006, 2.598645e-006, 
    -2.997982e-006, -6.677328e-006, -1.92659e-006, -1.723689e-006, 
    2.252189e-006, 3.891317e-006, 7.877628e-006, 7.545335e-006, 
    8.819388e-006, 8.138159e-006,
  4.347305e-006, 3.956648e-006, 4.421068e-006, 4.631666e-006, 5.442043e-006, 
    4.281988e-006, 2.696751e-006, 2.72233e-006, 3.52277e-006, 1.749037e-006, 
    2.206253e-006, 2.906359e-006, 3.233192e-006, 2.923248e-006, 
    3.851093e-006, 4.33116e-006, 2.260395e-006, 1.387685e-006, 1.532971e-006, 
    1.283874e-006, 9.679684e-007, 1.244137e-006, 2.560158e-006, 
    2.327698e-006, 2.405681e-006, 2.86886e-006, 2.918282e-006, 2.50552e-006, 
    2.405682e-006, 1.825779e-006, 1.395384e-006, 1.40805e-006, 1.08842e-006, 
    9.096057e-007, 7.116691e-007, 8.788097e-007, 1.355896e-006, 
    2.665708e-006, 4.945336e-006, 9.877623e-006, 9.126108e-006, 
    6.786413e-007, 1.254568e-006, 4.543006e-006, 5.26795e-006, 5.510832e-006, 
    2.731276e-006, 1.012426e-006, 1.228742e-006, 2.24599e-006, 4.259389e-006, 
    4.01302e-006, 6.673627e-006, 9.899477e-006, 8.942081e-006, 6.185113e-006, 
    6.086269e-006, 6.487109e-006, 5.93378e-006, 4.594411e-006, 4.360212e-006, 
    4.260633e-006, 5.568952e-006, 4.443158e-006, 1.90277e-006, 1.877932e-006, 
    2.285478e-006, 1.829998e-006, 1.689929e-006, 1.761456e-006, 
    1.598536e-006, 2.724318e-006, 3.506381e-006, 3.575671e-006, 
    4.982589e-006, 7.164118e-006, 7.29227e-006, 6.751856e-006, 6.403168e-006, 
    7.115443e-006, 7.708511e-006, 7.594268e-006, 3.870466e-006, 
    2.139193e-006, 3.216552e-006, 1.544144e-006, -2.253422e-006, 
    -4.059195e-006, -2.381323e-006, -1.907218e-006, -2.659232e-006, 
    1.975775e-006, 5.021822e-006, 5.652397e-006, 5.944457e-006, 5.404045e-006,
  3.350418e-006, 1.946228e-006, 3.019115e-006, 5.584845e-006, 7.065282e-006, 
    4.490108e-006, 5.959346e-007, 4.794574e-007, 2.338382e-006, 
    1.317401e-006, 1.925118e-006, 2.728042e-006, 2.928711e-006, 
    1.890349e-006, 2.235559e-006, 3.345447e-006, 2.605855e-006, 
    1.133124e-006, 8.346033e-007, 1.183539e-006, 1.281142e-006, 
    1.056383e-006, 1.017392e-006, 5.867473e-007, 1.090408e-006, 
    2.260395e-006, 2.481677e-006, 1.722464e-006, 1.813113e-006, 
    2.477704e-006, 2.323477e-006, 1.13362e-006, 7.362555e-007, 1.254319e-006, 
    1.624613e-006, 1.189002e-006, 1.542408e-006, 2.824653e-006, 
    5.566465e-006, 6.924955e-006, 4.148372e-006, 1.353907e-006, 
    1.203903e-006, 1.47113e-006, 1.102082e-006, 6.371738e-008, 1.472126e-006, 
    1.828266e-006, 4.118325e-006, 3.912688e-006, 4.047793e-006, 
    6.127251e-006, 7.868452e-006, 7.500394e-006, 6.989283e-006, 7.34095e-006, 
    1.003706e-005, 1.051439e-005, 6.11756e-006, 6.056714e-006, 9.75791e-006, 
    1.255536e-005, 9.938969e-006, 6.26608e-006, 3.490488e-006, 2.245245e-006, 
    2.30361e-006, 3.045686e-006, 5.236407e-006, 4.202265e-006, 4.057475e-006, 
    4.194318e-006, 5.016613e-006, 5.496927e-006, 7.212548e-006, 
    7.738807e-006, 6.508965e-006, 5.030273e-006, 3.353892e-006, 3.40083e-006, 
    5.383929e-006, 6.871067e-006, 5.440805e-006, 4.302605e-006, 5.12937e-006, 
    4.568341e-006, 1.861052e-006, 2.618981e-007, -1.809363e-006, 
    -1.759199e-006, 5.306138e-007, 2.368175e-006, 3.352892e-006, 
    2.587476e-006, 4.302352e-006, 2.973666e-006,
  1.101653e-007, -1.359344e-006, -1.983202e-006, 1.576187e-006, 
    3.354146e-006, 2.284985e-006, 2.015022e-006, 2.139198e-006, 
    1.359867e-006, 1.140076e-006, 1.440582e-006, 2.608833e-006, 
    2.691782e-006, 2.218423e-006, 1.366573e-006, 1.55731e-006, 2.426294e-006, 
    1.653172e-006, 7.196168e-007, 3.7987e-007, 1.037012e-006, 1.554827e-006, 
    1.766671e-006, 1.046447e-006, 7.434573e-007, 1.185525e-006, 
    1.738607e-006, 1.296043e-006, 1.048435e-006, 1.476595e-006, 
    1.206635e-006, 1.165161e-006, 1.133371e-006, 1.268972e-006, 
    1.475353e-006, 2.912075e-007, -5.325546e-009, 4.643093e-007, 
    1.574694e-006, 1.316656e-006, 1.346707e-006, 1.078486e-006, 4.21097e-007, 
    1.338012e-006, 9.769083e-007, 1.430152e-006, 2.271821e-006, 
    3.867239e-006, 4.645082e-006, 5.733611e-006, 6.738198e-006, 
    6.580742e-006, 5.483269e-006, 5.501895e-006, 7.931284e-006, 
    1.061722e-005, 1.462315e-005, 1.328055e-005, 1.102874e-005, 
    1.053328e-005, 1.071507e-005, 8.885951e-006, 6.18561e-006, 4.394986e-006, 
    3.457702e-006, 2.168505e-006, 2.149879e-006, 2.917041e-006, 
    3.560025e-006, 3.818809e-006, 4.076351e-006, 3.938266e-006, 3.71003e-006, 
    4.276027e-006, 4.608322e-006, 4.041581e-006, 3.60299e-006, 4.034876e-006, 
    3.31217e-006, 3.178555e-006, 3.477324e-006, 4.292914e-006, 3.208854e-006, 
    4.53655e-006, 7.834176e-006, 9.473304e-006, 5.857783e-006, 
    -3.356363e-007, -2.864363e-006, 4.320173e-007, 1.66037e-006, 
    -2.72107e-006, -6.582952e-006, -5.126116e-006, -1.714739e-006, 
    -1.575972e-008,
  -7.100265e-006, -7.366496e-006, -4.975107e-006, -1.642218e-006, 
    4.243229e-007, 1.121697e-006, 1.443563e-006, 1.241155e-006, 
    1.404075e-006, 5.552047e-007, -3.31429e-008, 1.45671e-007, 3.095847e-007, 
    9.699397e-008, 2.15211e-007, 2.628949e-007, 3.979985e-007, 1.176335e-006, 
    1.58711e-006, 1.678258e-006, 1.084943e-006, 4.538779e-007, 8.567067e-007, 
    9.823734e-007, 7.352628e-007, 1.170377e-006, 1.075754e-006, 
    8.544712e-007, 9.267419e-007, 1.001993e-006, 1.221785e-006, 
    8.010754e-007, 2.472484e-007, -1.600256e-009, 2.56935e-007, 
    3.756472e-007, 5.53468e-007, 8.375832e-007, 1.180061e-006, 1.745561e-006, 
    1.968334e-006, 1.818079e-006, 1.29356e-006, 1.188754e-006, 1.20912e-006, 
    1.442322e-006, 2.388048e-006, 3.173339e-006, 3.789502e-006, 
    4.132725e-006, 4.235048e-006, 4.666436e-006, 4.714615e-006, 
    4.328677e-006, 5.293527e-006, 7.034479e-006, 7.007658e-006, 
    4.703193e-006, 3.863513e-006, 4.344571e-006, 4.237034e-006, 
    3.679979e-006, 3.109265e-006, 3.058602e-006, 2.865632e-006, 
    2.101948e-006, 2.38954e-006, 2.299883e-006, 1.917918e-006, 2.401212e-006, 
    2.484659e-006, 2.777715e-006, 3.086665e-006, 3.511348e-006, 
    3.522028e-006, 2.73326e-006, 1.921891e-006, 2.136716e-006, 2.656271e-006, 
    2.411394e-006, 1.990436e-006, 2.195326e-006, 2.153106e-006, 
    2.654779e-006, 3.813846e-006, 5.090134e-006, 6.025173e-006, 
    4.313526e-006, 2.609577e-006, -1.227472e-006, -3.815061e-006, 
    -4.599347e-006, -4.141884e-006, -5.482992e-006, -4.71384e-006, 
    -4.577001e-006,
  -5.581091e-006, -7.4564e-006, -9.564916e-006, -9.039155e-006, 
    -6.040545e-006, -3.225468e-006, -1.736594e-006, -7.002182e-007, 
    6.605069e-007, 1.264997e-006, 1.763689e-006, 2.588717e-006, 
    2.709913e-006, 1.379736e-006, 5.234169e-007, 2.549486e-007, 
    -3.917617e-007, -3.194914e-007, 1.551107e-007, 1.317153e-006, 
    2.178192e-006, 2.166519e-006, 1.754502e-006, 1.197445e-006, 6.77147e-007, 
    5.368283e-007, 4.387293e-007, 6.77644e-007, 7.037211e-007, 6.513185e-007, 
    6.843493e-007, 6.8435e-007, 7.245831e-007, 1.129149e-006, 1.272946e-006, 
    1.282135e-006, 1.743823e-006, 1.948217e-006, 2.184897e-006, 
    2.167512e-006, 1.745064e-006, 1.684466e-006, 1.852849e-006, 
    1.602759e-006, 9.860992e-007, 1.336029e-006, 2.272566e-006, 
    3.317882e-006, 3.380963e-006, 3.239899e-006, 2.839306e-006, 
    2.607594e-006, 3.203887e-006, 3.44926e-006, 3.428647e-006, 3.597278e-006, 
    3.47509e-006, 2.395251e-006, 2.553701e-006, 2.494344e-006, 2.861658e-006, 
    3.030787e-006, 2.595672e-006, 2.368926e-006, 1.984973e-006, 
    1.770396e-006, 1.709798e-006, 1.642246e-006, 1.807897e-006, 
    2.064197e-006, 2.076118e-006, 2.05476e-006, 2.334653e-006, 2.218424e-006, 
    1.992424e-006, 1.793245e-006, 2.018501e-006, 2.551465e-006, 
    2.643356e-006, 2.507507e-006, 2.077112e-006, 1.71849e-006, 1.019875e-006, 
    1.314669e-006, 1.897303e-006, 3.06158e-006, 4.964957e-006, 5.770862e-006, 
    6.290416e-006, 5.786012e-006, 3.049914e-006, -3.438254e-007, 
    -1.483519e-006, -2.483386e-006, -3.564715e-006, -3.583591e-006,
  -3.303945e-006, -3.297488e-006, -4.288411e-006, -5.987145e-006, 
    -7.162598e-006, -5.869928e-006, -3.154439e-006, -1.25429e-006, 
    6.848441e-007, 2.12529e-006, 2.598898e-006, 2.829867e-006, 2.679365e-006, 
    2.645589e-006, 2.118833e-006, 7.769859e-007, 4.158805e-007, 
    8.087745e-007, 1.005221e-006, 1.000999e-006, 1.364091e-006, 
    1.304983e-006, 9.831183e-007, 1.02211e-006, 1.245379e-006, 1.325845e-006, 
    1.583884e-006, 1.552591e-006, 7.971023e-007, 7.60346e-007, 8.544714e-007, 
    1.014907e-006, 8.390739e-007, 8.306301e-007, 1.021861e-006, 
    1.229236e-006, 1.417487e-006, 1.321374e-006, 1.082956e-006, 
    8.748366e-007, 7.610902e-007, 7.891547e-007, 1.189499e-006, 
    1.357138e-006, 1.312186e-006, 1.28735e-006, 1.66584e-006, 2.178192e-006, 
    2.107659e-006, 2.036878e-006, 1.797715e-006, 1.377751e-006, 
    1.184284e-006, 1.304487e-006, 1.440584e-006, 1.957903e-006, 
    2.161303e-006, 2.031167e-006, 2.036879e-006, 1.743574e-006, 
    1.800447e-006, 1.632064e-006, 1.810878e-006, 2.358744e-006, 
    2.331176e-006, 2.070406e-006, 2.01403e-006, 1.84366e-006, 1.486777e-006, 
    1.646717e-006, 1.859804e-006, 1.802434e-006, 1.47138e-006, 1.596301e-006, 
    1.980503e-006, 2.053767e-006, 2.222647e-006, 2.255181e-006, 
    1.864274e-006, 1.407056e-006, 1.197447e-006, 9.843598e-007, 
    1.065323e-006, 1.292317e-006, 1.32957e-006, 1.111268e-006, 1.335282e-006, 
    2.607841e-006, 5.20387e-006, 6.569562e-006, 4.793842e-006, 2.591201e-006, 
    1.255066e-006, -4.59313e-007, -2.690263e-006, -3.488223e-006,
  -2.261111e-006, -2.441167e-006, -2.301844e-006, -2.161772e-006, 
    -2.234043e-006, -1.923354e-006, -1.149239e-006, -5.608917e-007, 
    -3.095593e-007, -1.059097e-007, 3.473342e-007, 8.403149e-007, 
    1.10183e-006, 1.351426e-006, 1.589844e-006, 1.698126e-006, 1.506397e-006, 
    1.535703e-006, 1.402834e-006, 1.17435e-006, 1.124928e-006, 1.123189e-006, 
    9.649884e-007, 7.295503e-007, 7.11917e-007, 8.87751e-007, 7.876647e-007, 
    5.994125e-007, 5.462659e-007, 5.65389e-007, 6.721805e-007, 8.057943e-007, 
    9.600215e-007, 8.966915e-007, 9.577861e-007, 1.133868e-006, 
    1.172114e-006, 1.177827e-006, 1.097609e-006, 1.062094e-006, 
    1.153736e-006, 1.18329e-006, 1.296291e-006, 1.444557e-006, 1.244634e-006, 
    1.142313e-006, 1.143554e-006, 1.147279e-006, 1.38545e-006, 1.625606e-006, 
    1.729418e-006, 1.707066e-006, 1.494974e-006, 1.301507e-006, 
    1.322368e-006, 1.515338e-006, 1.328329e-006, 1.043717e-006, 
    9.560474e-007, 9.736802e-007, 1.161187e-006, 1.286605e-006, 1.47734e-006, 
    1.538187e-006, 1.609215e-006, 1.544395e-006, 1.578171e-006, 
    1.475104e-006, 1.338263e-006, 1.27071e-006, 1.164913e-006, 1.149763e-006, 
    1.185029e-006, 1.204152e-006, 1.079728e-006, 1.004973e-006, 8.9992e-007, 
    7.57117e-007, 6.657235e-007, 6.356724e-007, 9.875889e-007, 1.156965e-006, 
    1.118719e-006, 9.848566e-007, 8.028139e-007, 8.154801e-007, 
    1.249104e-006, 2.103685e-006, 3.020853e-006, 2.973666e-006, 1.81212e-006, 
    6.905584e-007, 3.967561e-007, 6.629907e-007, 1.372282e-007, -1.547596e-006,
  5.11247e-007, 1.407043e-007, -5.823495e-009, 5.601669e-008, 1.464177e-007, 
    5.974289e-008, 7.017388e-008, 2.54453e-007, 5.825259e-007, 1.004725e-006, 
    1.284867e-006, 1.415252e-006, 1.465917e-006, 1.513352e-006, 
    1.431396e-006, 1.226752e-006, 1.072029e-006, 1.032044e-006, 
    9.813798e-007, 9.903206e-007, 1.111268e-006, 1.144051e-006, 
    1.127908e-006, 1.128653e-006, 1.167892e-006, 1.316159e-006, 
    1.456975e-006, 1.43512e-006, 1.235445e-006, 1.132875e-006, 1.146038e-006, 
    1.122196e-006, 1.195956e-006, 1.27096e-006, 1.190245e-006, 1.052409e-006, 
    9.543089e-007, 9.540609e-007, 9.987641e-007, 1.028318e-006, 
    1.057624e-006, 1.058866e-006, 1.017391e-006, 1.036265e-006, 1.16069e-006, 
    1.345217e-006, 1.440087e-006, 1.369803e-006, 1.404324e-006, 
    1.568237e-006, 1.623123e-006, 1.60698e-006, 1.58438e-006, 1.583138e-006, 
    1.610209e-006, 1.592079e-006, 1.562028e-006, 1.629331e-006, 
    1.759469e-006, 1.715262e-006, 1.487025e-006, 1.366078e-006, 
    1.432885e-006, 1.561283e-006, 1.66112e-006, 1.705824e-006, 1.636534e-006, 
    1.492738e-006, 1.402586e-006, 1.361856e-006, 1.398861e-006, 
    1.437852e-006, 1.361111e-006, 1.116732e-006, 9.210298e-007, 
    8.907309e-007, 9.942937e-007, 1.144796e-006, 1.334537e-006, 
    1.341243e-006, 1.17286e-006, 1.032789e-006, 8.075326e-007, 5.261492e-007, 
    3.331791e-007, 4.402191e-007, 1.103817e-006, 2.145657e-006, 
    2.998749e-006, 3.255297e-006, 2.885997e-006, 2.120575e-006, 
    1.255561e-006, 6.458549e-007, 5.502388e-007, 6.331875e-007,
  1.803676e-006, 1.535951e-006, 1.292566e-006, 1.066068e-006, 8.298848e-007, 
    5.765651e-007, 3.696869e-007, 2.805282e-007, 3.152977e-007, 
    4.186127e-007, 5.422926e-007, 6.692007e-007, 8.365905e-007, 
    9.826213e-007, 1.04918e-006, 1.077989e-006, 1.082708e-006, 1.048932e-006, 
    9.697069e-007, 8.698694e-007, 8.020688e-007, 8.311263e-007, 
    9.125856e-007, 9.977707e-007, 9.952878e-007, 9.108473e-007, 
    7.956112e-007, 7.183737e-007, 7.253279e-007, 7.710248e-007, 
    8.055463e-007, 8.507461e-007, 9.110959e-007, 9.600215e-007, 
    1.014907e-006, 1.098105e-006, 1.191486e-006, 1.302996e-006, 
    1.376757e-006, 1.375267e-006, 1.339256e-006, 1.278409e-006, 
    1.257796e-006, 1.289337e-006, 1.346955e-006, 1.401592e-006, 1.38992e-006, 
    1.306224e-006, 1.200178e-006, 1.082211e-006, 9.885816e-007, 
    1.016149e-006, 1.153737e-006, 1.311937e-006, 1.456975e-006, 
    1.575687e-006, 1.660624e-006, 1.742084e-006, 1.755743e-006, 
    1.712033e-006, 1.664349e-006, 1.65516e-006, 1.711785e-006, 1.809387e-006, 
    1.93108e-006, 1.983979e-006, 1.895814e-006, 1.746802e-006, 1.594066e-006, 
    1.479078e-006, 1.373032e-006, 1.264253e-006, 1.182794e-006, 
    1.152743e-006, 1.147527e-006, 1.137593e-006, 1.113006e-006, 
    1.052657e-006, 9.597729e-007, 8.932143e-007, 8.924692e-007, 
    9.178013e-007, 9.292253e-007, 9.51329e-007, 9.317089e-007, 8.624188e-007, 
    7.685412e-007, 7.111719e-007, 7.705275e-007, 9.461137e-007, 
    1.218308e-006, 1.556565e-006, 1.913945e-006, 2.165526e-006, 
    2.179434e-006, 2.03514e-006,
  2.287218e-006, 2.171982e-006, 2.058237e-006, 1.959144e-006, 1.881162e-006, 
    1.825034e-006, 1.773128e-006, 1.722464e-006, 1.67478e-006, 1.625855e-006, 
    1.575191e-006, 1.518318e-006, 1.454988e-006, 1.389423e-006, 
    1.331557e-006, 1.280645e-006, 1.230974e-006, 1.182545e-006, 
    1.144299e-006, 1.120953e-006, 1.113999e-006, 1.123685e-006, 
    1.150756e-006, 1.191734e-006, 1.230477e-006, 1.262763e-006, 
    1.290331e-006, 1.314669e-006, 1.332302e-006, 1.330067e-006, 
    1.313427e-006, 1.283873e-006, 1.242647e-006, 1.19844e-006, 1.151501e-006, 
    1.104563e-006, 1.06582e-006, 1.040984e-006, 1.032044e-006, 1.039743e-006, 
    1.064081e-006, 1.101582e-006, 1.153488e-006, 1.203903e-006, 1.24811e-006, 
    1.281141e-006, 1.302251e-006, 1.321374e-006, 1.342484e-006, 
    1.365084e-006, 1.388429e-006, 1.413017e-006, 1.443564e-006, 
    1.479327e-006, 1.519063e-006, 1.554329e-006, 1.59183e-006, 1.624613e-006, 
    1.645475e-006, 1.649697e-006, 1.637279e-006, 1.616169e-006, 
    1.589844e-006, 1.56178e-006, 1.54514e-006, 1.534461e-006, 1.523286e-006, 
    1.508136e-006, 1.489758e-006, 1.480817e-006, 1.48032e-006, 1.499195e-006, 
    1.537442e-006, 1.594563e-006, 1.657893e-006, 1.709302e-006, 
    1.748293e-006, 1.768161e-006, 1.7699e-006, 1.7622e-006, 1.752018e-006, 
    1.745313e-006, 1.744319e-006, 1.761456e-006, 1.799205e-006, 
    1.865516e-006, 1.957654e-006, 2.071896e-006, 2.194831e-006, 
    2.308576e-006, 2.403944e-006, 2.477208e-006, 2.516696e-006, 
    2.516945e-006, 2.474725e-006, 2.392768e-006,
  4.246988e-007, 4.934925e-007, 5.478819e-007, 5.84638e-007, 6.097216e-007, 
    6.199041e-007, 6.15682e-007, 6.010293e-007, 5.853831e-007, 5.784291e-007, 
    5.794227e-007, 5.891081e-007, 5.960621e-007, 5.948204e-007, 
    5.764423e-007, 5.391894e-007, 4.86787e-007, 4.254439e-007, 3.690677e-007, 
    3.226257e-007, 2.9034e-007, 2.781708e-007, 2.784191e-007, 2.945621e-007, 
    3.251096e-007, 3.670807e-007, 4.135227e-007, 4.607098e-007, 
    5.118704e-007, 5.607958e-007, 6.050025e-007, 6.420071e-007, 
    6.742932e-007, 7.058338e-007, 7.346425e-007, 7.666802e-007, 
    8.133704e-007, 8.767011e-007, 9.70578e-007, 1.101708e-006, 1.267359e-006, 
    1.458342e-006, 1.67118e-006, 1.901652e-006, 2.150253e-006, 2.408291e-006, 
    2.669558e-006, 2.922879e-006, 3.146644e-006, 3.332661e-006, 
    3.477202e-006, 3.572073e-006, 3.617025e-006, 3.613548e-006, 3.56487e-006, 
    3.468758e-006, 3.336882e-006, 3.179924e-006, 3.006076e-006, 2.81857e-006, 
    2.626842e-006, 2.435113e-006, 2.255058e-006, 2.09338e-006, 1.945611e-006, 
    1.809513e-006, 1.679376e-006, 1.546756e-006, 1.411156e-006, 1.27034e-006, 
    1.117106e-006, 9.489715e-007, 7.805882e-007, 6.295897e-007, 5.03923e-007, 
    4.045821e-007, 3.338016e-007, 2.987838e-007, 2.928234e-007, 
    3.010189e-007, 3.042476e-007, 3.007706e-007, 2.915815e-007, 
    2.732036e-007, 2.434012e-007, 2.118604e-007, 1.746075e-007, 1.34871e-007, 
    1.025851e-007, 8.669053e-008, 8.917414e-008, 1.070555e-007, 
    1.448052e-007, 2.021748e-007, 2.739489e-007, 3.516832e-007,
  5.198181e-007, 5.545864e-007, 5.473848e-007, 5.250336e-007, 5.006948e-007, 
    4.924991e-007, 5.086422e-007, 5.324839e-007, 5.036752e-007, 
    4.249467e-007, 3.365335e-007, 3.151754e-007, 3.564019e-007, 
    4.192352e-007, 4.912577e-007, 5.560777e-007, 6.037615e-007, 
    6.427526e-007, 6.643592e-007, 6.745418e-007, 6.708162e-007, 
    6.457327e-007, 6.054994e-007, 5.714753e-007, 5.431632e-007, 
    4.962245e-007, 4.110395e-007, 3.107053e-007, 2.441466e-007, 
    2.478719e-007, 3.288346e-007, 4.44567e-007, 5.339742e-007, 5.948206e-007, 
    6.439941e-007, 7.465636e-007, 9.392857e-007, 1.182671e-006, 
    1.357263e-006, 1.399235e-006, 1.350309e-006, 1.330689e-006, 
    1.385824e-006, 1.505778e-006, 1.721347e-006, 2.082204e-006, 
    2.629325e-006, 3.318753e-006, 3.996758e-006, 4.513827e-006, 
    4.797445e-006, 4.914171e-006, 4.823522e-006, 4.518794e-006, 4.03674e-006, 
    3.433989e-006, 2.829996e-006, 2.327331e-006, 1.939155e-006, 
    1.555202e-006, 1.254944e-006, 1.125552e-006, 1.0503e-006, 1.045581e-006, 
    1.150385e-006, 1.283999e-006, 1.360491e-006, 1.393771e-006, 
    1.460577e-006, 1.525646e-006, 1.531855e-006, 1.570101e-006, 1.72259e-006, 
    1.941637e-006, 2.070532e-006, 1.994784e-006, 1.687572e-006, 
    1.259661e-006, 8.245465e-007, 5.208117e-007, 3.722967e-007, 
    2.920788e-007, 2.068937e-007, 8.470397e-008, -1.353369e-007, 
    -3.772329e-007, -5.406487e-007, -6.114287e-007, -6.111804e-007, 
    -5.923057e-007, -5.33943e-007, -4.15479e-007, -2.088491e-007, 
    3.801415e-008, 2.719621e-007, 4.393514e-007,
  5.568222e-007, 3.360365e-007, 1.840449e-007, 3.621137e-007, 7.666804e-007, 
    1.145667e-006, 1.319265e-006, 1.290705e-006, 1.207258e-006, 1.0878e-006, 
    8.886215e-007, 7.021085e-007, 6.606339e-007, 5.943239e-007, 
    4.197318e-007, 3.156722e-007, 3.357887e-007, 4.09798e-007, 4.19732e-007, 
    3.119471e-007, 2.982877e-007, 3.631077e-007, 4.21222e-007, 4.470508e-007, 
    4.813235e-007, 4.885255e-007, 4.117848e-007, 2.627729e-007, 
    2.890985e-007, 4.487893e-007, 4.723828e-007, 3.501933e-007, 3.10457e-007, 
    4.142684e-007, 5.516072e-007, 6.991282e-007, 7.567461e-007, 
    7.430867e-007, 8.734717e-007, 1.070664e-006, 1.349564e-006, 
    1.653796e-006, 1.840557e-006, 1.834846e-006, 1.711662e-006, 
    1.906619e-006, 2.396619e-006, 2.954421e-006, 3.362465e-006, 
    3.856685e-006, 4.478561e-006, 4.797445e-006, 4.491226e-006, 
    3.800806e-006, 3.026692e-006, 2.102571e-006, 1.226879e-006, 
    5.297525e-007, -1.092585e-007, -5.731818e-007, -8.307234e-007, 
    -9.553969e-007, -8.965362e-007, -7.293957e-007, -4.745871e-007, 
    -1.927065e-007, -1.97133e-009, 3.601267e-007, 1.087055e-006, 
    1.853968e-006, 2.282874e-006, 2.436107e-006, 2.552584e-006, 2.51558e-006, 
    2.338008e-006, 2.275423e-006, 2.37526e-006, 2.49447e-006, 2.860542e-006, 
    3.189858e-006, 3.091759e-006, 2.377e-006, 1.608348e-006, 1.071409e-006, 
    8.235529e-007, 6.136952e-007, 3.285877e-007, -8.427378e-009, 
    -4.164713e-007, -6.630853e-007, -4.745862e-007, -1.27141e-007, 
    1.88516e-007, 4.527624e-007, 6.579021e-007, 7.252056e-007,
  2.689819e-007, 2.72707e-007, 3.241162e-007, 5.091388e-007, 8.404411e-007, 
    1.05626e-006, 1.103695e-006, 1.001125e-006, 1.023974e-006, 1.1104e-006, 
    8.401928e-007, 6.509481e-007, 5.208115e-007, 3.092148e-007, 
    2.158343e-007, 2.011817e-007, 2.369445e-007, 2.669951e-007, 
    3.578921e-007, 3.668328e-007, 1.085459e-007, -1.70106e-007, 
    -2.043785e-007, 3.925516e-008, 1.982014e-007, 3.606237e-007, 
    4.895189e-007, 5.893567e-007, 6.723064e-007, 6.713128e-007, 
    4.957276e-007, 4.517694e-007, 4.947342e-007, 3.531734e-007, 
    6.011715e-008, -1.929545e-007, -1.333499e-007, 2.436495e-007, 
    6.534317e-007, 1.133497e-006, 1.27034e-006, 1.316781e-006, 1.21297e-006, 
    5.920883e-007, 2.01429e-007, 6.91678e-007, 1.012302e-006, 7.915178e-007, 
    8.454099e-007, 8.747156e-007, 1.081594e-006, 1.394518e-006, 1.85869e-006, 
    2.329317e-006, 2.544639e-006, 2.184775e-006, 1.363224e-006, 
    2.652569e-007, -1.162026e-006, -2.496923e-006, -3.195043e-006, 
    -2.77135e-006, -1.698962e-006, -8.811367e-007, -4.485082e-007, 
    3.268506e-007, 1.746185e-006, 2.731153e-006, 3.074872e-006, 
    3.858425e-006, 4.554558e-006, 4.281121e-006, 3.613301e-006, 
    2.794482e-006, 2.291318e-006, 2.175089e-006, 2.13138e-006, 2.021361e-006, 
    1.581529e-006, 1.291452e-006, 1.561411e-006, 1.804549e-006, 
    1.353788e-006, 1.137225e-006, 1.344101e-006, 1.312809e-006, 
    8.235538e-007, -1.956869e-007, -1.235789e-006, -1.808986e-006, 
    -1.195803e-006, 3.601281e-007, 1.832859e-006, 2.056873e-006, 
    1.244014e-006, 5.79174e-007,
  1.885151e-007, 3.012674e-007, 1.023368e-007, 3.780085e-007, 1.478955e-006, 
    2.09785e-006, 2.5352e-006, 3.290691e-006, 3.682094e-006, 2.977268e-006, 
    2.034272e-006, 1.436487e-006, 1.530613e-006, 2.01341e-006, 1.259163e-006, 
    4.850485e-007, -5.448101e-009, -3.238367e-007, -3.078003e-008, 
    4.496769e-008, -3.798209e-008, -1.065273e-007, -4.661429e-007, 
    -1.100683e-006, -8.374295e-007, -2.23502e-007, -2.904108e-008, 
    1.482827e-007, 2.374404e-007, 1.711305e-007, 6.632536e-008, 
    3.700607e-007, 3.154241e-007, 3.751757e-008, -5.498373e-007, 
    -7.616818e-007, -5.257475e-007, -9.30313e-007, -1.148119e-006, 
    -9.494365e-007, -3.658083e-007, 4.366198e-007, 1.204031e-006, 
    -2.890656e-007, -1.852943e-006, -2.906205e-006, -3.245455e-006, 
    -3.337594e-006, -2.053859e-006, -1.116576e-006, -7.388317e-007, 
    1.651706e-007, 7.329063e-007, 8.81917e-007, 1.611578e-006, 1.692789e-006, 
    7.406043e-007, 9.966561e-007, 1.058495e-006, -4.453796e-009, 
    4.80828e-007, 6.260143e-008, -6.54888e-007, -8.125917e-007, 
    -1.196546e-006, -1.118315e-006, 2.257693e-007, 1.349564e-006, 
    9.869691e-007, -3.773312e-008, 2.230372e-007, 2.06398e-007, 
    -9.022488e-007, -1.879871e-007, 7.366307e-007, 1.191861e-006, 
    1.249382e-007, 4.321491e-007, 1.136974e-006, 1.042353e-006, 7.76864e-007, 
    -4.400636e-007, -1.381571e-006, -5.749207e-007, 5.873717e-007, 
    9.248815e-007, 9.817541e-007, 1.411654e-006, 1.405198e-006, 
    1.863159e-006, 2.760456e-006, 2.386686e-006, 1.861171e-006, 
    1.733519e-006, 8.873794e-007, 1.172375e-007,
  -1.003191e-007, 3.62752e-008, 3.536697e-007, 3.077239e-007, 3.318164e-007, 
    7.824838e-008, 1.506524e-006, 2.733386e-006, 2.224512e-006, 2.68471e-006, 
    2.528247e-006, 2.252327e-006, 3.182906e-006, 5.812464e-006, 
    6.594774e-006, 4.587838e-006, 2.861288e-006, 2.065316e-006, 
    2.419218e-006, 1.512733e-006, 7.530207e-007, -2.506931e-008, 
    -2.282204e-007, -1.201513e-006, -2.269184e-006, -1.658731e-006, 
    -7.125082e-007, 1.063462e-006, 2.058861e-006, 2.058612e-006, 
    2.166149e-006, 2.633301e-006, 1.954553e-006, 3.206396e-007, 
    -1.217159e-006, -3.150089e-006, -5.102886e-006, -5.45679e-006, 
    -6.179744e-006, -5.028382e-006, -2.068763e-006, 9.211544e-007, 
    1.358256e-006, -5.761631e-007, -3.447003e-007, -1.404669e-006, 
    -1.684313e-006, -3.524854e-006, -2.883358e-006, -8.811376e-007, 
    8.300121e-007, 3.842206e-007, -1.932012e-007, -2.696934e-007, 
    1.111645e-006, 1.56588e-006, 1.961258e-006, 2.532469e-006, 3.389037e-006, 
    3.737229e-006, 2.009191e-006, 1.383839e-006, 1.49833e-006, 1.962998e-006, 
    2.240657e-006, 2.084443e-006, 2.188751e-006, 1.266368e-006, 
    1.255688e-006, 1.982367e-006, 2.087172e-006, 8.07162e-007, 
    -8.034031e-007, -1.278255e-006, -1.086277e-006, -4.8129e-007, 
    7.408526e-007, 8.389525e-007, 1.604622e-006, 2.780074e-006, 
    3.042085e-006, 1.855211e-006, 1.418111e-006, 2.524771e-006, 
    2.211351e-006, 1.979637e-006, 3.16552e-006, 3.155834e-006, 3.88773e-006, 
    4.217293e-006, 2.655403e-006, 7.830722e-007, 7.601102e-008, 
    3.328087e-007, 9.442529e-007, 2.876086e-007,
  3.863142e-006, 2.639757e-006, 2.164162e-006, 9.385421e-007, 1.363624e-007, 
    2.992838e-007, 8.08157e-007, -8.237694e-007, -1.926457e-006, 
    -6.387472e-007, 2.150002e-006, 4.685935e-006, 5.421554e-006, 
    6.901488e-006, 8.169576e-006, 6.929056e-006, 5.936389e-006, 
    6.612156e-006, 7.763767e-006, 7.006789e-006, 4.688418e-006, 
    3.971425e-006, 2.724694e-006, 2.251334e-006, 1.303371e-006, 1.94884e-006, 
    2.31814e-006, 2.446042e-006, 4.08815e-006, 4.24784e-006, 5.485628e-006, 
    6.188715e-006, 5.233303e-006, 1.753387e-006, 2.251083e-006, 
    2.569719e-006, 1.955299e-006, -1.652274e-006, -3.614263e-006, 
    -2.734099e-006, -4.544709e-007, 1.867378e-006, 1.00758e-006, 
    -5.299717e-007, 9.027808e-007, 1.418266e-007, -7.664003e-007, 
    -7.112649e-007, -7.647395e-008, -4.216854e-007, 1.251716e-006, 
    1.981127e-006, 2.834465e-006, 3.678617e-006, 5.556909e-006, 
    6.075221e-006, 7.250174e-006, 6.53318e-006, 4.934285e-006, 3.478692e-006, 
    1.492616e-006, 1.340376e-006, 1.228123e-006, 1.892713e-006, 
    2.271449e-006, 3.867116e-006, 4.604971e-006, 3.205009e-006, 
    1.949088e-006, 1.927481e-006, 1.023975e-006, -2.418801e-007, 
    9.119667e-007, 3.064797e-007, -7.534891e-007, 1.099967e-006, 
    2.201659e-006, 1.483175e-006, 2.359611e-006, 2.892828e-006, 
    1.968956e-006, 2.903756e-006, 2.330557e-006, 1.204527e-006, 
    2.391653e-006, 2.970066e-006, 2.661612e-006, 2.840427e-006, 
    3.717111e-006, 2.744562e-006, 2.549606e-006, 2.767162e-006, 
    3.868606e-006, 4.704562e-006, 4.046178e-006, 4.370031e-006,
  7.033858e-006, 4.230705e-006, 1.510249e-006, 2.511359e-006, 4.203634e-006, 
    4.703317e-006, 3.500547e-006, 2.688188e-006, 2.516326e-006, 
    3.979867e-006, 5.494072e-006, 5.754347e-006, 5.220638e-006, 
    8.071476e-006, 9.01919e-006, 5.700454e-006, 4.162655e-006, 4.52972e-006, 
    6.096827e-006, 6.913162e-006, 6.633267e-006, 5.796815e-006, 4.44081e-006, 
    4.904731e-006, 5.977864e-006, 3.471983e-006, 4.233931e-006, 
    4.526244e-006, 4.473593e-006, 3.3945e-006, 3.526871e-006, 2.836452e-006, 
    2.220786e-006, 2.775605e-006, 2.181298e-006, 2.153731e-006, 
    2.766665e-006, 1.780953e-006, 3.114359e-006, 4.710273e-006, 
    2.027566e-006, 2.306218e-006, 2.550847e-006, 2.46566e-006, 3.183646e-006, 
    2.446039e-006, 1.056256e-006, 1.226999e-007, 1.861916e-006, 
    1.574321e-006, 2.071029e-006, 4.584605e-006, 4.849848e-006, 
    3.975396e-006, 4.822776e-006, 8.614874e-006, 6.85902e-006, 6.016606e-006, 
    5.323949e-006, 6.04765e-006, 7.447863e-006, 3.543262e-006, 7.890321e-007, 
    1.844777e-006, 4.399832e-006, 5.1963e-006, 4.806632e-006, 4.574918e-006, 
    5.017981e-006, 3.478443e-006, 2.032531e-006, 3.798817e-006, 
    3.788637e-006, 3.319994e-006, 2.701845e-006, 4.005447e-006, 3.32074e-006, 
    2.813103e-006, 1.863655e-006, -9.137875e-008, 1.331928e-006, 
    3.30832e-006, 4.252308e-006, 3.823156e-006, 5.414598e-006, 4.679723e-006, 
    3.954536e-006, 6.190703e-006, 7.749116e-006, 7.430726e-006, 
    5.364435e-006, 3.966458e-006, 5.414848e-006, 7.84324e-006, 8.170322e-006, 
    7.722044e-006,
  6.841388e-006, 3.930691e-006, 2.07674e-006, 3.790125e-006, 7.797793e-006, 
    8.65014e-006, 7.264827e-006, 5.064176e-006, 4.562751e-006, 7.116065e-006, 
    7.685288e-006, 8.313373e-006, 7.770968e-006, 7.617988e-006, 
    6.660335e-006, 5.186115e-006, 4.379466e-006, 5.237525e-006, 
    5.955511e-006, 6.992881e-006, 6.359831e-006, 6.291533e-006, 
    6.701564e-006, 7.970399e-006, 8.026525e-006, 5.548216e-006, 
    3.479438e-006, 5.77645e-006, 7.625436e-006, 8.039939e-006, 7.789595e-006, 
    5.736962e-006, 6.719198e-006, 4.011408e-006, 2.739594e-006, 
    5.784277e-007, -2.13071e-007, 1.322245e-006, 3.137953e-006, 4.86574e-006, 
    5.899881e-006, 4.528973e-006, 4.902746e-006, 7.45879e-006, 6.691382e-006, 
    2.086923e-006, 1.771765e-006, 2.955414e-006, 4.442798e-006, 
    3.450876e-006, 2.604242e-006, 4.078709e-006, 5.358472e-006, 4.60845e-006, 
    5.795571e-006, 6.522998e-006, 6.745524e-006, 8.046145e-006, 
    7.491326e-006, 6.462398e-006, 6.674991e-006, 6.16959e-006, 5.12378e-006, 
    6.136561e-006, 5.480912e-006, 5.338108e-006, 5.542006e-006, 
    3.507748e-006, 5.858903e-006, 5.732989e-006, 7.517401e-006, 
    9.085748e-006, 7.625187e-006, 5.618247e-006, 4.589572e-006, 
    5.393988e-006, 5.02096e-006, 5.275027e-006, 4.754973e-006, 3.188616e-006, 
    8.829102e-007, 1.926239e-006, 3.64484e-006, 5.888705e-006, 6.609675e-006, 
    5.859152e-006, 5.379334e-006, 7.188584e-006, 8.257992e-006, 
    8.658335e-006, 7.874534e-006, 8.655106e-006, 1.018272e-005, 
    1.161547e-005, 9.475911e-006, 7.772462e-006,
  8.368754e-006, 7.479402e-006, 8.400544e-006, 6.662571e-006, 4.530961e-006, 
    4.95614e-006, 6.699578e-006, 6.048151e-006, 7.832814e-006, 7.8425e-006, 
    7.066645e-006, 6.97724e-006, 3.8994e-006, 5.250331e-007, -3.330279e-007, 
    1.129774e-006, 3.906358e-006, 4.918142e-006, 5.245967e-006, 8.04441e-006, 
    9.547439e-006, 7.219627e-006, 7.20249e-006, 7.403407e-006, 6.761913e-006, 
    6.616383e-006, 5.73895e-006, 5.949056e-006, 7.479408e-006, 9.474919e-006, 
    1.017204e-005, 7.804001e-006, 5.100434e-006, 3.838553e-006, 
    5.236281e-006, 6.439055e-006, 7.113087e-006, 6.707272e-006, 
    6.493698e-006, 6.555036e-006, 6.154445e-006, 5.090002e-006, 
    7.168464e-006, 5.721568e-006, 5.900878e-006, 4.236417e-006, 
    3.289446e-006, 6.322078e-006, 4.467631e-006, 2.445548e-006, 
    3.689296e-006, 3.743931e-006, 3.960746e-006, 5.742924e-006, 7.59762e-006, 
    7.433957e-006, 7.197279e-006, 5.63862e-006, 5.847731e-006, 5.502769e-006, 
    7.220373e-006, 5.407153e-006, 4.322843e-006, 6.809099e-006, 
    7.109362e-006, 4.807131e-006, 7.655239e-006, 1.015491e-005, 
    9.143119e-006, 4.761929e-006, 4.252563e-006, 6.160904e-006, 
    6.449738e-006, 6.716466e-006, 6.103774e-006, 3.566609e-006, 
    3.677873e-006, 5.398961e-006, 4.563746e-006, 1.458591e-006, 
    1.010563e-006, 1.117352e-006, 4.505629e-006, 4.239646e-006, 
    4.401321e-006, 6.189957e-006, 7.215409e-006, 6.998343e-006, 
    7.410858e-006, 6.671269e-006, 3.266852e-006, 4.361837e-006, 6.88758e-006, 
    7.480399e-006, 9.043031e-006, 9.471936e-006,
  3.371901e-006, 2.972552e-006, 2.478824e-006, 1.987835e-006, 5.903457e-007, 
    2.183289e-006, 4.175075e-006, 4.90672e-006, 4.217043e-006, 2.576679e-006, 
    4.763919e-006, 4.884372e-006, 1.197328e-006, -2.59759e-007, 
    1.224893e-006, 5.490601e-006, 7.272276e-006, 8.912401e-006, 
    1.015118e-005, 1.093176e-005, 8.241597e-006, 9.464493e-006, 
    9.410101e-006, 6.649418e-006, 7.400678e-006, 6.168601e-006, 
    3.864883e-006, 2.760207e-006, 3.291934e-006, 3.23506e-006, 1.898425e-006, 
    1.266617e-006, 1.450644e-006, 2.20216e-006, 3.606594e-006, 2.46815e-006, 
    1.920525e-006, 9.499636e-007, 1.057007e-006, 4.361282e-007, 3.23233e-006, 
    4.740581e-006, 2.68521e-006, 1.114622e-006, 3.210971e-006, 4.123667e-006, 
    2.66459e-006, 1.774992e-006, -3.660498e-007, 5.240363e-007, 
    1.283999e-006, 2.706813e-006, 5.710888e-006, 5.558148e-006, 
    1.039879e-005, 1.220258e-005, 7.989518e-006, 6.844864e-006, 
    8.153926e-006, 8.175535e-006, 7.740418e-006, 6.068516e-006, 
    3.542766e-006, 1.888988e-006, -1.203003e-006, 2.515331e-006, 
    4.287827e-006, 4.978243e-006, 2.814846e-006, 3.679856e-006, 
    4.412501e-006, 3.41214e-006, 2.174347e-006, 2.626595e-006, 1.272572e-006, 
    -2.002449e-006, -1.140419e-006, -4.781021e-006, -1.961222e-006, 
    -2.915531e-007, 5.896036e-007, 1.015776e-006, 2.488265e-006, 
    2.469638e-006, 3.101446e-006, 2.845143e-006, 1.091525e-006, 2.40705e-006, 
    6.879134e-006, 9.54992e-006, 8.830197e-006, 7.266815e-006, 8.157407e-006, 
    6.04691e-006, 1.807028e-006, 1.906621e-006,
  1.244764e-006, 1.872591e-006, 7.656854e-007, -1.575783e-006, 
    -2.337481e-006, 7.13786e-007, -7.424023e-008, 1.023478e-006, 
    1.479701e-006, 2.141067e-006, 3.567606e-006, -1.022705e-006, 
    -1.863373e-006, 7.4524e-008, 3.830115e-006, 6.706287e-006, 8.570667e-006, 
    7.675357e-006, 5.239763e-006, 1.205524e-006, -6.926348e-007, 
    1.451142e-006, 3.293353e-007, 5.672555e-007, 8.041861e-007, 
    -1.154822e-006, -3.443394e-006, -2.012388e-006, -3.419555e-006, 
    -5.726746e-006, -6.031478e-006, -2.481029e-006, -3.915757e-006, 
    -4.240606e-006, -4.17827e-006, -3.552424e-006, -3.52833e-006, 
    -4.241352e-006, -2.642708e-006, -5.001639e-007, 7.582366e-007, 
    -1.405413e-006, -3.643068e-006, -2.578381e-006, 4.977155e-007, 
    3.79503e-007, -1.338849e-006, 2.027817e-006, 1.372911e-006, 
    3.273308e-006, 6.096579e-006, 7.433213e-006, 8.690618e-006, 
    8.376704e-006, 9.261086e-006, 8.448482e-006, 7.399685e-006, 
    7.063412e-006, 5.092737e-006, -5.083602e-007, -3.845969e-006, 
    -2.256762e-006, -4.452944e-006, -5.288402e-006, -1.646556e-006, 
    1.348817e-006, -6.740083e-007, -4.504946e-007, -1.089509e-006, 
    -1.281234e-006, -2.962828e-006, -4.100286e-006, -5.427728e-006, 
    -6.145967e-006, -8.459623e-006, -1.141328e-005, -1.139565e-005, 
    -1.461752e-005, -6.321055e-006, -2.493307e-007, 1.154356e-006, 
    5.011916e-007, 1.099972e-006, 2.472116e-006, 2.737113e-006, 
    6.887021e-007, 4.520225e-007, 3.259152e-006, 4.219033e-006, 3.02694e-006, 
    3.403442e-006, 5.328675e-006, 4.444541e-006, 2.852848e-006, 
    3.176199e-006, 1.713153e-006,
  -7.805575e-007, -2.47432e-006, -5.71135e-006, -7.450319e-006, 
    -6.856753e-006, -6.012602e-006, -2.971276e-006, -2.510333e-006, 
    -1.17544e-006, -1.076343e-006, -3.328156e-006, -1.572056e-006, 
    8.496318e-007, 3.423806e-006, 1.759847e-006, -3.302921e-007, 
    -2.447498e-006, -2.678968e-006, -4.369505e-006, -8.481973e-006, 
    -1.307277e-005, -1.174259e-005, -9.933345e-006, -9.831519e-006, 
    -1.05736e-005, -8.730078e-006, -8.085852e-006, -6.867927e-006, 
    -8.256224e-006, -8.150921e-006, -7.240213e-006, -7.336821e-006, 
    -6.391343e-006, -5.205458e-006, -2.371506e-006, -2.531691e-006, 
    -5.281207e-006, -5.119777e-006, -4.015104e-006, -4.133813e-006, 
    -2.474319e-006, -2.268687e-006, -3.661198e-006, -3.530571e-006, 
    -8.808303e-006, -9.25261e-006, -3.339577e-006, 2.294051e-006, 
    2.255547e-009, 1.988581e-006, 2.053897e-006, 3.028683e-006, 
    4.396108e-006, 7.204977e-006, 5.691763e-006, 6.167113e-006, 
    3.897916e-006, -1.974386e-006, -6.347876e-006, -4.281825e-006, 
    -2.680947e-006, -2.502144e-006, -2.619356e-006, -3.53553e-006, 
    -1.661712e-006, -3.050503e-006, -8.020288e-006, -5.957467e-006, 
    -6.646645e-006, -9.591859e-006, -9.46123e-006, -9.124215e-006, 
    -8.146202e-006, -8.27013e-006, -8.837615e-006, -1.079985e-005, 
    -1.348975e-005, -1.465701e-005, -6.992602e-006, -1.167738e-006, 
    1.938655e-006, 3.261879e-006, 6.948427e-006, 8.610157e-006, 
    6.325066e-006, 6.716964e-006, 1.547254e-006, -4.127432e-007, 
    -1.826367e-006, -1.335622e-006, -1.591761e-007, -3.388504e-006, 
    -3.457302e-006, -2.747511e-006, -2.004435e-006, -6.409791e-007,
  -6.299204e-006, -7.397914e-006, -4.610152e-006, -3.58123e-006, 
    -4.179758e-006, -3.022189e-006, -2.781037e-006, -2.216034e-006, 
    -2.258999e-006, -4.331141e-007, 2.074505e-006, 7.820781e-007, 
    -3.95612e-007, -9.419873e-007, -3.775194e-006, -2.977236e-006, 
    -2.957864e-006, -4.372976e-006, -8.335195e-006, -8.515253e-006, 
    -7.444109e-006, -7.399651e-006, -7.810428e-006, -8.473775e-006, 
    -6.830925e-006, -6.030483e-006, -6.044393e-006, -5.611515e-006, 
    -5.060916e-006, -4.04242e-006, -2.36008e-006, -3.237757e-006, 
    -3.058198e-006, -3.948297e-006, -3.895397e-006, -2.800906e-006, 
    -2.885346e-006, -6.487949e-006, -7.839732e-006, -4.858757e-006, 
    -1.397715e-006, -2.080682e-006, -2.679462e-006, -3.055964e-006, 
    -3.227069e-008, 1.400227e-006, 5.804519e-006, 3.399466e-006, 
    5.307065e-006, 1.949338e-006, 6.435828e-006, 6.873921e-006, 
    6.830458e-006, 3.592191e-006, 3.013531e-006, -1.552686e-006, 
    -4.663549e-006, -9.73516e-006, -5.777911e-006, -4.34914e-006, 
    -4.914633e-006, -6.949385e-006, -8.181465e-006, -9.063364e-006, 
    -8.525187e-006, -8.356556e-006, -6.232645e-006, -6.68862e-006, 
    -7.395682e-006, -7.289136e-006, -6.656335e-006, -6.078168e-006, 
    -6.421639e-006, -6.148452e-006, -5.776171e-006, -5.058185e-006, 
    -7.068847e-006, -5.347514e-006, -4.096091e-008, 2.989686e-006, 
    4.592799e-006, 7.547453e-006, 4.309926e-006, 3.262623e-006, 
    3.142919e-006, -1.551944e-006, -2.152454e-006, 9.022879e-007, 
    -1.113596e-006, -1.276265e-006, -4.012123e-006, -6.244565e-006, 
    -5.46374e-006, -2.602719e-006, -3.051246e-006, -6.101267e-006,
  -3.228818e-006, -2.126876e-006, -1.01972e-006, -9.732785e-007, 
    -9.802329e-007, -1.283223e-006, -4.482617e-007, -5.120855e-007, 
    8.583229e-007, -8.426487e-007, -3.645308e-006, -2.850576e-006, 
    -4.336071e-007, -4.427984e-007, 4.651793e-007, 3.522153e-006, 
    4.325077e-006, -1.180153e-006, -6.376436e-006, -1.92894e-006, 
    -4.253274e-006, -5.666647e-006, -4.71943e-006, -7.311337e-007, 
    -1.281333e-007, -3.66393e-006, -4.18249e-006, -1.451854e-006, 
    -6.496739e-007, 1.539059e-006, 3.116097e-006, 1.700736e-006, 
    -7.308863e-007, -1.26832e-006, 4.53756e-007, -3.275609e-007, 
    -3.237261e-006, -1.888458e-006, -2.023908e-007, 2.715755e-006, 
    6.337978e-006, 9.247922e-006, 5.765027e-006, 1.730785e-006, 
    1.825656e-006, 6.720935e-006, 1.368971e-005, 1.24261e-005, 6.730123e-006, 
    9.301075e-006, 1.548729e-005, 9.813422e-006, 1.444683e-006, 
    -1.095217e-006, -3.492072e-006, -8.216235e-006, -9.916208e-006, 
    -9.948e-006, -4.276366e-006, -3.449848e-006, -4.754693e-006, 
    -6.148201e-006, -6.289018e-006, -5.877002e-006, -5.341803e-006, 
    -6.683653e-006, -3.680077e-006, -5.542226e-006, -7.057423e-006, 
    -5.572273e-006, -5.217624e-006, -2.945445e-006, -2.377962e-006, 
    -3.386026e-006, -3.441904e-006, -2.275888e-006, -2.155685e-006, 
    -1.125022e-006, -6.707833e-007, 1.786415e-006, 4.0749e-008, 
    -4.524845e-007, -9.571359e-007, 8.789357e-007, -6.841965e-007, 
    1.382346e-006, -5.314541e-007, -2.859018e-006, -2.17804e-006, 
    -9.288269e-007, -2.259747e-006, -2.193687e-006, -2.406276e-006, 
    -3.863855e-006, -4.365279e-006, -3.533296e-006,
  -1.216772e-007, 4.833091e-007, 4.273215e-008, -1.092488e-006, 
    -7.346114e-007, -1.370643e-006, 1.323239e-006, 8.270308e-007, 
    -5.911523e-006, -6.078666e-006, -2.190205e-006, 1.983362e-006, 
    7.287179e-006, 2.996887e-006, -2.146002e-006, 1.107424e-006, 
    9.598105e-006, 6.21554e-006, -2.207838e-006, -1.983082e-006, 
    -2.272911e-006, -2.500783e-007, 6.517286e-006, 3.531592e-006, 
    -1.259627e-006, -1.342081e-006, 1.558428e-006, 1.974669e-006, 
    5.034271e-007, 2.254315e-006, 1.886255e-006, 5.367065e-007, 
    2.185652e-007, -1.260374e-006, -1.621725e-006, -4.141762e-006, 
    -3.711367e-006, 7.54264e-007, 3.790128e-006, 2.300505e-006, 6.71423e-006, 
    1.419884e-005, 3.396734e-006, -5.989261e-006, 2.761844e-007, 
    9.670122e-006, 2.041038e-005, 1.082869e-005, 7.858398e-006, 
    1.327323e-005, 8.073963e-006, 4.62782e-006, 6.663468e-007, 
    -4.103513e-006, -7.084489e-006, -3.61972e-006, -3.991754e-006, 
    -3.592402e-006, 7.795988e-007, -4.681182e-006, -7.788074e-006, 
    -5.768719e-006, -4.660073e-006, -3.986044e-006, -5.780146e-006, 
    -7.807201e-006, -8.3876e-006, -8.495136e-006, -5.39793e-006, 
    -4.097554e-006, -1.312032e-006, -3.131572e-007, -1.537137e-007, 
    7.00511e-008, -4.668875e-007, 3.318148e-007, -1.686153e-007, 
    -3.551287e-007, 5.024349e-007, 8.967534e-006, 7.009279e-006, 
    1.010797e-005, 6.448994e-006, 4.295525e-006, 2.639757e-006, 
    1.168766e-006, 9.242707e-006, 1.273504e-005, 1.183129e-005, 
    5.853439e-006, 2.920147e-006, -1.313523e-006, -2.151462e-006, 
    -2.311402e-006, -1.130486e-006, -1.392747e-006,
  9.513496e-008, 2.568122e-007, -9.95879e-007, -4.994213e-007, 3.405073e-007, 
    2.76766e-006, 3.911072e-006, -5.93561e-006, -7.92442e-006, 
    -1.163766e-006, 2.51707e-006, 6.01785e-006, 8.503615e-006, 4.152971e-006, 
    -5.520364e-006, -4.809579e-006, -2.461409e-006, 8.693103e-006, 
    2.364583e-006, -1.001257e-005, -9.730693e-006, -4.656598e-006, 
    -2.158169e-006, 8.508741e-007, -8.011684e-007, 2.322611e-006, 
    2.073921e-007, -1.90783e-006, -1.772477e-006, 4.105535e-006, 1.6538e-006, 
    3.16254e-006, -2.947772e-007, -2.314381e-006, 1.247245e-006, 
    1.018016e-006, 4.679141e-007, 4.115718e-006, 1.219215e-005, 
    7.773951e-006, 3.203764e-006, 8.242592e-006, -3.257132e-006, 
    -1.738203e-006, 5.656995e-006, 3.70196e-006, 2.092025e-005, 
    1.391323e-005, 2.979257e-006, 5.933656e-006, 3.80478e-006, 2.587101e-006, 
    4.941492e-006, -1.849963e-006, -1.703438e-006, 3.564019e-007, 
    -4.770718e-007, -3.938854e-006, -9.532505e-006, -1.104696e-005, 
    -1.370607e-005, -8.887782e-006, -5.096927e-006, -7.853145e-006, 
    -1.188292e-005, -1.015513e-005, -8.214744e-006, -5.387747e-006, 
    -1.655504e-006, -7.197095e-007, 7.356357e-007, 4.974672e-007, 
    -6.803339e-008, 2.587994e-007, -2.798779e-007, 1.071657e-006, 
    -2.354225e-007, -3.017327e-007, -8.483557e-007, 1.189958e-005, 
    9.790328e-006, 6.023562e-006, -2.392368e-006, -9.856958e-007, 
    -3.49628e-006, 1.38335e-005, 1.932359e-005, 1.524192e-005, 1.246004e-006, 
    2.009328e-007, -1.066412e-006, -3.220966e-007, -8.811403e-007, 
    -3.772311e-007, 9.052619e-007, 3.8695e-007,
  -7.442968e-007, -4.817894e-007, -2.679571e-007, -3.275612e-007, 
    1.860672e-006, 4.273177e-006, -1.597637e-006, -4.809335e-006, 
    -6.784234e-006, -1.285458e-006, -1.3838e-006, 6.960843e-006, 
    1.700895e-005, 3.827376e-006, -7.734179e-006, -1.442332e-005, 
    8.644201e-008, 1.03742e-005, 2.431516e-007, -1.072658e-005, 
    -1.215164e-005, -3.57204e-006, 7.808376e-007, -5.086094e-007, 
    -1.482401e-006, -1.068894e-006, -4.718549e-007, 1.803219e-007, 
    -9.784926e-007, 1.031671e-006, -3.680452e-007, 3.920011e-006, 
    -3.476676e-006, 2.94697e-006, 7.583216e-006, 4.221018e-006, 3.13646e-006, 
    7.86584e-006, 9.614989e-006, 2.182045e-006, 4.838423e-006, 1.018223e-005, 
    1.048994e-005, 2.230606e-005, 3.887231e-006, 8.666288e-006, 
    1.544905e-005, 5.540933e-007, -3.611029e-006, 3.851219e-006, 
    1.839625e-005, 1.837911e-005, 1.780517e-005, 3.796584e-006, 
    5.888069e-008, 6.329035e-006, 2.255303e-006, -2.718203e-006, 
    -7.915478e-006, -8.936702e-006, -6.682902e-006, -1.035331e-005, 
    -1.04827e-005, -1.127272e-005, -9.287878e-006, -4.967285e-006, 
    -2.321583e-006, -3.176256e-007, 4.607118e-007, 4.597186e-007, 
    7.34397e-007, -3.213518e-007, -3.784735e-007, 6.3282e-007, 7.377616e-008, 
    1.087942e-007, -7.013321e-007, -6.938137e-009, -6.863709e-006, 
    3.307323e-006, 1.043009e-005, 2.707166e-007, -7.110324e-006, 
    -5.48461e-006, -3.104156e-006, -4.300709e-006, 3.462046e-006, 
    -7.531024e-006, -9.109806e-006, -2.651648e-006, -1.100185e-006, 
    -3.004889e-007, -1.134786e-007, -6.529899e-008, 4.845542e-007, 
    -9.521682e-007,
  -3.722644e-007, -3.871664e-007, 3.449777e-007, 1.703854e-007, 
    -1.590932e-006, -2.026045e-006, -1.077054e-005, -1.243922e-005, 
    -7.423496e-006, -4.471076e-006, 1.330191e-006, 1.747983e-005, 
    2.102928e-005, 1.373765e-005, 8.836505e-007, -7.460258e-006, 
    5.513699e-006, 1.138948e-005, 1.04732e-006, -6.004902e-006, 
    -1.188341e-005, -1.613284e-006, -2.156181e-006, 9.437554e-007, 
    1.292194e-006, -4.922185e-007, 1.562401e-006, -2.321834e-006, 
    -2.589559e-006, -3.313005e-006, -4.348476e-007, 8.1486e-007, 
    -1.122353e-007, -1.050519e-006, 7.212178e-006, 1.142151e-005, 
    8.898989e-006, 7.611779e-006, 1.257734e-005, 1.709537e-005, 
    5.851205e-006, -1.516426e-006, 5.618251e-006, 2.435646e-005, 
    1.519224e-005, 1.68649e-005, 3.197394e-005, 2.182377e-005, 2.355875e-005, 
    8.681935e-006, 2.414537e-005, 3.130687e-005, 4.060767e-005, 
    3.842042e-005, 1.622763e-005, 1.535343e-005, 1.02555e-005, 9.869764e-007, 
    -7.32117e-006, -9.585154e-006, -1.226091e-005, -1.90695e-005, 
    -1.659615e-005, -1.067244e-005, -4.530434e-006, -1.216416e-006, 
    2.006855e-007, 7.9847e-007, 1.207163e-007, -7.796643e-008, 
    -1.139779e-007, -3.263185e-007, -9.218675e-007, -4.37085e-007, 
    -2.163881e-006, -5.833635e-007, -3.372472e-007, -4.010739e-007, 
    -1.244121e-005, 1.568472e-005, 1.546245e-005, 3.428024e-006, 
    -3.485617e-006, -4.66207e-006, -2.220258e-007, 3.328169e-007, 
    -3.009271e-006, -1.504493e-005, -1.060166e-005, -1.87803e-006, 
    1.050548e-006, 8.295146e-007, 1.151629e-006, 1.704958e-006, 
    -4.735903e-007, -4.631602e-007,
  -2.2816e-006, -6.551395e-007, -8.392772e-008, 6.119581e-007, 3.586731e-006, 
    -1.574295e-006, -8.308376e-006, -1.484502e-005, -5.300575e-006, 
    -3.809961e-006, 6.500897e-006, 1.311999e-005, 9.390475e-006, 
    4.766407e-006, -3.937617e-006, -1.072832e-005, 2.20356e-005, 
    2.913228e-005, 1.424528e-005, -1.475736e-005, -1.97999e-005, 
    -1.101889e-005, -9.702373e-006, -1.621556e-007, -3.957477e-006, 
    1.357021e-006, 6.115701e-006, -2.30455e-007, 1.450397e-006, 
    6.208837e-006, 4.132853e-006, -1.555665e-006, -5.656962e-006, 
    7.589879e-007, 1.392018e-005, 1.535293e-005, 1.762337e-005, 
    2.973553e-006, 3.777818e-005, 3.611275e-005, 2.436963e-005, 
    5.038586e-006, 1.499977e-005, 2.387267e-005, 3.911531e-005, 
    2.753959e-005, 3.098723e-005, 4.202924e-005, 1.842927e-005, 
    -2.278612e-006, 5.509472e-006, 2.346786e-005, 3.337836e-005, 
    4.612085e-005, 2.178005e-005, 2.089641e-005, 1.742395e-005, 
    6.179274e-006, 2.209366e-006, -6.242328e-006, -1.80125e-005, 
    -1.971074e-005, -1.439947e-005, -6.761138e-006, -2.122158e-006, 
    1.147555e-007, 1.283503e-006, 5.856327e-007, 3.583909e-007, 
    -3.275582e-007, -1.113596e-006, -1.599125e-006, -9.665719e-007, 
    -2.114459e-006, -1.733238e-006, 4.549978e-007, 2.456367e-007, 
    -9.900066e-006, -8.85893e-006, 1.45649e-005, 1.068514e-005, 
    3.576548e-006, -1.887725e-006, -1.497465e-007, -1.860135e-006, 
    8.086627e-006, -1.067691e-005, -1.657852e-005, -5.142127e-006, 
    -3.489837e-006, -1.368157e-006, -1.721673e-009, -6.017417e-007, 
    -4.470176e-007, -7.033168e-007, -9.109399e-007,
  -1.079573e-006, -1.075104e-006, 7.22971e-007, -1.338602e-006, 
    1.639419e-007, 8.854287e-006, 3.174704e-006, 8.955365e-006, 
    -5.913171e-007, 3.906753e-007, 9.5832e-006, 2.285914e-005, 8.197145e-006, 
    -4.741785e-006, -2.355606e-006, -4.488713e-006, 2.010516e-005, 
    2.753364e-005, 1.115503e-005, 4.892063e-006, -7.930386e-006, 
    -2.414708e-006, -4.873647e-006, -7.225026e-008, 2.94052e-006, 
    1.633915e-005, 7.314993e-006, 3.139688e-006, 3.915542e-006, 4.88064e-006, 
    6.199647e-006, 2.477827e-006, -6.913629e-006, -1.027176e-006, 
    9.290961e-007, 1.725779e-005, 1.576047e-005, 1.343292e-005, 
    3.192775e-005, 3.642441e-005, 2.749613e-005, 2.717651e-005, 2.86865e-005, 
    4.549303e-005, 4.313019e-005, 3.287099e-005, 3.43569e-005, 6.12669e-005, 
    3.014805e-005, 1.541825e-005, -5.03211e-006, 2.807108e-005, 
    4.097224e-005, 1.558862e-005, 1.367904e-005, 1.917357e-005, 
    1.069731e-005, 1.026021e-005, 9.062656e-006, -1.616259e-006, 
    -8.990843e-006, -1.331491e-005, -1.209426e-005, -6.452932e-006, 
    -7.574599e-007, 1.84792e-007, -2.232509e-007, -6.149048e-007, 
    -1.477681e-006, -2.301467e-006, -2.365046e-006, -2.262477e-006, 
    -2.817794e-006, -1.533065e-006, 8.518655e-007, 1.611079e-006, 
    9.842406e-007, -1.071616e-005, 1.482667e-005, 6.307928e-006, 
    4.424423e-006, 7.715586e-006, -7.845942e-006, -1.616575e-005, 
    -2.243847e-006, 2.302828e-005, -2.661589e-006, -3.973619e-006, 
    -3.302328e-006, -6.141599e-007, 1.570845e-006, 4.227131e-007, 
    -8.674797e-007, -1.623216e-006, -1.305077e-006, -1.486127e-006,
  3.722079e-006, 3.21842e-006, 7.28122e-006, 8.163515e-007, 3.652531e-008, 
    1.403592e-005, 1.798621e-005, 9.510681e-006, 4.129368e-006, 
    2.256662e-005, 2.3938e-005, 2.578225e-005, 1.352183e-005, 4.78304e-006, 
    9.800744e-006, 2.08229e-005, 2.105858e-005, 2.070717e-005, 9.826086e-006, 
    -3.720816e-006, -9.716285e-006, 4.060334e-006, -3.356967e-006, 
    6.806658e-008, 1.016335e-005, 1.924927e-007, 2.923123e-006, 
    5.402188e-006, 1.646306e-005, 9.905067e-006, 3.787893e-006, 
    1.527515e-007, 2.904751e-006, 9.391726e-006, 6.500151e-006, 
    -5.570284e-006, -6.29299e-006, 1.672359e-005, 1.972146e-005, 
    7.823124e-006, 5.862661e-006, 4.047755e-005, 5.290411e-005, 
    4.389288e-005, 4.527894e-005, 2.055918e-005, 2.180516e-005, 
    3.533445e-005, 4.192593e-005, -8.543138e-007, -1.622881e-005, 
    1.679266e-005, 2.9253e-005, 1.197959e-005, 1.207717e-005, 2.336629e-005, 
    2.131663e-005, 2.095255e-005, 1.702459e-005, 1.283215e-005, 
    7.597373e-006, -9.943833e-007, -1.173713e-005, -8.583298e-006, 
    -1.808987e-006, -8.210409e-007, -1.164013e-006, -2.179031e-006, 
    -2.2441e-006, -9.792388e-007, -8.359398e-007, -1.934513e-007, 
    -1.406654e-006, 1.028692e-006, 5.663453e-006, 1.326528e-005, 
    -2.627276e-006, 5.025431e-006, 7.146115e-006, 9.698851e-009, 
    1.127039e-006, -8.481147e-007, -7.411574e-006, -1.435875e-005, 
    -8.322531e-006, 2.003711e-005, 7.469476e-006, 4.321351e-006, 
    -3.81071e-006, -5.400165e-006, -5.617549e-007, 5.918515e-006, 
    9.366389e-006, 1.098813e-005, 4.689661e-006, 4.717227e-006,
  1.300103e-005, 1.330303e-005, 8.782015e-006, 3.009802e-006, -3.193303e-006, 
    -2.348155e-006, -3.388268e-006, -3.121677e-007, 1.206921e-005, 
    2.756046e-005, 2.320882e-005, 1.74689e-005, 1.866918e-005, 1.71063e-005, 
    1.590725e-005, 8.277362e-006, 1.323796e-005, 9.011746e-006, 
    3.591456e-006, 2.261513e-006, 1.325971e-006, 4.55902e-006, 4.769383e-006, 
    3.555433e-006, 6.190952e-006, 8.442519e-006, 1.29901e-005, 8.755182e-006, 
    1.102638e-005, 2.257999e-005, 1.573293e-005, 1.166962e-005, 
    1.407019e-005, 1.378619e-006, -1.574753e-005, -7.071838e-006, 
    8.147486e-006, 5.938188e-005, 2.327614e-005, 1.851126e-005, 
    9.124269e-006, 9.613301e-006, 3.692068e-006, 1.479985e-005, 2.65961e-005, 
    -2.353321e-006, -2.200202e-005, -3.016515e-005, -2.295891e-005, 
    -2.637679e-005, -1.449631e-005, -6.892733e-006, -8.660296e-006, 
    -8.113901e-006, 8.434319e-006, 1.687558e-005, 1.725258e-005, 
    1.666324e-005, 2.106404e-005, 2.560891e-005, 2.570055e-005, 
    2.249258e-005, 2.019506e-005, 1.546643e-005, 1.275591e-005, 
    1.465878e-005, 1.322405e-005, 1.055004e-005, 7.908558e-006, 
    1.031981e-005, 4.988429e-006, 6.590799e-006, 8.386638e-006, 
    9.747114e-006, 6.459171e-006, 6.488233e-006, 5.280986e-006, 
    2.671793e-006, -8.777519e-006, -1.747394e-006, 4.78006e-006, 
    4.780799e-006, -8.024144e-007, -8.408464e-006, -4.418675e-006, 
    3.186542e-007, -6.757658e-006, -6.195143e-006, 7.338967e-007, 
    -9.315481e-007, -5.608777e-006, 1.181928e-006, 2.944489e-006, 
    8.280596e-006, 1.242486e-005, 9.680556e-006,
  -1.949054e-006, -4.171812e-006, -2.107012e-006, 2.060104e-006, 
    -4.385392e-006, -6.767339e-006, -5.624934e-006, -1.169764e-005, 
    1.033332e-007, 1.679462e-005, 1.022619e-005, 2.118465e-006, 
    7.941839e-006, 7.715336e-006, 1.139096e-005, 7.860624e-006, 
    1.016137e-005, 4.714238e-006, -1.434484e-006, -5.073569e-006, 
    -2.104774e-006, 1.226384e-006, 1.066677e-005, 7.863608e-006, 
    7.953764e-006, 9.088973e-006, 1.743164e-005, 1.394019e-006, 
    9.350733e-006, 2.461749e-005, 2.054598e-005, 2.369584e-005, 
    7.176903e-006, -7.316936e-006, -2.930436e-005, -1.290564e-005, 
    1.710505e-005, 2.835617e-005, 2.614361e-005, 2.419554e-005, 
    5.197799e-006, -1.765834e-005, -2.433681e-005, -2.334116e-005, 
    -3.182761e-005, -4.801054e-005, -4.971596e-005, -3.701025e-005, 
    -2.621262e-005, -2.939129e-005, -2.690453e-005, -2.447415e-005, 
    -1.598446e-005, -1.15531e-005, -5.400663e-006, -9.839569e-007, 
    1.991939e-007, -1.392253e-006, 5.48127e-007, 1.168019e-006, 4.08964e-006, 
    4.854315e-006, 6.046161e-006, 9.164476e-006, 9.046013e-006, 
    1.056543e-005, 1.208734e-005, 1.290243e-005, 1.13013e-005, 1.353648e-005, 
    1.292429e-005, 1.608185e-005, 1.589484e-005, 1.696101e-005, 
    4.200905e-006, 4.413378e-007, 1.221872e-005, 6.7726e-006, 5.851456e-006, 
    8.51305e-006, 5.641101e-006, -2.291533e-006, -7.403232e-007, 
    -9.325131e-006, -6.636217e-006, -4.052847e-006, -9.578947e-006, 
    -7.120252e-006, -8.558218e-006, -5.32069e-006, -2.846107e-006, 
    9.910946e-008, 7.612216e-007, 6.049995e-007, -1.236782e-006, 2.940687e-007,
  -8.232622e-006, -6.553855e-007, -2.630284e-006, -1.163481e-005, 
    -1.270521e-005, -1.161991e-005, -4.398556e-006, -4.520249e-006, 
    -2.626313e-006, 4.130618e-006, 2.698368e-006, 5.131125e-007, 
    1.281764e-006, 2.500431e-006, 1.178708e-005, 1.230713e-005, 
    1.749249e-005, 9.220606e-006, 1.997021e-006, 3.370413e-006, 
    2.555065e-006, 4.343856e-007, 5.997863e-007, 1.792872e-006, 
    8.052353e-006, 1.011542e-005, 5.643582e-006, -3.366898e-006, 
    9.979325e-006, 6.73061e-006, -3.575406e-008, 1.157821e-005, 
    1.661134e-005, 1.843284e-006, -1.117442e-007, 1.511246e-006, 
    -4.811074e-006, -2.940236e-006, 5.575777e-006, 4.245609e-006, 
    4.866983e-006, 2.838191e-006, -7.090348e-007, 6.534319e-007, 
    -4.545087e-006, -7.416034e-006, -3.360936e-006, -2.108936e-008, 
    -6.07891e-006, -1.00456e-005, -8.187177e-006, -6.754181e-006, 
    -7.171668e-006, -6.582575e-006, -3.492072e-006, -1.961476e-006, 
    -4.278954e-007, -2.885718e-007, -1.65153e-006, -2.148236e-006, 
    -9.733685e-008, 8.600618e-007, 2.145536e-006, 4.601993e-006, 
    6.762661e-006, 6.957369e-006, 5.734233e-006, 4.627822e-006, 
    5.789864e-006, 1.10229e-005, 1.127126e-005, 1.307901e-005, 1.041915e-005, 
    1.585211e-005, 1.390602e-005, 2.220226e-005, 2.012304e-005, 
    9.579229e-006, 1.046759e-005, 6.090867e-006, 4.733758e-007, 
    -1.141165e-006, -3.924205e-006, -1.134101e-005, -1.103653e-005, 
    -1.079712e-005, -7.967884e-006, -5.846205e-006, -4.804863e-006, 
    -2.807361e-006, -2.109495e-006, -2.258257e-006, -2.533052e-007, 
    3.963731e-006, 2.50242e-006, -6.941191e-007,
  -3.542986e-006, -3.916255e-006, -4.040683e-006, -5.434934e-006, 
    -5.286171e-006, -7.235493e-006, -6.883575e-006, -3.547454e-006, 
    -2.855904e-007, -9.357766e-007, 2.939023e-006, 8.399443e-007, 
    1.296559e-007, -8.803945e-007, 2.365328e-006, 9.002801e-006, 
    1.327372e-005, 1.221276e-005, 8.235886e-006, 4.417712e-006, 
    1.076113e-005, 6.136808e-006, -6.42227e-007, -1.905595e-006, 
    5.049522e-006, 6.293281e-006, 2.958041e-007, 8.384523e-007, 
    5.111859e-006, 9.065079e-007, 2.15671e-006, 5.521142e-006, 2.060162e-005, 
    9.060168e-006, 4.473099e-006, 1.581413e-005, 1.487882e-005, 
    1.491435e-005, 1.327968e-005, 1.347911e-005, 1.503008e-005, 
    1.198279e-005, 1.00198e-005, 9.277977e-006, 8.511064e-006, 1.004116e-005, 
    9.169198e-006, 8.283574e-006, 6.096077e-006, 8.238867e-006, 
    8.484738e-006, 8.02628e-006, 7.066395e-006, 4.859532e-006, 2.114743e-006, 
    -4.367761e-006, -5.255621e-006, -6.59077e-006, -7.0686e-006, 
    -7.475897e-006, -4.459904e-006, -1.513399e-008, 3.374382e-006, 
    1.336655e-006, 6.876904e-006, 1.067595e-005, 1.199272e-005, 
    1.483884e-005, 9.45381e-006, 9.134676e-006, 5.206731e-006, 5.826367e-006, 
    8.5878e-006, 1.467592e-005, 2.063067e-005, 1.057065e-005, 8.125372e-006, 
    2.32559e-006, 3.377861e-006, 2.915815e-007, -1.117572e-006, 
    -7.668973e-007, -1.54424e-006, -2.551808e-006, -3.887698e-006, 
    -2.607439e-006, -2.03896e-006, -1.833573e-006, -1.543496e-006, 
    -9.914093e-007, -2.554043e-006, -1.38455e-006, -2.224231e-006, 
    -4.254758e-006, -3.49853e-006, -2.635008e-006,
  2.727068e-007, -3.352607e-007, -1.013263e-006, -9.690564e-007, 
    -6.504199e-007, -1.22635e-006, -1.183633e-006, -9.347838e-007, 
    -4.281443e-007, -5.836134e-007, 9.228952e-007, 7.820781e-007, 
    3.983735e-007, -3.450538e-008, -2.468611e-006, -1.580749e-006, 
    -2.282097e-006, 2.061343e-006, 5.360958e-006, 1.233048e-005, 
    4.288323e-006, -3.638211e-007, 2.198432e-006, 8.121278e-007, 
    -6.685495e-007, -9.03492e-007, -9.313071e-007, -3.186206e-007, 
    -4.882459e-007, -2.433708e-007, 3.286963e-006, 2.516823e-006, 
    3.85296e-006, 3.92796e-006, 1.605552e-005, 1.719645e-005, 7.267308e-006, 
    6.442531e-006, 5.059703e-006, 5.151842e-006, 1.906123e-006, 
    -2.110837e-007, -8.024108e-007, 3.652349e-008, -1.994751e-006, 
    -2.205604e-006, -1.50053e-006, -2.055349e-006, -1.503509e-006, 
    -1.366668e-006, -1.329663e-006, -5.063748e-007, 1.760836e-006, 
    1.404947e-006, -9.213727e-007, -2.700321e-006, -3.49356e-006, 
    -5.387747e-006, -5.351736e-006, -1.262524e-005, -1.384664e-005, 
    -1.37771e-005, -1.545025e-005, -1.244617e-005, -1.082418e-005, 
    -9.382249e-006, -1.197539e-006, 4.16092e-006, 4.700587e-006, 
    4.219528e-006, 5.756085e-006, 7.75632e-006, 3.621495e-006, 1.853721e-006, 
    2.866749e-006, -2.669622e-007, 1.59295e-006, 8.188331e-007, 
    -3.290513e-007, -3.901464e-007, -4.172152e-007, -5.313086e-008, 
    -1.666294e-007, -5.48097e-007, -8.982743e-007, -1.508726e-006, 
    -8.95544e-007, -1.611297e-006, -1.178914e-006, -1.285706e-006, 
    -8.185547e-007, -5.540594e-007, 4.596041e-008, 2.034158e-007, 
    5.891079e-007, 7.666804e-007,
  -3.014844e-007, -3.084383e-007, -2.312006e-007, -2.716821e-007, 
    -1.887323e-007, -9.485495e-008, -2.334359e-007, -3.054581e-007, 
    -1.435321e-007, -4.369431e-008, -2.843478e-007, -7.076483e-008, 
    7.625999e-008, -1.087627e-007, -1.792842e-006, -1.54598e-006, 
    -2.832943e-006, -1.665685e-006, 8.185862e-007, 4.19196e-006, 
    9.688397e-007, -1.738454e-006, 1.664724e-006, 9.628789e-007, 
    -2.382649e-008, -2.020086e-006, -9.062232e-007, -5.168058e-007, 
    -1.613283e-006, -7.184681e-007, 2.747543e-006, 2.622374e-006, 
    1.783686e-006, 3.754612e-006, 9.540234e-006, 8.837896e-006, 
    4.843142e-006, 2.902267e-006, 5.491256e-007, 6.514465e-007, 
    -2.917986e-007, 4.778476e-007, -2.682045e-007, -5.468555e-007, 
    -1.511707e-006, -2.004935e-006, -2.440545e-006, -3.304069e-006, 
    -2.382184e-006, -2.260739e-006, -2.739066e-006, -3.679826e-006, 
    -3.611033e-006, -2.758685e-006, -1.160535e-006, -2.451972e-006, 
    -5.044027e-006, -1.069306e-005, -9.239448e-006, -7.730703e-006, 
    -1.139838e-005, -1.096624e-005, -1.262871e-005, -1.084555e-005, 
    -1.333727e-005, -1.310208e-005, -9.400133e-006, -3.61451e-006, 
    2.535697e-006, 3.137455e-006, 6.388643e-006, 2.962366e-006, 
    9.129601e-007, -1.14787e-006, 4.619533e-007, 6.107166e-007, 5.79671e-007, 
    1.129026e-006, -1.455192e-007, 7.835715e-007, -1.760654e-007, 
    -6.228529e-007, -1.207722e-006, -1.385295e-006, -1.282726e-006, 
    -1.616511e-006, -1.224362e-006, -1.57007e-006, -1.597638e-006, 
    -1.137688e-006, -5.202832e-007, -3.789705e-007, -4.090211e-007, 
    -4.865072e-007, -4.798017e-007, -3.894013e-007,
  -6.33532e-007, -5.339426e-007, -5.520723e-007, -7.127566e-007, 
    -4.728478e-007, -5.858483e-007, -2.550425e-007, -3.782254e-007, 
    -2.235016e-007, -6.579768e-008, 3.751703e-008, -9.775931e-010, 
    6.111048e-008, 1.271723e-007, -1.857521e-007, -9.90912e-007, 
    -8.647485e-007, -2.158026e-007, -5.511851e-008, 1.460471e-007, 
    2.034769e-006, -1.6489e-007, 9.7629e-007, 1.73153e-006, 1.244263e-006, 
    -9.792388e-007, -6.936336e-007, 4.400963e-007, -1.100931e-006, 
    5.066559e-007, 2.282874e-006, 3.312296e-006, 1.845772e-006, 5.89392e-006, 
    5.685307e-006, 4.814829e-006, 2.570218e-006, 1.129772e-006, 
    6.648588e-007, 4.224648e-007, -9.042351e-007, -1.099937e-006, 
    5.901029e-007, 1.887647e-007, -2.198899e-006, -2.818042e-006, 
    -2.862993e-006, -3.040317e-006, -2.018843e-006, -7.005847e-007, 
    -1.85344e-006, -1.693998e-006, -1.700951e-006, -4.999323e-006, 
    -2.545601e-006, -6.588634e-007, -2.627403e-007, -1.048121e-005, 
    -1.398199e-005, -8.445464e-006, -8.323275e-006, -1.051424e-005, 
    -1.14858e-005, -1.015835e-005, -1.015438e-005, -7.43194e-006, 
    -9.813393e-006, -1.513683e-005, -6.282563e-006, -1.81743e-006, 
    1.534981e-007, -1.01525e-006, -1.601114e-006, -1.167242e-006, 
    1.828141e-006, 1.248984e-006, 8.292664e-007, 9.98396e-007, 1.208998e-006, 
    -1.984163e-007, -1.388116e-007, -1.552035e-007, -2.152456e-006, 
    -2.333504e-006, -2.506855e-006, -2.058083e-006, -2.356106e-006, 
    -1.802528e-006, -1.475447e-006, -1.247211e-006, -7.383366e-007, 
    -1.076841e-006, -3.672979e-007, -8.446316e-007, -1.285706e-006, 
    -9.439727e-007,
  -1.310293e-006, -1.193567e-006, -4.485091e-007, -2.642314e-007, 
    -7.058024e-007, -7.716161e-007, -7.346114e-007, -5.046369e-007, 
    -2.307039e-007, -2.148093e-007, -7.904908e-007, -2.135676e-007, 
    -2.220115e-007, 6.930611e-008, 5.142471e-008, -3.04713e-007, 
    -8.73192e-007, -5.834715e-008, -1.134814e-007, 8.718757e-008, 
    9.641209e-007, 1.99851e-006, 2.181794e-006, 1.64262e-006, 1.586493e-006, 
    6.516934e-007, 2.164162e-006, 5.389411e-007, -8.997631e-007, 
    -1.692756e-006, -8.411544e-007, 1.513727e-006, 2.832725e-006, 
    -6.628397e-007, -3.213518e-007, 2.209114e-006, 2.445545e-006, 
    1.059986e-006, -1.577272e-006, -2.281598e-006, -2.23888e-006, 
    -2.62383e-006, -1.61651e-006, -9.833002e-008, -3.285541e-007, 
    -2.056096e-006, -2.133086e-006, -3.106626e-006, -2.642704e-006, 
    -2.120667e-006, -2.152207e-006, -1.418823e-006, -4.142357e-007, 
    -1.801782e-006, -2.715722e-006, -2.596016e-006, -5.927996e-007, 
    -3.553163e-006, -8.137504e-006, -2.948174e-006, -4.36255e-006, 
    -5.867316e-006, -1.01581e-005, -9.94502e-006, -8.359289e-006, 
    -6.829435e-006, -6.05507e-006, -7.230526e-006, -6.620569e-006, 
    -5.782628e-006, -3.625188e-006, -9.775013e-007, 1.117751e-007, 
    -5.51825e-007, 1.178694e-006, 1.427545e-006, 2.814595e-006, 
    1.540298e-006, 1.266762e-007, -4.355943e-007, -1.4139e-008, 
    7.445778e-007, -2.321832e-006, -2.821271e-006, -3.552172e-006, 
    -2.038213e-006, -2.867711e-006, -2.61489e-006, -1.606081e-006, 
    -1.065666e-006, -1.147232e-007, -7.646621e-007, -8.272469e-007, 
    -8.218899e-008, -8.299789e-007, -1.222625e-006,
  -1.325443e-006, -1.845741e-006, -1.50674e-006, -4.713575e-007, 
    -3.357569e-007, -6.3229e-007, -9.154122e-007, -1.001342e-006, 
    -7.579566e-007, -3.779771e-007, -6.464463e-007, -1.092594e-007, 
    -3.732584e-007, -9.956302e-007, -2.85838e-007, 2.669949e-007, 
    -2.092356e-006, -8.277435e-007, 3.329495e-008, 8.520075e-008, 
    4.969695e-007, 9.34567e-007, 2.162422e-006, 3.097719e-006, 2.539423e-006, 
    8.06665e-007, 9.636242e-007, 1.8947e-006, 9.344783e-006, 2.461311e-007, 
    -1.039094e-006, -2.377217e-006, -3.223849e-006, -8.345374e-006, 
    -7.669858e-006, -6.05855e-006, -3.490333e-006, -2.483357e-007, 
    7.302879e-008, 1.840453e-007, -6.243445e-007, -1.133712e-006, 
    -3.226333e-006, -2.532434e-006, -2.306931e-006, -4.185968e-006, 
    -3.535782e-006, -3.529075e-006, -3.008528e-006, -1.35425e-006, 
    -2.826485e-006, -4.302941e-006, -4.145983e-006, -4.546329e-006, 
    -5.975848e-006, -7.12423e-006, -6.083137e-006, -2.165871e-006, 
    -1.437447e-006, 5.838901e-007, 4.559897e-007, -4.733447e-007, 
    -4.821502e-006, -8.08312e-006, -6.078914e-006, -4.982438e-006, 
    -5.534524e-006, -4.511061e-006, -6.344651e-006, -9.388712e-006, 
    -5.621694e-006, 2.545748e-007, 2.519057e-006, 3.720337e-006, 
    7.223105e-006, 5.905593e-006, 1.919534e-006, 1.013792e-006, 
    3.329182e-006, -9.411087e-008, -1.581991e-006, -2.245092e-006, 
    -2.272163e-006, -2.752227e-006, -3.502255e-006, -2.949668e-006, 
    -1.366171e-006, -2.564225e-006, -1.595899e-006, -1.523876e-006, 
    -7.51003e-007, -6.819608e-007, -8.034051e-007, -5.488436e-007, 
    -1.497407e-007, -1.31973e-006,
  -6.305515e-007, -9.623508e-007, -1.483892e-006, -1.534059e-006, 
    -1.160537e-006, -9.807291e-007, -1.501276e-006, -1.401935e-006, 
    -1.113597e-006, -7.452908e-007, -1.038843e-006, -9.544035e-007, 
    -2.398931e-007, -2.148732e-006, -4.665786e-006, -4.114444e-006, 
    -4.115436e-006, -3.87975e-006, -2.255275e-006, -1.231565e-006, 
    1.428184e-007, 1.337644e-006, 7.334011e-007, -7.498716e-008, 
    7.731373e-007, 9.950268e-006, 2.479818e-006, 2.518311e-006, 
    5.612786e-006, 4.867976e-006, -1.137305e-007, -7.423077e-007, 
    1.211232e-006, -4.133071e-006, -8.349354e-006, -1.231107e-005, 
    -1.472406e-005, -1.262996e-005, -1.093644e-005, -5.937851e-006, 
    -2.584587e-006, -1.602109e-006, -7.564686e-007, -1.905844e-006, 
    -3.713852e-006, -3.160772e-006, -3.402416e-006, -3.098929e-006, 
    -4.675225e-006, -5.265065e-006, -4.880614e-006, -3.30283e-006, 
    -2.916144e-006, -3.45035e-006, -5.359932e-006, -4.769841e-006, 
    8.988027e-007, 1.204775e-006, -2.389386e-006, -1.178172e-006, 
    2.64261e-007, -1.823639e-006, -3.460033e-006, -5.371854e-006, 
    -5.039807e-006, -3.119542e-006, -3.436192e-006, -5.75829e-006, 
    -4.961572e-006, -5.367383e-006, -5.549176e-006, -2.447745e-006, 
    -7.532326e-007, 2.887864e-006, 9.189565e-006, 9.714826e-006, 
    6.499155e-006, 3.98856e-006, 2.118213e-006, 1.746183e-006, 1.492119e-006, 
    2.322609e-006, 1.402708e-006, -1.819168e-006, -3.704661e-006, 
    -5.545589e-007, 9.387886e-007, -8.346979e-007, -7.383351e-007, 
    -8.982752e-007, -1.978362e-006, -1.219397e-006, -1.208965e-006, 
    -1.296882e-006, -4.569529e-007, -4.457772e-007,
  -1.36965e-006, -7.028225e-007, -9.15413e-007, -1.045053e-006, 
    -7.706226e-007, -1.41932e-006, -2.319847e-006, -2.897266e-006, 
    -2.920363e-006, -3.728752e-006, -3.12898e-006, -2.040698e-006, 
    -1.606826e-006, -3.737444e-006, -3.926687e-006, -3.401422e-006, 
    -4.110221e-006, -6.334716e-006, -9.00724e-006, -4.828954e-006, 
    -2.781782e-006, -2.358588e-006, -1.214266e-007, 1.875223e-007, 
    -6.635826e-007, -1.455579e-006, -2.523093e-007, 3.357497e-006, 
    5.237279e-006, 7.249928e-006, 4.861522e-006, 3.15435e-006, 4.819594e-008, 
    3.203932e-007, -4.358408e-007, 1.541412e-008, -4.156409e-006, 
    -7.97235e-006, -1.238906e-005, -1.255023e-005, -1.410194e-005, 
    -1.254104e-005, -6.692837e-006, -5.309761e-006, -1.81072e-006, 
    8.449169e-007, 4.987123e-007, -6.203663e-007, 1.604603e-007, 
    -2.710753e-006, -3.372115e-006, -2.282843e-006, -4.178513e-006, 
    -1.657976e-006, 3.507997e-006, 3.12852e-006, 1.716635e-006, 
    9.261239e-007, 3.945344e-006, 3.323968e-006, 2.804414e-006, 5.27516e-007, 
    -2.25602e-006, -2.016361e-006, -3.024425e-006, -2.322827e-006, 
    -4.04267e-006, -5.082026e-006, -5.669876e-006, -4.897251e-006, 
    -3.880246e-006, -4.660076e-006, -6.320057e-006, -6.312614e-006, 
    2.232846e-007, 1.010747e-005, 1.432202e-005, 5.65749e-006, 
    -2.655725e-008, -2.030021e-006, -1.759807e-006, 8.960342e-009, 
    1.677392e-006, 1.492299e-008, -6.332848e-007, -4.68377e-007, 
    3.904279e-007, 9.132109e-007, 3.211335e-007, -8.51338e-007, 
    -1.263601e-006, -1.829844e-006, -2.329036e-006, -3.348773e-006, 
    -4.454686e-006, -3.435695e-006,
  -2.939735e-006, -2.406768e-006, -4.588795e-006, -5.160506e-006, 
    -2.999341e-006, -2.120421e-006, -3.423529e-006, -3.907564e-006, 
    -5.983298e-006, -6.659313e-006, -3.232292e-006, -3.696465e-006, 
    -4.933014e-006, -5.416804e-006, -3.386021e-006, -5.205311e-007, 
    -5.746697e-007, -1.301598e-006, -4.222478e-006, -3.847465e-006, 
    -1.078579e-006, -7.008357e-007, 3.496971e-007, 1.440603e-007, 
    1.472886e-007, 4.006088e-007, 2.771772e-007, 7.726408e-007, 
    2.454488e-006, 4.456707e-006, 4.765656e-006, 5.424038e-006, 
    6.038958e-006, 6.488477e-006, 7.562852e-006, 8.232164e-006, 
    9.161249e-006, 7.760547e-006, 3.451372e-006, -2.572182e-006, 
    -3.245965e-006, -3.457062e-006, -5.448601e-006, -7.36439e-006, 
    -4.9956e-006, -4.219743e-006, 9.94427e-007, 2.706322e-006, 2.167646e-006, 
    1.473989e-006, 1.417615e-006, 3.583744e-006, 1.021242e-006, 
    -1.303706e-007, 3.216435e-006, 4.227226e-006, -7.194612e-007, 
    -3.285688e-006, -3.772257e-007, 5.303093e-006, 5.327682e-006, 
    3.800555e-006, 1.916305e-006, -1.475699e-006, -2.421422e-006, 
    -1.207226e-006, -2.386496e-007, -4.703625e-007, -5.622551e-007, 
    -5.349357e-007, -2.712741e-006, -1.148865e-006, -3.916008e-006, 
    -9.675678e-007, -2.110828e-007, 2.024834e-006, 9.110339e-006, 
    9.785603e-006, 1.138749e-005, -1.274529e-006, -6.390852e-006, 
    -3.429741e-006, -2.628789e-006, -3.45608e-009, 1.899665e-006, 
    2.214576e-006, 2.128148e-006, 1.312317e-006, -1.547465e-006, 
    1.416993e-008, 1.507018e-006, -1.25193e-006, -1.168484e-006, 
    -2.556526e-006, -6.492669e-006, -4.484737e-006,
  -2.678466e-006, -3.726269e-006, -3.242478e-006, -4.877882e-006, 
    -2.716717e-006, -3.055467e-006, -1.217164e-006, -2.480282e-006, 
    -5.195521e-006, -6.439275e-006, -3.039819e-006, -1.678352e-006, 
    -2.836014e-007, 9.201631e-007, 1.22207e-007, 2.758497e-008, 
    -3.824462e-007, -8.923053e-009, 1.795111e-006, 2.776724e-007, 
    1.77549e-006, 1.352048e-006, 8.667666e-007, 1.40743e-006, 1.00634e-006, 
    1.020745e-006, 1.218682e-006, 5.138575e-007, 9.566704e-007, 
    1.677887e-006, 1.675651e-006, 1.575565e-006, 1.88998e-006, 3.093746e-006, 
    3.598398e-006, 2.690173e-006, -2.443769e-006, 4.45819e-006, 
    6.667538e-006, 7.449602e-006, 1.06248e-005, 1.16865e-005, 1.002203e-005, 
    6.553048e-006, 6.034737e-006, 4.862508e-006, 6.31711e-006, 5.927934e-006, 
    2.639747e-006, 3.166759e-006, 7.302326e-006, 1.091288e-005, 
    9.911029e-006, 6.487986e-006, 9.852916e-006, 9.382038e-006, 
    8.108978e-006, 4.951424e-006, 3.383822e-006, 4.091133e-006, 
    6.496677e-006, 2.240908e-006, 2.160938e-006, 6.65438e-006, 4.642479e-006, 
    2.303734e-006, 3.913307e-006, 3.462053e-006, 4.457701e-006, 
    5.902119e-006, 3.665453e-006, 3.233814e-006, 1.338636e-006, 
    -1.718472e-007, 2.126664e-006, 7.075585e-006, 8.213286e-006, 
    6.985181e-006, 6.241866e-006, 5.849717e-006, 2.649693e-006, 9.93663e-007, 
    -9.372743e-007, -6.361537e-006, -4.809328e-006, -3.136171e-006, 
    1.85621e-006, 2.677258e-006, -7.810522e-007, -5.82615e-007, 
    1.494107e-006, 2.52129e-006, 7.726376e-007, 9.948053e-009, 
    -2.974752e-006, -3.600604e-006,
  3.925379e-008, -2.407342e-008, -6.695427e-007, -2.983696e-006, 
    -7.470317e-007, 2.841316e-007, 4.741196e-007, -6.059636e-007, 
    -6.990949e-007, -6.963655e-007, 1.330191e-006, 2.00596e-006, 
    -1.693606e-007, 1.987833e-006, 2.255557e-006, 1.757361e-006, 
    4.957278e-007, 1.142687e-006, 2.719479e-006, 2.814102e-006, 
    3.325708e-006, 2.117967e-006, 8.77694e-007, 3.12195e-007, 2.073904e-007, 
    3.462195e-007, 4.040857e-007, 3.900743e-008, 3.87588e-008, 2.6625e-007, 
    6.235223e-008, -1.122398e-007, -8.367897e-008, 3.410041e-007, 
    1.138961e-006, 1.049802e-006, -4.683743e-007, 1.933695e-006, 
    4.022339e-006, 5.602107e-006, 5.775957e-006, 5.602109e-006, 
    6.678965e-006, 5.877777e-006, 6.236649e-006, 6.071998e-006, 
    4.063317e-006, 6.11024e-006, 6.173323e-006, 6.33052e-006, 6.427385e-006, 
    9.884952e-006, 1.083912e-005, 9.165971e-006, 1.38129e-005, 1.330923e-005, 
    1.366215e-005, 8.746996e-006, 6.566956e-006, 2.60002e-006, 3.402201e-006, 
    4.721704e-006, 5.75485e-006, 5.377849e-006, 6.880135e-006, 8.307168e-006, 
    6.445511e-006, 4.341222e-006, 4.705059e-006, 4.20885e-006, 5.448131e-006, 
    5.770737e-006, 4.685187e-006, 2.604489e-006, 3.950809e-006, 
    5.044061e-006, 9.515654e-006, 1.217799e-005, 1.235159e-005, 
    8.452451e-006, 1.886503e-006, 1.904384e-006, -1.011278e-006, 
    -2.595767e-006, -3.065648e-006, -5.865822e-006, -5.672104e-006, 
    -2.506105e-006, 1.260654e-006, 4.798196e-006, 6.351391e-006, 
    5.756086e-006, 3.906851e-006, 2.817578e-006, 3.381589e-006, -4.395697e-007,
  4.31266e-006, 3.236546e-006, 2.965351e-006, 1.512979e-006, 5.687416e-007, 
    9.314681e-008, 5.861275e-007, 1.494355e-006, 5.381962e-007, 5.25034e-007, 
    3.434735e-006, 3.696248e-006, 4.777327e-006, 3.789631e-006, 
    3.692775e-006, 1.836334e-006, 1.324232e-006, 1.719858e-006, 
    9.983928e-007, 2.130882e-006, 2.537434e-006, 2.535199e-006, 
    2.044703e-006, 1.362479e-006, 1.272575e-006, 7.845613e-007, 
    6.069895e-007, 2.441466e-007, 1.984499e-007, 3.151752e-007, 
    8.133708e-007, 7.140299e-007, 6.131986e-007, 4.929957e-007, 
    3.946477e-007, 6.027674e-007, 7.36381e-007, -1.116579e-006, 
    7.475537e-007, 2.908473e-006, 1.971934e-006, 3.616224e-007, 
    1.790639e-006, 3.859914e-006, 3.94907e-006, 3.110883e-006, 2.299264e-006, 
    2.485282e-006, 3.273057e-006, 3.969686e-006, 6.029277e-006, 
    2.966837e-006, 8.642939e-006, 8.175288e-006, 1.069979e-005, 9.91649e-006, 
    8.632505e-006, 8.592026e-006, 8.996591e-006, 4.678735e-006, 
    3.435733e-006, 6.824921e-007, 1.662742e-006, 4.4505e-006, 7.880248e-006, 
    7.726518e-006, 3.712143e-006, 2.531973e-006, 3.371158e-006, 
    3.872083e-006, 5.377101e-006, 5.265342e-006, 4.845874e-006, 
    6.391867e-006, 6.050881e-006, 3.84948e-006, 6.486987e-006, 9.144613e-006, 
    1.068887e-005, 9.538497e-006, 6.817547e-006, 2.734134e-006, 
    2.461442e-006, -1.547218e-006, -1.005064e-006, -1.406403e-006, 
    -4.413705e-006, -6.369984e-006, -7.806448e-006, -3.141897e-006, 
    -1.47197e-006, 8.789393e-007, 6.486494e-006, 8.161878e-006, 
    6.777318e-006, 6.77259e-006,
  5.846485e-006, 7.545714e-006, 8.16138e-006, 5.806998e-006, 4.081941e-006, 
    5.579011e-006, 4.641729e-006, 2.98472e-006, 4.067786e-006, 2.412515e-006, 
    2.449024e-006, 3.09027e-006, 3.130008e-006, 2.422943e-006, 2.203651e-006, 
    3.14615e-006, 3.46106e-006, 2.954419e-006, 2.187258e-006, 1.580035e-006, 
    1.62449e-006, 2.115483e-006, 2.332048e-006, 1.887496e-006, 1.715635e-006, 
    1.4648e-006, 1.047568e-006, 1.040862e-006, 1.323239e-006, 1.156594e-006, 
    7.579881e-007, 7.284341e-007, 1.078612e-006, 6.482161e-007, 6.41511e-007, 
    1.25072e-006, 9.887076e-007, 1.60959e-006, 2.825029e-006, 4.405793e-006, 
    6.260738e-006, 4.376734e-006, 4.2836e-006, 5.267326e-006, 3.806515e-006, 
    3.068417e-006, 3.20873e-006, 4.717975e-006, 6.055852e-006, 7.782895e-006, 
    6.992883e-006, 2.642242e-006, 3.344088e-006, 4.65415e-006, 8.500134e-006, 
    8.294253e-006, 6.697341e-006, 6.390375e-006, 8.529936e-006, 
    7.203489e-006, 6.356855e-006, 4.883375e-006, 3.670175e-006, 
    5.180402e-006, 6.946189e-006, 4.538164e-006, 3.412136e-006, 
    1.559422e-006, 1.951818e-006, 3.13373e-006, 3.698735e-006, 3.914553e-006, 
    3.911572e-006, 3.876058e-006, 5.027421e-006, 5.436706e-006, 
    6.975994e-006, 7.718816e-006, 8.135801e-006, 8.133564e-006, 
    7.096443e-006, 6.837168e-006, 6.591301e-006, 2.947221e-006, 
    1.931956e-006, -5.693437e-009, -3.745139e-006, -8.553248e-006, 
    -1.051275e-005, -5.149577e-006, -7.225026e-008, 1.113633e-006, 
    3.93964e-006, 7.226332e-006, 8.729869e-006, 7.462517e-006,
  3.634905e-006, 3.617022e-006, 3.433737e-006, 3.586974e-006, 3.797578e-006, 
    3.665951e-006, 3.135469e-006, 4.271434e-006, 6.500149e-006, 
    6.178287e-006, 2.763935e-006, 2.385693e-006, 1.988825e-006, 
    2.926358e-006, 3.921259e-006, 4.938014e-006, 3.094741e-006, 
    2.199676e-006, 3.582751e-006, 2.929336e-006, 1.32001e-006, 1.661495e-006, 
    3.507007e-006, 4.010417e-006, 2.851602e-006, 2.108282e-006, 
    2.265489e-006, 2.484038e-006, 2.114987e-006, 1.744693e-006, 
    1.611328e-006, 1.527633e-006, 1.096492e-006, 1.142686e-006, 1.23855e-006, 
    1.549736e-006, 8.175925e-007, 1.216447e-006, 3.268092e-006, 9.26059e-006, 
    1.248471e-005, 5.703683e-006, 1.837578e-006, 1.444929e-006, 
    9.852338e-007, 2.343226e-006, 1.699245e-006, 2.382216e-006, 
    6.119571e-007, 3.056495e-006, 3.508745e-006, 4.64396e-006, 6.518037e-006, 
    5.431491e-006, 7.273025e-006, 7.337845e-006, 6.225473e-006, 
    5.339602e-006, 6.398826e-006, 7.194296e-006, 1.022022e-005, 
    1.299234e-005, 1.341454e-005, 7.874038e-006, 5.923475e-006, 
    4.021592e-006, 3.185639e-006, 1.563644e-006, 7.718954e-007, 
    7.830713e-007, 1.100218e-006, 2.255309e-006, 2.789017e-006, 
    2.575185e-006, 3.12479e-006, 4.037486e-006, 5.370644e-006, 6.017355e-006, 
    5.159296e-006, 6.263965e-006, 5.56982e-006, 3.254429e-006, 6.021075e-006, 
    4.324582e-006, -3.963578e-007, -9.961259e-007, -7.996787e-007, 
    -2.195913e-006, -6.033708e-006, -6.625782e-006, -3.685287e-006, 
    -1.974633e-006, 4.448193e-007, 5.191338e-006, 2.851357e-006, 1.837578e-006,
  2.328074e-006, 3.940875e-006, 5.174443e-006, 6.993627e-006, 7.998711e-006, 
    7.328902e-006, 3.802546e-006, 3.986823e-006, 6.533181e-006, 
    5.055977e-006, 3.024456e-006, 2.307213e-006, 2.862532e-006, 
    3.231085e-006, 3.43399e-006, 4.259017e-006, 4.454473e-006, 3.729032e-006, 
    3.432251e-006, 2.384201e-006, 2.304232e-006, 2.502416e-006, 
    2.284612e-006, 1.543776e-006, 1.313056e-006, 2.162424e-006, 
    2.319134e-006, 1.098479e-006, 5.493721e-007, 8.508719e-007, 
    9.519522e-007, 1.069174e-006, 1.134987e-006, 1.086807e-006, 
    1.067932e-006, 1.669194e-006, 1.767293e-006, 1.767789e-006, 
    3.176694e-006, 5.190092e-006, 5.284218e-006, 2.620139e-006, 
    1.760838e-006, 2.291816e-006, 2.866127e-007, -1.770604e-007, 
    2.168385e-006, 4.751004e-006, 7.026159e-006, 5.97538e-006, 4.724179e-006, 
    4.24188e-006, 3.910081e-006, 4.562751e-006, 5.979851e-006, 6.61489e-006, 
    9.19776e-006, 1.043902e-005, 1.089326e-005, 1.513612e-005, 1.883533e-005, 
    1.58315e-005, 8.910911e-006, 4.310425e-006, 3.70097e-006, 2.871472e-006, 
    2.076988e-006, 2.118217e-006, 2.446044e-006, 1.438475e-006, 
    1.646594e-006, 1.853968e-006, 1.576806e-006, 1.685833e-006, 
    1.953061e-006, 2.341981e-006, 4.236914e-006, 5.137192e-006, 
    2.956656e-006, 3.592686e-006, 6.022568e-006, 5.069142e-006, 2.48677e-006, 
    -1.213684e-006, -5.173168e-006, -2.771598e-006, 4.492867e-007, 
    -6.198716e-007, -1.860146e-006, -4.497149e-006, -1.124521e-006, 
    4.123172e-006, 5.425532e-006, 5.600621e-006, 6.087635e-006, 3.578776e-006,
  4.843389e-006, 3.695503e-006, 5.435462e-006, 5.539523e-006, 3.551457e-006, 
    2.441073e-006, 3.189113e-006, 2.866505e-006, 2.436108e-006, 
    2.359368e-006, 2.227493e-006, 2.530731e-006, 3.197807e-006, 
    3.601131e-006, 2.384949e-006, 1.616792e-006, 2.056377e-006, 
    2.170123e-006, 2.305227e-006, 2.203649e-006, 2.301996e-006, 
    2.195455e-006, 1.448906e-006, 1.417862e-006, 1.579787e-006, 1.95033e-006, 
    1.619524e-006, 1.312063e-006, 8.543484e-007, 1.006837e-006, 
    1.456107e-006, 1.133498e-006, 9.551804e-007, 9.010391e-007, 1.46331e-006, 
    1.623497e-006, 1.037136e-006, 1.555945e-006, 2.808387e-006, 3.92051e-006, 
    3.150121e-006, 2.236928e-006, 2.344962e-006, 2.076744e-006, 4.84305e-007, 
    -1.27885e-007, 7.423423e-007, 1.980629e-006, 3.150121e-006, 
    5.364184e-006, 5.24125e-006, 3.012784e-006, 1.847015e-006, 4.406289e-006, 
    6.077205e-006, 5.715356e-006, 8.778787e-006, 1.197061e-005, 
    1.375751e-005, 1.478445e-005, 1.382854e-005, 6.542617e-006, 
    2.541907e-006, 1.471009e-006, 1.015034e-006, 1.386817e-006, 
    1.841302e-006, 2.415992e-006, 3.278273e-006, 1.702224e-006, 
    9.889559e-007, 1.324729e-006, 2.183533e-006, 2.021109e-006, 
    1.377876e-006, 1.03962e-006, 2.125169e-006, 3.094987e-006, 3.186629e-006, 
    3.610817e-006, 2.717245e-006, 3.417508e-007, 1.839544e-008, 
    4.855465e-007, 9.598971e-007, 8.312491e-007, 2.136097e-006, 
    2.979006e-006, 1.827397e-006, 3.656016e-006, 3.411888e-006, 
    1.842543e-006, -1.9123e-006, -1.336368e-006, 4.908215e-006, 6.957858e-006,
  -1.450857e-006, -6.019909e-007, 1.611326e-006, 4.494206e-006, 
    5.161034e-006, 3.687805e-006, 3.5455e-006, 3.404931e-006, 2.356636e-006, 
    1.779961e-006, 1.288967e-006, 1.789151e-006, 1.977402e-006, 
    1.902896e-006, 1.749413e-006, 1.629955e-006, 2.160188e-006, 
    2.986707e-006, 2.790509e-006, 1.931703e-006, 1.727309e-006, 1.87185e-006, 
    1.243767e-006, 9.901978e-007, 1.227623e-006, 1.53558e-006, 1.317278e-006, 
    8.161028e-007, 7.771114e-007, 8.441666e-007, 1.053776e-006, 
    1.181926e-006, 1.106675e-006, 1.133497e-006, 1.120583e-006, 
    1.024222e-006, 1.172737e-006, 1.046326e-006, 1.409914e-006, 
    2.630071e-006, 3.64012e-006, 3.271814e-006, 1.985844e-006, 1.071409e-006, 
    1.233584e-006, 1.41215e-006, 1.200307e-006, 1.338141e-006, 1.543776e-006, 
    1.633683e-006, 8.183397e-007, 1.016027e-006, 1.488146e-006, 
    1.676151e-006, 2.374518e-006, 3.856686e-006, 4.562505e-006, 
    4.852829e-006, 4.394618e-006, 3.326703e-006, 2.424435e-006, 1.49485e-006, 
    1.001869e-006, 7.87541e-007, 6.506989e-007, 8.528586e-007, 1.44369e-006, 
    2.460693e-006, 1.654044e-006, 1.396751e-006, 8.267816e-007, 
    1.084324e-006, 1.233831e-006, 1.454121e-006, 1.134739e-006, 
    7.515309e-007, 1.059985e-006, 2.043462e-006, 1.92003e-006, 1.470512e-006, 
    8.83655e-007, 4.035892e-007, 7.562512e-007, 4.713911e-007, 1.383836e-006, 
    -3.640707e-007, -4.567937e-006, -5.645536e-006, -1.355493e-006, 
    1.886008e-006, 7.912677e-007, -2.843481e-007, 4.430767e-007, 
    1.982862e-006, 2.537186e-006, 4.242065e-007,
  -1.61577e-006, -3.350511e-006, -3.321453e-006, -2.459423e-006, 
    -1.327679e-006, 7.477047e-008, 7.428398e-007, 1.441952e-006, 
    2.235688e-006, 1.88129e-006, 1.658516e-006, 2.437848e-006, 3.35849e-006, 
    3.208485e-006, 2.614425e-006, 2.280639e-006, 1.907364e-006, 2.13709e-006, 
    2.123183e-006, 1.837577e-006, 1.440461e-006, 8.816678e-007, 
    7.507861e-007, 1.493609e-006, 1.895941e-006, 1.937662e-006, 1.16628e-006, 
    9.459909e-007, 9.184239e-007, 1.068677e-006, 1.332925e-006, 
    1.268849e-006, 1.147405e-006, 9.452458e-007, 8.74217e-007, 8.054235e-007, 
    1.101957e-006, 2.037998e-006, 2.480313e-006, 1.983609e-006, 
    1.346087e-006, 1.240537e-006, 1.870856e-006, 2.189493e-006, 
    1.946106e-006, 2.535696e-006, 2.606725e-006, 1.74668e-006, 1.463806e-006, 
    1.768535e-006, 1.505033e-006, 1.674409e-006, 1.880294e-006, 
    1.929964e-006, 1.84304e-006, 2.350674e-006, 2.025579e-006, 1.702474e-006, 
    1.433507e-006, 9.651139e-007, 1.254942e-006, 1.487152e-006, 
    1.397744e-006, 1.204774e-006, 7.711506e-007, 8.07659e-007, 5.081451e-007, 
    9.427624e-007, 1.223152e-006, 1.605367e-006, 1.853968e-006, 
    1.918788e-006, 1.867875e-006, 1.863902e-006, 1.7437e-006, 1.533345e-006, 
    1.184906e-006, 1.294678e-006, 9.283576e-007, 4.204762e-007, 
    7.098074e-007, 1.453127e-006, 1.694278e-006, 8.911061e-007, 
    4.743706e-007, -7.589488e-007, -2.205107e-006, -1.951539e-006, 
    -2.014003e-007, 9.854775e-007, 1.134988e-006, 1.404949e-006, 
    3.276282e-006, 1.575068e-006, 8.324951e-007, 6.497066e-007,
  8.178431e-007, 7.24458e-007, -1.234794e-006, -3.603582e-006, -4.13779e-006, 
    -3.539259e-006, -1.407152e-006, 1.544522e-006, 3.78044e-006, 
    3.775971e-006, 3.218421e-006, 3.014025e-006, 2.600269e-006, 
    2.000746e-006, 1.683848e-006, 1.588479e-006, 1.302625e-006, 
    1.385327e-006, 1.568362e-006, 1.397248e-006, 1.401469e-006, 
    1.566872e-006, 2.056624e-006, 2.26673e-006, 1.970446e-006, 1.572833e-006, 
    1.122321e-006, 1.011556e-006, 7.480539e-007, 7.584849e-007, 
    8.928437e-007, 1.121328e-006, 1.081592e-006, 1.158333e-006, 
    1.479701e-006, 1.454121e-006, 1.646842e-006, 1.60636e-006, 9.946682e-007, 
    9.693363e-007, 1.341865e-006, 1.882281e-006, 2.1356e-006, 2.335772e-006, 
    2.063578e-006, 1.688814e-006, 1.83559e-006, 2.01192e-006, 2.172108e-006, 
    2.19446e-006, 1.95927e-006, 1.636411e-006, 1.195337e-006, 1.186148e-006, 
    9.869693e-007, 9.554285e-007, 1.336898e-006, 1.552468e-006, 
    1.400476e-006, 1.132752e-006, 7.281853e-007, 7.552562e-007, 
    9.613889e-007, 1.119838e-006, 1.354283e-006, 1.230603e-006, 
    1.084075e-006, 1.156843e-006, 1.078115e-006, 1.278038e-006, 
    1.734758e-006, 2.057866e-006, 1.865392e-006, 1.642371e-006, 1.68186e-006, 
    1.964734e-006, 1.948342e-006, 1.615549e-006, 6.529344e-007, 
    6.011692e-008, 1.495239e-007, 3.459711e-007, 1.487792e-007, 
    -3.628284e-007, 2.311162e-008, 4.912574e-007, 6.991286e-007, 
    1.020745e-006, 1.980628e-006, 2.471126e-006, 2.087421e-006, 
    1.955545e-006, 2.284363e-006, 9.603937e-007, -5.063757e-007, 
    -3.640689e-007,
  -1.129243e-006, -3.00739e-007, 3.159203e-007, 2.096258e-007, 2.578072e-007, 
    9.134583e-007, 1.431771e-006, 1.192608e-006, 5.08644e-007, 
    -1.000699e-007, -1.92209e-007, 9.438918e-008, 6.084792e-007, 
    9.673495e-007, 9.34815e-007, 9.368018e-007, 1.217192e-006, 1.412894e-006, 
    1.393771e-006, 1.471753e-006, 1.788651e-006, 2.071773e-006, 
    1.905625e-006, 1.495347e-006, 1.438971e-006, 1.523411e-006, 
    1.479204e-006, 1.403954e-006, 1.201297e-006, 8.680083e-007, 
    7.609683e-007, 7.132846e-007, 7.597266e-007, 8.771972e-007, 
    8.126253e-007, 8.732236e-007, 9.797668e-007, 1.002864e-006, 
    1.074638e-006, 1.206761e-006, 1.248236e-006, 1.254693e-006, 
    1.367694e-006, 1.311318e-006, 1.074638e-006, 8.901118e-007, 
    9.775317e-007, 1.251962e-006, 1.565382e-006, 1.901404e-006, 
    1.934186e-006, 1.695022e-006, 1.41811e-006, 1.285737e-006, 1.226133e-006, 
    1.485661e-006, 1.712904e-006, 1.779214e-006, 1.719858e-006, 1.48293e-006, 
    1.272326e-006, 1.040862e-006, 8.801771e-007, 9.38292e-007, 1.176959e-006, 
    1.309082e-006, 1.11959e-006, 1.104937e-006, 1.382098e-006, 1.81597e-006, 
    1.863902e-006, 1.410908e-006, 1.320755e-006, 1.593447e-006, 
    1.902646e-006, 2.135848e-006, 2.054885e-006, 1.796847e-006, 1.65777e-006, 
    1.407431e-006, 7.425904e-007, -2.714337e-007, -9.439727e-007, 
    -8.798984e-007, -2.207701e-007, 4.311557e-007, 8.84648e-007, 
    1.205023e-006, 1.729792e-006, 2.629078e-006, 3.458079e-006, 
    3.593182e-006, 3.093251e-006, 2.127655e-006, 4.030926e-007, -1.052751e-006,
  2.509869e-006, 1.887745e-006, 1.280274e-006, 1.084571e-006, 1.206761e-006, 
    1.091525e-006, 6.586461e-007, 3.206378e-007, 1.465423e-007, 1.34125e-007, 
    4.47546e-007, 9.862229e-007, 1.521672e-006, 1.857693e-006, 2.061095e-006, 
    2.042965e-006, 1.887992e-006, 1.774495e-006, 1.608844e-006, 
    1.461075e-006, 1.334166e-006, 1.267359e-006, 1.18888e-006, 1.065697e-006, 
    9.710745e-007, 1.058495e-006, 1.207506e-006, 1.332676e-006, 
    1.318024e-006, 1.164541e-006, 1.005099e-006, 9.318351e-007, 
    9.867208e-007, 1.053031e-006, 9.58905e-007, 8.851446e-007, 8.901118e-007, 
    9.62134e-007, 1.083082e-006, 1.111394e-006, 1.040365e-006, 1.037385e-006, 
    1.079605e-006, 1.168267e-006, 1.227126e-006, 1.128778e-006, 
    1.009321e-006, 9.472326e-007, 1.055266e-006, 1.299397e-006, 
    1.449898e-006, 1.442945e-006, 1.330937e-006, 1.186893e-006, 
    1.025216e-006, 9.581604e-007, 9.978967e-007, 1.06222e-006, 1.185403e-006, 
    1.240537e-006, 1.134988e-006, 1.020497e-006, 1.005099e-006, 
    9.884591e-007, 9.785251e-007, 1.032666e-006, 1.137223e-006, 
    1.202788e-006, 1.288966e-006, 1.426802e-006, 1.468525e-006, 
    1.305606e-006, 1.190122e-006, 1.245256e-006, 1.231845e-006, 
    1.155849e-006, 1.104688e-006, 1.085813e-006, 1.020496e-006, 
    9.154433e-007, 8.352258e-007, 6.874559e-007, 5.056618e-007, 
    4.838064e-007, 6.715613e-007, 9.554284e-007, 1.284744e-006, 
    1.783933e-006, 2.312428e-006, 2.601758e-006, 2.557055e-006, 
    2.437597e-006, 2.452251e-006, 2.554323e-006, 2.60921e-006, 2.656645e-006,
  3.286219e-006, 3.084308e-006, 2.796964e-006, 2.420212e-006, 2.055382e-006, 
    1.759097e-006, 1.49783e-006, 1.268352e-006, 1.115368e-006, 1.021987e-006, 
    9.740552e-007, 1.00808e-006, 1.141941e-006, 1.304116e-006, 1.424815e-006, 
    1.477714e-006, 1.441703e-006, 1.440462e-006, 1.517699e-006, 
    1.581774e-006, 1.586741e-006, 1.52962e-006, 1.44667e-006, 1.327213e-006, 
    1.188632e-006, 1.037633e-006, 9.445012e-007, 9.298481e-007, 
    9.579121e-007, 1.0652e-006, 1.193599e-006, 1.258667e-006, 1.253203e-006, 
    1.21744e-006, 1.183913e-006, 1.177456e-006, 1.178946e-006, 1.177207e-006, 
    1.161313e-006, 1.129275e-006, 1.117603e-006, 1.156594e-006, 
    1.210983e-006, 1.262889e-006, 1.301135e-006, 1.317775e-006, 
    1.316782e-006, 1.289711e-006, 1.213467e-006, 1.15411e-006, 1.112387e-006, 
    1.072402e-006, 1.009569e-006, 9.422658e-007, 9.055098e-007, 
    9.216526e-007, 9.440043e-007, 9.363055e-007, 9.137054e-007, 
    9.402791e-007, 1.00187e-006, 1.048312e-006, 1.091774e-006, 1.158581e-006, 
    1.265373e-006, 1.336402e-006, 1.312063e-006, 1.24923e-006, 1.167025e-006, 
    1.067932e-006, 1.004354e-006, 9.901978e-007, 1.028444e-006, 
    1.116113e-006, 1.207258e-006, 1.241779e-006, 1.222904e-006, 
    1.186148e-006, 1.147902e-006, 1.12108e-006, 1.159326e-006, 1.265869e-006, 
    1.390046e-006, 1.466042e-006, 1.481688e-006, 1.517202e-006, 
    1.574075e-006, 1.630699e-006, 1.66373e-006, 1.691049e-006, 1.805539e-006, 
    2.060845e-006, 2.475346e-006, 2.901769e-006, 3.213451e-006, 3.348307e-006,
  2.001242e-006, 1.928474e-006, 1.840557e-006, 1.747922e-006, 1.661247e-006, 
    1.57929e-006, 1.493609e-006, 1.402215e-006, 1.306103e-006, 1.210983e-006, 
    1.12257e-006, 1.039868e-006, 9.685909e-007, 9.13705e-007, 8.77694e-007, 
    8.6776e-007, 8.816676e-007, 9.20659e-007, 9.772837e-007, 1.040613e-006, 
    1.103447e-006, 1.164045e-006, 1.226133e-006, 1.281764e-006, 
    1.328206e-006, 1.371171e-006, 1.409169e-006, 1.441455e-006, 
    1.463061e-006, 1.470512e-006, 1.457349e-006, 1.426802e-006, 
    1.370674e-006, 1.2989e-006, 1.217937e-006, 1.13002e-006, 1.042352e-006, 
    9.536898e-007, 8.737202e-007, 8.213178e-007, 8.051747e-007, 8.24298e-007, 
    8.635379e-007, 9.122152e-007, 9.594021e-007, 1.003609e-006, 
    1.039123e-006, 1.066442e-006, 1.083578e-006, 1.088545e-006, 
    1.086807e-006, 1.079356e-006, 1.06669e-006, 1.045828e-006, 1.014784e-006, 
    9.780282e-007, 9.31338e-007, 8.843994e-007, 8.46898e-007, 8.220629e-007, 
    8.111354e-007, 8.061684e-007, 8.128741e-007, 8.282721e-007, 
    8.496304e-007, 8.657732e-007, 8.719821e-007, 8.707405e-007, 
    8.697468e-007, 8.72727e-007, 8.821644e-007, 8.935888e-007, 9.005423e-007, 
    9.012874e-007, 8.89615e-007, 8.76204e-007, 8.595644e-007, 8.324939e-007, 
    8.007048e-007, 7.728893e-007, 7.552562e-007, 7.512826e-007, 
    7.656872e-007, 8.086522e-007, 8.848963e-007, 9.864727e-007, 
    1.110152e-006, 1.246001e-006, 1.39849e-006, 1.557932e-006, 1.715884e-006, 
    1.852727e-006, 1.957532e-006, 2.027567e-006, 2.057121e-006, 2.048429e-006,
  -1.688461e-007, -2.080858e-007, -2.286993e-007, -2.334179e-007, 
    -2.177715e-007, -1.820088e-007, -1.305996e-007, -6.230266e-008, 
    1.468675e-008, 9.266932e-008, 1.632018e-007, 2.250415e-007, 
    2.729735e-007, 3.097296e-007, 3.3382e-007, 3.435057e-007, 3.400287e-007, 
    3.30343e-007, 3.19912e-007, 3.07743e-007, 2.990507e-007, 2.913516e-007, 
    2.856393e-007, 2.858876e-007, 3.000439e-007, 3.273624e-007, 
    3.641187e-007, 4.127958e-007, 4.738906e-007, 5.397042e-007, 
    6.089947e-007, 6.807691e-007, 7.470792e-007, 8.081734e-007, 
    8.568504e-007, 8.903783e-007, 9.109917e-007, 9.21671e-007, 9.266375e-007, 
    9.266373e-007, 9.231603e-007, 9.122327e-007, 8.923644e-007, 
    8.623142e-007, 8.193488e-007, 7.714166e-007, 7.185172e-007, 
    6.611481e-007, 6.00302e-007, 5.362258e-007, 4.65694e-007, 3.882078e-007, 
    2.997931e-007, 1.992112e-007, 9.291671e-008, -1.611079e-008, 
    -1.109802e-007, -1.805201e-007, -2.110673e-007, -1.946764e-007, 
    -1.298567e-007, -1.014996e-008, 1.510311e-007, 3.534392e-007, 
    5.742245e-007, 7.81351e-007, 9.519699e-007, 1.066212e-006, 1.123829e-006, 
    1.132026e-006, 1.098498e-006, 1.044605e-006, 9.730795e-007, 
    8.913719e-007, 8.029581e-007, 7.065973e-007, 6.000539e-007, 
    4.940075e-007, 3.976465e-007, 3.134551e-007, 2.488835e-007, 2.02193e-007, 
    1.753708e-007, 1.696587e-007, 1.907688e-007, 2.245447e-007, 2.61301e-007, 
    2.873778e-007, 2.901097e-007, 2.722284e-007, 2.352238e-007, 1.78848e-007, 
    1.07819e-007, 3.05813e-008, -4.615981e-008, -1.149535e-007,
  -1.68543e-008, 5.020115e-008, 1.26694e-007, 1.71646e-007, 1.748742e-007, 
    1.783512e-007, 2.446611e-007, 3.88706e-007, 5.585791e-007, 6.869775e-007, 
    7.262173e-007, 6.685992e-007, 5.695068e-007, 4.835762e-007, 
    4.279452e-007, 4.095673e-007, 4.023651e-007, 4.060904e-007, 
    3.998815e-007, 3.730595e-007, 3.303427e-007, 2.839008e-007, 
    2.513668e-007, 2.550922e-007, 2.82411e-007, 3.281076e-007, 3.829933e-007, 
    4.155278e-007, 4.28442e-007, 4.031102e-007, 3.181735e-007, 1.964806e-007, 
    1.175047e-007, 1.271906e-007, 2.228062e-007, 3.474793e-007, 
    4.244687e-007, 4.502972e-007, 4.470689e-007, 3.874643e-007, 
    2.719803e-007, 1.944945e-007, 2.724769e-007, 5.044376e-007, 
    8.022121e-007, 1.072669e-006, 1.29246e-006, 1.404964e-006, 1.315308e-006, 
    9.365704e-007, 3.122123e-007, -3.558562e-007, -1.039817e-006, 
    -1.663929e-006, -2.083149e-006, -2.267672e-006, -2.141757e-006, 
    -1.756066e-006, -1.329646e-006, -9.57366e-007, -7.537164e-007, 
    -6.504015e-007, -5.341726e-007, -2.617289e-007, 1.27191e-007, 
    4.706617e-007, 6.536984e-007, 7.336671e-007, 7.955068e-007, 
    8.677785e-007, 9.291216e-007, 9.810267e-007, 9.830135e-007, 
    9.668709e-007, 9.584269e-007, 8.83673e-007, 7.068459e-007, 4.207434e-007, 
    1.098056e-007, -1.333315e-007, -2.932702e-007, -4.04284e-007, 
    -4.311059e-007, -3.931086e-007, -3.40458e-007, -2.897937e-007, 
    -1.807666e-007, 1.027729e-009, 1.478038e-007, 1.925073e-007, 
    1.569929e-007, 1.023554e-007, 4.920776e-008, 2.08961e-008, -1.95223e-009, 
    -2.927163e-008,
  3.760397e-007, 5.329985e-007, 5.960801e-007, 6.243927e-007, 5.59573e-007, 
    4.969875e-007, 4.507942e-007, 3.76785e-007, 3.196639e-007, 2.858878e-007, 
    2.126238e-007, 1.470582e-007, 1.373725e-007, 2.501249e-007, 
    4.152794e-007, 5.476516e-007, 6.266276e-007, 6.435152e-007, 
    5.958316e-007, 4.654466e-007, 3.23637e-007, 2.54595e-007, 2.237995e-007, 
    2.382039e-007, 3.435055e-007, 4.689238e-007, 5.272864e-007, 
    5.089084e-007, 4.229786e-007, 3.752946e-007, 3.685891e-007, 
    3.971498e-007, 3.998819e-007, 2.960705e-007, 9.962355e-008, 
    -9.781706e-008, -2.028701e-007, -1.966616e-007, -9.955556e-008, 
    4.473736e-008, 1.388635e-007, 2.468964e-007, 3.295972e-007, 
    3.201599e-007, 2.1908e-007, 1.130329e-007, 3.164332e-007, 1.360014e-006, 
    2.639775e-006, 3.153118e-006, 2.693168e-006, 1.691068e-006, 
    5.081629e-007, -3.66038e-007, -6.141418e-007, -4.579288e-007, 
    7.255312e-008, 8.315174e-007, 1.403722e-006, 1.78246e-006, 1.903656e-006, 
    1.970215e-006, 2.019141e-006, 1.956058e-006, 1.942399e-006, 
    1.919302e-006, 1.939667e-006, 1.930232e-006, 1.670951e-006, 
    1.343125e-006, 9.591727e-007, 6.551886e-007, 6.161972e-007, 8.41701e-007, 
    1.089061e-006, 1.176481e-006, 1.109177e-006, 9.412902e-007, 
    8.205907e-007, 6.857344e-007, 6.586647e-007, 6.67108e-007, 3.549289e-007, 
    3.281593e-008, 1.523858e-009, 1.358826e-007, 3.827454e-007, 
    4.778631e-007, 4.520352e-007, 2.588167e-007, 8.496954e-008, 
    -2.450179e-009, -1.35567e-007, -2.232355e-007, -1.432654e-007, 
    1.214789e-007,
  4.87302e-007, 1.997096e-007, 1.02852e-007, 3.670993e-007, 6.224057e-007, 
    7.72659e-007, 6.243924e-007, 3.894509e-007, 2.685033e-007, 3.385385e-007, 
    4.62715e-007, 4.71159e-007, 4.649503e-007, 4.798512e-007, 6.708347e-007, 
    8.978291e-007, 9.206774e-007, 8.412046e-007, 8.680267e-007, 
    1.058016e-006, 1.286501e-006, 1.110419e-006, 6.566786e-007, 
    3.904445e-007, 4.075805e-007, 5.652844e-007, 5.538604e-007, 
    3.894511e-007, 3.66354e-007, 4.17763e-007, 3.92679e-007, 3.795165e-007, 
    4.068354e-007, 3.117163e-007, 7.379435e-008, -3.299738e-008, 
    9.838141e-008, 2.188881e-008, 9.987184e-008, 2.595623e-007, 
    1.949911e-007, -1.427684e-007, -5.1505e-007, -1.009023e-006, 
    -1.24794e-006, -8.113357e-007, -2.771303e-007, 8.749776e-007, 
    1.473013e-006, 9.055275e-007, 5.421871e-007, -2.537854e-007, 
    -7.105027e-007, -2.960023e-007, 5.732327e-007, 1.467052e-006, 
    1.920294e-006, 1.487912e-006, 1.115135e-006, 1.049571e-006, 
    7.210001e-007, 7.242306e-007, 1.728318e-006, 3.013296e-006, 
    3.392282e-006, 3.901903e-006, 5.59517e-006, 8.071742e-006, 8.907697e-006, 
    7.607569e-006, 6.049407e-006, 5.673649e-006, 5.915297e-006, 
    6.091876e-006, 5.661977e-006, 4.80218e-006, 3.935927e-006, 2.992932e-006, 
    2.156231e-006, 1.707706e-006, 1.850261e-006, 2.308223e-006, 
    2.455992e-006, 2.351188e-006, 1.745952e-006, 6.636319e-007, 
    -7.819926e-008, -3.434416e-007, -2.61236e-007, -4.303629e-007, 
    -3.168652e-007, 3.790201e-007, 9.777978e-007, 1.098993e-006, 
    9.360751e-007, 7.282038e-007,
  1.701746e-006, 1.06795e-006, 1.087571e-006, 1.14494e-006, 6.519604e-007, 
    1.195531e-008, -4.050298e-007, -1.393722e-006, -2.180503e-006, 
    -1.716332e-006, -5.503161e-007, 5.419392e-007, 1.123085e-006, 
    8.990701e-007, 6.395419e-007, 6.320913e-007, 4.835767e-007, 
    3.186703e-007, 3.675959e-007, 7.214985e-007, 1.293951e-006, 
    2.060616e-006, 1.81549e-006, 8.079246e-007, 3.680916e-007, 3.882092e-007, 
    5.431812e-007, 1.185918e-006, 1.417631e-006, 1.114392e-006, 
    1.218452e-006, 1.490895e-006, 1.486424e-006, 1.153384e-006, 
    7.644635e-007, 3.154414e-007, 4.577473e-007, 6.176865e-007, 
    6.720763e-007, 5.939046e-008, -7.822764e-007, -1.109358e-006, 
    -7.812851e-007, -9.297992e-007, -2.164608e-006, -2.23713e-006, 
    -2.843335e-007, 1.937478e-007, -1.693443e-007, 3.869645e-007, 
    4.008743e-007, 9.51969e-007, 1.800839e-006, 5.431793e-007, 2.829074e-007, 
    1.03343e-006, 2.737625e-006, 4.441571e-006, 5.511226e-006, 4.767657e-006, 
    2.94922e-006, 1.677652e-006, 1.015049e-006, 8.481566e-007, 1.914084e-006, 
    3.090532e-006, 4.624605e-006, 5.243504e-006, 4.69787e-006, 3.92922e-006, 
    3.024225e-006, 2.620402e-006, 3.152868e-006, 3.663484e-006, 
    3.712908e-006, 3.565882e-006, 2.0405e-006, 1.136994e-006, 1.566394e-006, 
    1.280043e-006, 1.118614e-006, 1.850508e-006, 2.766681e-006, 
    3.173732e-006, 2.684227e-006, 1.324002e-006, 5.096517e-007, 
    9.470004e-007, 1.539323e-006, 1.229379e-006, 9.872365e-007, 
    1.298421e-006, 2.537699e-006, 4.525264e-006, 4.469883e-006, 2.781087e-006,
  3.767293e-006, 3.551476e-006, 3.658516e-006, 4.616412e-006, 4.361603e-006, 
    2.117982e-006, 1.006156e-007, -1.844978e-006, -1.272774e-006, 
    -8.734232e-007, -1.894596e-007, 7.003873e-007, 3.392528e-006, 
    5.899401e-006, 7.031397e-006, 5.84104e-006, 3.6985e-006, 2.211614e-006, 
    2.335542e-006, 2.591841e-006, 3.461573e-006, 4.476094e-006, 
    6.326317e-006, 5.638879e-006, 2.270222e-006, -4.574331e-007, 
    -8.816187e-007, -4.7308e-007, 9.099958e-007, 3.018513e-006, 
    4.431886e-006, 4.524025e-006, 3.834598e-006, 2.330823e-006, 
    1.535847e-006, 1.561179e-006, 1.093529e-006, 1.527696e-007, 
    -3.655423e-007, 1.639473e-007, 1.892235e-006, 3.797591e-006, 
    3.512981e-006, 1.407449e-006, 1.368735e-007, -5.379006e-007, 
    -2.061042e-007, 1.640896e-006, 2.845909e-006, 3.67292e-006, 
    3.914814e-006, 3.06818e-006, 2.871486e-006, 2.821322e-006, 2.636049e-006, 
    1.637669e-006, 3.70744e-006, 5.450627e-006, 4.725192e-006, 2.336535e-006, 
    8.516345e-007, 1.356784e-006, 2.810392e-006, 3.260159e-006, 3.85372e-006, 
    3.69552e-006, 2.409301e-006, 1.395525e-006, 1.297924e-006, 2.316419e-006, 
    3.921026e-006, 4.215321e-006, 2.789283e-006, 2.764446e-006, 
    2.837711e-006, 2.615436e-006, 1.621031e-006, 1.204045e-006, 
    9.072646e-007, 6.939281e-007, -3.277928e-007, 8.198731e-008, 
    2.043479e-006, 2.455992e-006, 2.740604e-006, 3.445181e-006, 
    4.127901e-006, 5.228103e-006, 5.292674e-006, 4.920893e-006, 
    3.670684e-006, 3.67441e-006, 4.614427e-006, 5.302114e-006, 4.728421e-006, 
    3.824913e-006,
  7.092238e-006, 6.265967e-006, 4.333288e-006, 5.97341e-006, 6.612672e-006, 
    6.387168e-006, 6.314152e-006, 7.235538e-006, 7.179164e-006, 
    6.198665e-006, 5.135467e-006, 4.54389e-006, 6.34718e-006, 7.123786e-006, 
    8.378463e-006, 1.037423e-005, 9.873294e-006, 6.85432e-006, 5.890464e-006, 
    6.484024e-006, 7.509223e-006, 7.984321e-006, 8.405281e-006, 
    7.924968e-006, 7.274528e-006, 7.310789e-006, 5.625219e-006, 
    2.975048e-006, 2.051922e-006, 5.106906e-006, 6.027301e-006, 
    6.405295e-006, 6.730637e-006, 6.065799e-006, 6.030285e-006, 
    5.670916e-006, 7.607576e-006, 7.280243e-006, 7.481911e-006, 
    8.651401e-006, 9.59514e-006, 7.665192e-006, 6.954902e-006, 7.573051e-006, 
    6.502152e-006, 4.921139e-006, 4.117717e-006, 4.745803e-006, 
    5.023461e-006, 5.855441e-006, 4.108286e-006, 3.091778e-006, 
    5.004586e-006, 6.127637e-006, 6.935777e-006, 4.732394e-006, 
    4.656644e-006, 5.789629e-006, 4.83198e-006, 4.064574e-006, 5.11287e-006, 
    4.518062e-006, 3.616544e-006, 4.614672e-006, 5.976639e-006, 
    6.382945e-006, 6.496939e-006, 6.445034e-006, 4.591826e-006, 
    3.887249e-006, 3.527632e-006, 3.545265e-006, 2.805671e-006, 2.95543e-006, 
    3.405197e-006, 2.215587e-006, 9.41287e-007, -7.497474e-007, 
    -1.269547e-006, 1.708977e-007, 1.335671e-006, 2.563529e-006, 
    4.009189e-006, 4.97379e-006, 5.735985e-006, 4.840425e-006, 4.721713e-006, 
    5.829615e-006, 5.424552e-006, 4.995647e-006, 5.017502e-006, 
    5.968444e-006, 5.424055e-006, 5.327449e-006, 5.960252e-006, 6.136826e-006,
  4.464171e-006, 5.905113e-006, 6.976257e-006, 5.32372e-006, 4.148018e-006, 
    3.894698e-006, 5.513461e-006, 5.999485e-006, 6.233433e-006, 
    6.015876e-006, 3.579042e-006, 3.600648e-006, 5.754115e-006, 
    8.741306e-006, 8.493698e-006, 9.167727e-006, 1.021999e-005, 
    9.426258e-006, 7.833329e-006, 7.862385e-006, 8.678719e-006, 
    6.689164e-006, 5.001109e-006, 6.039472e-006, 6.546361e-006, 
    8.254285e-006, 8.925084e-006, 6.351403e-006, 6.858043e-006, 6.98694e-006, 
    7.059954e-006, 7.976128e-006, 7.333643e-006, 8.659841e-006, 
    9.991012e-006, 9.122527e-006, 7.172956e-006, 4.866999e-006, 
    5.756598e-006, 6.801671e-006, 5.778209e-006, 6.778322e-006, 8.30271e-006, 
    7.093733e-006, 7.088018e-006, 7.194065e-006, 5.701218e-006, 
    6.413244e-006, 6.676995e-006, 7.826618e-006, 5.94535e-006, 6.344699e-006, 
    7.810229e-006, 8.709017e-006, 7.792847e-006, 6.392878e-006, 
    5.500295e-006, 6.959619e-006, 8.023066e-006, 6.886106e-006, 
    6.485512e-006, 5.853955e-006, 4.932315e-006, 6.465147e-006, 
    6.252065e-006, 4.847878e-006, 6.872942e-006, 6.527982e-006, 
    5.802294e-006, 5.123797e-006, 3.038871e-006, 4.303734e-006, 
    4.579406e-006, 5.131991e-006, 4.382213e-006, 2.471141e-006, 
    1.522494e-009, 4.142839e-007, 2.622135e-006, 2.833738e-006, 
    3.124307e-006, 2.457482e-006, 3.349316e-006, 4.365824e-006, 
    3.990066e-006, 5.320493e-006, 7.352515e-006, 7.370396e-006, 
    5.280755e-006, 4.862528e-006, 5.621991e-006, 5.878042e-006, 
    4.696876e-006, 4.328322e-006, 4.121692e-006, 4.16888e-006,
  5.910331e-006, 4.76443e-006, 5.173219e-006, 6.143036e-006, 5.831849e-006, 
    4.592323e-006, 3.521176e-006, 4.787775e-006, 4.133368e-006, 
    3.364219e-006, 4.178819e-006, 6.250326e-006, 8.66779e-006, 7.92695e-006, 
    5.132242e-006, 4.565749e-006, 4.198686e-006, 5.985825e-006, 
    6.698358e-006, 4.546378e-006, 5.116592e-006, 4.872965e-006, 
    5.404439e-006, 8.958114e-006, 1.141855e-005, 1.037671e-005, 
    7.716597e-006, 8.051633e-006, 8.541632e-006, 6.210097e-006, 
    5.814471e-006, 6.450751e-006, 6.854325e-006, 6.212083e-006, 
    5.672162e-006, 5.677128e-006, 5.525388e-006, 5.117337e-006, 
    3.293188e-006, 5.198059e-006, 5.612559e-006, 5.556929e-006, 
    7.837547e-006, 6.504142e-006, 6.707298e-006, 7.010038e-006, 
    8.367035e-006, 1.002156e-005, 9.703921e-006, 8.214052e-006, 
    7.032639e-006, 7.72678e-006, 7.471974e-006, 7.682573e-006, 6.432612e-006, 
    5.47249e-006, 6.818058e-006, 8.271918e-006, 6.979988e-006, 4.636031e-006, 
    6.612676e-006, 8.217528e-006, 9.821886e-006, 1.030071e-005, 
    9.244468e-006, 7.629182e-006, 6.904986e-006, 6.671535e-006, 
    6.905728e-006, 7.419074e-006, 9.52138e-006, 1.105694e-005, 7.012271e-006, 
    4.714266e-006, 2.975303e-006, 1.584271e-006, 2.835477e-006, 
    5.215687e-006, 4.815593e-006, 3.706205e-006, 3.137011e-007, 
    -4.877347e-007, 9.842533e-007, 3.804797e-006, 4.911459e-006, 
    3.527883e-006, 2.87745e-006, 3.209496e-006, 3.573086e-006, 5.744183e-006, 
    7.821158e-006, 7.432734e-006, 5.986576e-006, 4.162177e-006, 
    3.902394e-006, 5.941374e-006,
  6.44429e-006, 6.932052e-006, 6.227478e-006, 5.243503e-006, 4.553582e-006, 
    3.168268e-006, 2.283141e-006, 2.288107e-006, 6.243936e-007, 
    1.428063e-006, 1.581546e-006, 2.743091e-006, 2.139837e-006, 
    2.663863e-006, 4.802179e-006, 4.983227e-006, 7.039594e-006, 
    8.683935e-006, 7.873063e-006, 4.913447e-006, 7.472718e-006, 
    9.766507e-006, 1.016933e-005, 8.450483e-006, 6.480797e-006, 
    6.601997e-006, 7.757579e-006, 8.785759e-006, 5.92498e-006, 2.478839e-006, 
    5.257971e-007, 7.612362e-007, 2.888872e-006, 2.103829e-006, 
    4.344001e-007, 3.058449e-008, 2.958259e-007, -1.39869e-006, 
    -2.374716e-006, -7.33351e-007, 2.311201e-006, 4.369795e-006, 
    5.659251e-006, 7.787628e-006, 7.697232e-006, 7.358227e-006, 
    9.505236e-006, 6.078717e-006, 3.947847e-006, 2.84144e-006, 3.07216e-006, 
    4.28388e-006, 2.395402e-006, 1.517714e-006, 3.526642e-006, 3.122321e-006, 
    2.097371e-006, 3.035897e-006, 3.49585e-006, 3.417616e-006, 4.966092e-006, 
    6.057853e-006, 8.627809e-006, 7.513947e-006, 4.134614e-006, 
    4.366822e-006, 6.667804e-006, 9.444888e-006, 9.700194e-006, 
    7.040584e-006, 4.9343e-006, 2.618664e-006, 4.860631e-007, 8.387178e-007, 
    2.496225e-006, 1.718894e-006, -1.606459e-007, 2.264758e-006, 
    1.613831e-006, -1.023431e-006, 7.152867e-007, 2.600285e-006, 
    3.505529e-006, 4.523281e-008, -5.816109e-007, 1.141463e-006, 
    2.854849e-006, 3.975416e-006, 3.516707e-006, 3.511246e-006, 
    5.361224e-006, 7.920251e-006, 7.446639e-006, 7.244482e-006, 
    9.250674e-006, 7.33836e-006,
  8.081435e-006, 4.593072e-006, 3.056015e-006, 1.036162e-006, 1.102719e-006, 
    -9.091855e-007, -2.009139e-006, -1.685534e-006, 2.039342e-007, 
    4.083267e-007, -2.877277e-008, 2.133711e-007, -3.819332e-007, 
    2.071542e-006, 2.01293e-006, 1.962268e-006, 3.190373e-006, 3.046574e-006, 
    3.59767e-006, 6.769384e-006, 8.899009e-006, 9.051993e-006, 6.425664e-006, 
    2.702112e-006, 1.582543e-006, 3.261899e-006, 1.458604e-006, 
    -3.484056e-007, -1.429482e-006, -1.340075e-006, -1.948043e-006, 
    -1.740918e-006, -4.461872e-006, -5.939572e-006, -6.38462e-006, 
    -5.407601e-006, -5.917718e-006, -4.680911e-006, -3.959449e-006, 
    -1.897872e-006, 1.321514e-006, 3.820445e-006, 3.403213e-006, 
    3.310328e-006, 7.582603e-007, 1.540575e-006, 1.862431e-006, 
    4.371359e-007, -2.227316e-007, 1.419117e-006, 2.111337e-007, 
    -2.101766e-006, -1.87055e-006, -1.723274e-006, -1.777171e-006, 
    -2.577472e-007, 6.010559e-007, 1.336673e-006, -4.191716e-007, 
    1.242552e-006, 4.517329e-006, 3.987592e-006, 3.627723e-006, 8.89886e-007, 
    7.125673e-007, 9.835167e-007, -1.837434e-007, -5.434413e-008, 
    7.152958e-007, -1.646222e-007, 8.695242e-007, -6.839218e-007, 
    -1.754324e-006, -8.70441e-007, -1.219621e-006, -7.775488e-007, 
    3.775385e-007, -7.462622e-007, -1.336604e-006, -2.587805e-006, 
    -1.059441e-006, 3.705718e-007, -1.822882e-006, -3.171117e-007, 
    -1.049753e-006, 7.113158e-007, 4.205638e-006, 5.406178e-006, 
    1.600674e-006, 7.624876e-007, 1.783959e-006, 3.08036e-006, 3.893223e-006, 
    4.995411e-006, 7.234299e-006, 9.336116e-006,
  -1.959474e-006, -3.141628e-006, -4.49242e-006, -4.545071e-006, 
    -5.382766e-006, -7.472407e-006, -9.379011e-006, -8.522939e-006, 
    -6.032209e-006, -6.051579e-006, -3.123751e-006, -7.604212e-007, 
    -1.362925e-006, -6.536357e-007, 2.395893e-006, 3.807279e-006, 
    4.806894e-006, 2.898807e-006, 2.63704e-006, 3.658017e-006, 1.421351e-006, 
    1.311335e-006, -1.069369e-006, -2.181496e-006, -4.48621e-006, 
    -5.727976e-006, -6.867171e-006, -8.71864e-006, -9.956928e-006, 
    -9.801706e-006, -9.802201e-006, -1.082715e-005, -1.030387e-005, 
    -9.765196e-006, -7.44906e-006, -7.761988e-006, -8.721367e-006, 
    -6.135519e-006, -6.014821e-006, -4.834405e-006, -3.061661e-006, 
    -3.286914e-006, -2.85701e-006, -2.13207e-006, -1.447119e-006, 
    -3.042282e-006, -4.057052e-006, -2.79344e-006, -1.782639e-006, 
    -4.355323e-006, -3.839003e-006, -4.517249e-006, -6.314582e-006, 
    -4.466834e-006, -1.607794e-006, 1.15524e-007, 1.623775e-006, 
    -8.128118e-007, -1.834538e-006, -2.048127e-006, -2.812059e-006, 
    -3.47168e-006, -6.880076e-006, -1.152998e-005, -6.757389e-006, 
    -6.215978e-006, -6.238581e-006, -4.492413e-006, -3.458023e-006, 
    -3.681787e-006, -1.540993e-006, -3.529552e-006, -4.066493e-006, 
    -4.698799e-006, -5.588896e-006, -8.629228e-006, -1.019136e-005, 
    -9.24911e-006, -4.76809e-006, -3.506956e-006, -1.940103e-006, 
    -2.657094e-006, -5.153015e-007, 1.502816e-006, 2.580418e-006, 
    5.644844e-006, 4.554335e-006, -5.863185e-007, -1.62841e-006, 
    -6.215851e-007, 2.227018e-006, 2.059631e-006, 2.84542e-006, 
    2.699879e-006, 5.787006e-007, 4.731519e-007,
  -8.443712e-006, -6.919821e-006, -6.231387e-006, -6.023516e-006, 
    -6.315577e-006, -4.600206e-006, -2.206085e-006, -1.058943e-006, 
    -1.534043e-006, 1.742475e-006, 1.421353e-006, -1.894652e-006, 
    -2.756433e-006, -8.741717e-007, 1.465312e-006, 1.602402e-006, 
    6.800219e-007, 5.916081e-007, 1.928242e-006, 9.052783e-007, 
    -1.339584e-006, -6.625278e-006, -1.056887e-005, -1.235229e-005, 
    -1.360821e-005, -1.178952e-005, -8.649102e-006, -8.479477e-006, 
    -9.616931e-006, -8.487918e-006, -9.10706e-006, -7.565784e-006, 
    -5.9207e-006, -5.320924e-006, -4.383888e-006, -1.96419e-006, 
    -1.24695e-006, -1.258126e-006, -3.413079e-006, -7.040508e-007, 
    -1.028398e-006, -3.821879e-007, 4.694175e-007, -1.98182e-006, 
    -7.767196e-006, -1.16631e-005, -7.87498e-006, -4.691849e-006, 
    -2.749977e-006, -3.102385e-006, -4.464597e-006, -4.220714e-006, 
    -5.31297e-006, -2.126853e-006, 2.747183e-007, 1.680393e-006, 
    6.325972e-007, -3.501485e-006, 1.158845e-006, 2.351942e-006, 
    1.023502e-006, 2.235574e-007, -8.949108e-006, -8.480456e-006, 
    -6.765586e-006, -4.931255e-006, -5.437643e-006, -6.632221e-006, 
    -8.666968e-006, -4.032961e-006, -4.465102e-006, -5.353957e-006, 
    -7.45055e-006, -8.513996e-006, -8.58155e-006, -1.043649e-005, 
    -1.415111e-005, -1.299204e-005, -3.754313e-006, 9.263886e-007, 
    2.378754e-006, 5.457579e-006, 4.59729e-006, 2.022371e-006, 1.653072e-006, 
    1.784447e-006, 3.10022e-006, 5.859001e-007, 1.220938e-006, 4.163667e-006, 
    7.691888e-007, -2.070919e-007, -7.293784e-007, -4.059792e-006, 
    -6.348855e-006, -8.321769e-006,
  -6.290991e-006, -5.581444e-006, -5.304531e-006, -4.33074e-006, 
    -2.832429e-006, -1.283206e-006, 6.318414e-007, 1.757624e-006, 
    6.40331e-006, 7.318238e-006, 7.237286e-007, -1.689265e-006, 
    -1.05994e-006, -3.66019e-006, -2.753206e-006, 1.67343e-006, 
    1.342378e-006, 4.65292e-006, 2.814364e-006, -2.416182e-007, 
    -5.070835e-006, -5.996691e-006, -7.430186e-006, -6.533379e-006, 
    -5.974834e-006, -5.999424e-006, -5.282182e-006, -7.399884e-006, 
    -7.556347e-006, -5.512405e-006, -2.171066e-006, -1.77842e-006, 
    -2.237321e-007, 2.492003e-006, 4.520547e-006, 3.608597e-006, 
    2.364597e-006, 3.99381e-007, -1.63239e-006, -9.451978e-007, 
    1.176977e-006, 1.023242e-006, 3.004106e-006, 2.231729e-006, 
    -5.018919e-007, 2.155732e-006, 1.08707e-006, 2.125431e-006, 
    4.977019e-006, 9.167015e-007, 2.20615e-006, 5.140191e-006, 7.205243e-006, 
    8.262974e-006, 8.996612e-006, 3.839326e-006, -1.442495e-007, 
    2.925884e-006, 5.447899e-006, 5.069913e-006, 3.633682e-006, 
    -1.64282e-006, -5.544931e-006, -4.395813e-006, 4.209905e-007, 
    -1.240238e-006, -3.812183e-006, -6.858721e-006, -6.005637e-006, 
    -5.920201e-006, -7.477869e-006, -1.078518e-005, -1.024948e-005, 
    -8.081611e-006, -5.183336e-006, -3.710604e-006, -6.130306e-006, 
    -6.266402e-006, -2.056326e-006, 4.235439e-006, 6.112488e-006, 
    7.012271e-006, 9.005056e-006, 7.800048e-006, 8.505864e-006, 
    3.923013e-006, 8.595816e-007, 1.226397e-006, 5.522406e-006, 
    4.871717e-006, 2.048691e-006, -1.520382e-006, -3.449091e-006, 
    -5.990238e-006, -6.086597e-006, -6.487193e-006,
  -4.444488e-006, -4.841354e-006, -3.387002e-006, -1.701432e-006, 
    -4.611579e-007, 5.071702e-007, 1.730555e-006, 8.638026e-007, 
    9.827618e-007, -4.06178e-006, -9.304003e-006, -7.234479e-006, 
    -4.875131e-006, -2.812067e-006, 2.0929e-006, 9.328656e-006, 
    1.334203e-005, 1.020012e-005, 6.199907e-006, -2.185207e-007, 
    -5.134163e-006, -3.309517e-006, -4.984902e-006, -5.437648e-006, 
    -5.513396e-006, -4.676201e-006, -1.818405e-006, -2.233403e-006, 
    -2.854285e-006, 1.040135e-006, 1.443956e-006, 2.997402e-006, 
    9.680074e-006, 1.017901e-005, 8.63103e-006, 4.304481e-006, 3.434255e-006, 
    2.419486e-006, 7.540311e-007, 3.352297e-006, 8.871935e-006, 
    1.405978e-005, 1.234862e-005, 3.494606e-006, -3.086747e-006, 
    2.734141e-006, 6.941755e-007, 7.602466e-008, 5.719598e-006, 
    6.805392e-006, 9.542237e-006, 1.04306e-005, 8.352392e-006, 8.884115e-006, 
    1.287886e-005, 9.880005e-006, 5.549478e-006, 4.851852e-006, 
    2.892593e-006, 1.435263e-006, 2.064153e-007, 3.245503e-006, 
    4.696874e-006, 5.529608e-006, 2.937799e-006, 1.441225e-006, 
    -2.063498e-007, -2.64815e-006, -6.187427e-006, -4.577605e-006, 
    -6.177494e-006, -5.656696e-006, -3.414568e-006, -2.06825e-006, 
    -1.198518e-006, -2.016093e-006, -1.962449e-006, -8.475939e-007, 
    -2.329211e-007, 5.609327e-006, 6.39909e-006, 7.334384e-006, 
    6.113734e-006, 5.883012e-006, 5.130503e-006, 1.584025e-006, 
    -8.259867e-007, 1.343369e-006, 1.298666e-006, -2.508059e-007, 
    -2.056577e-006, -1.86535e-006, -3.544459e-006, -4.207312e-006, 
    -2.355344e-006, -3.843224e-006,
  -2.272396e-006, -1.382547e-006, -1.320459e-006, -8.786378e-007, 
    -1.681009e-007, -4.119192e-008, 2.972564e-006, 6.20912e-007, 
    -2.783258e-006, -6.780492e-006, -2.627046e-006, 4.341546e-007, 
    1.172257e-006, 6.741073e-006, 1.209978e-005, 1.376697e-005, 
    1.267422e-005, 5.180671e-006, -1.666913e-006, -3.098419e-006, 
    -5.885431e-006, -9.420733e-006, -4.908907e-006, -2.796914e-006, 
    -2.356319e-008, 2.280904e-006, 3.336652e-006, 2.933823e-006, 
    -1.58665e-007, 2.871293e-007, 9.278765e-007, 4.75996e-006, 8.062058e-006, 
    7.764279e-006, 2.244147e-006, 1.664494e-006, 3.921772e-006, 
    2.185287e-006, 1.077139e-006, 2.622885e-006, 1.149702e-005, 
    1.071422e-005, -1.653698e-007, -3.637593e-006, -3.467967e-006, 
    -8.76902e-007, 4.515332e-007, 2.725954e-006, 6.943725e-006, 
    1.469382e-005, 1.499731e-005, 6.460192e-006, 6.728409e-006, 
    1.064518e-005, 1.16972e-005, -1.685949e-007, -1.117223e-007, 
    7.845811e-007, -5.205147e-007, 3.388057e-006, 8.099061e-006, 
    3.060482e-006, 4.051912e-006, 1.809531e-006, 6.102382e-007, 
    -2.138284e-006, -8.555226e-006, -8.768558e-006, -5.954967e-006, 
    -3.987767e-006, -3.78486e-006, -4.06023e-007, 5.570882e-007, 
    -5.845886e-007, -1.111592e-006, -6.218409e-007, -2.530373e-007, 
    -1.402855e-007, -1.921721e-006, 1.999775e-006, 6.473347e-006, 
    6.546867e-006, 3.584264e-006, 6.486509e-006, 9.491836e-006, 
    5.582508e-006, -1.817414e-006, 1.956556e-006, 1.156612e-006, 
    -2.7316e-006, -3.574263e-006, -3.335843e-006, -2.75867e-006, 
    -3.552403e-006, -4.521724e-006, -3.455547e-006,
  -2.517963e-007, 1.47058e-007, 7.520453e-007, 3.370487e-007, -4.015524e-007, 
    9.487394e-007, 1.802076e-006, 1.154138e-006, -7.58926e-007, 
    -2.063782e-006, -1.440168e-006, 4.200172e-006, 6.335511e-006, 
    8.182516e-006, 1.94833e-005, 2.209001e-005, 1.320172e-005, 1.025477e-005, 
    -2.653618e-006, -4.64665e-006, -8.740988e-006, -8.452655e-006, 
    -3.447354e-006, 1.151144e-006, 9.743198e-007, -1.41632e-006, 
    2.536017e-007, -1.685536e-006, -2.300952e-006, -7.397648e-008, 
    -1.186818e-007, 3.819943e-006, 9.280722e-006, 9.059688e-006, 
    1.023887e-005, 4.425182e-006, 1.158103e-006, 3.189626e-006, 
    1.100733e-006, 3.696019e-006, -3.379799e-006, -1.152104e-005, 
    -7.666618e-006, -6.328988e-006, -5.453796e-006, 7.342831e-006, 
    4.343226e-006, 8.369769e-006, 1.754193e-005, 2.334196e-005, 
    1.490343e-005, 6.197184e-006, 5.145164e-006, 1.262231e-005, 
    5.949576e-006, -5.041267e-006, -3.176392e-006, 2.122459e-006, 
    6.319868e-006, 9.101917e-006, 3.392041e-006, -4.448706e-006, 
    -3.284182e-006, -5.829541e-006, -7.151775e-006, -9.001018e-006, 
    -1.091879e-005, -8.174e-006, -4.173531e-006, -3.083761e-006, 
    6.181835e-007, 2.794295e-007, -3.538694e-007, -4.740732e-007, 
    -1.974067e-007, 4.085741e-007, -3.690185e-007, -2.698044e-009, 
    -3.467716e-006, -5.173206e-009, 3.139539e-007, -5.086986e-008, 
    -4.271315e-007, -3.119523e-006, 9.498046e-006, 6.009181e-006, 
    -5.284401e-006, -2.926754e-008, -3.587669e-006, -5.573998e-006, 
    -3.695211e-006, -4.422138e-006, -3.183599e-006, -9.807118e-007, 
    -1.378822e-006, -1.561239e-008,
  6.67108e-007, 1.40104e-007, -3.739847e-007, -4.700979e-007, -1.773455e-006, 
    -5.788326e-006, -2.651381e-006, 3.459882e-007, 1.727078e-006, 
    3.124596e-007, 6.551083e-006, 1.2594e-005, 1.453463e-005, 9.713862e-006, 
    1.785287e-005, 1.076663e-005, -3.435664e-006, 4.592828e-006, 
    2.347471e-006, -2.485649e-007, -6.891754e-006, -5.443613e-006, 
    -4.060041e-006, -1.34579e-006, -1.668399e-006, -5.579709e-006, 
    -1.699195e-006, -3.432448e-006, -2.681929e-006, -6.086346e-006, 
    7.38927e-006, 1.272587e-005, 6.792229e-006, 4.77337e-006, 8.158666e-006, 
    7.481905e-006, 4.994155e-006, 3.718865e-006, 2.523593e-007, 
    5.799066e-006, 4.311696e-007, -7.706843e-006, -1.364023e-005, 
    -3.774676e-006, -1.955494e-006, 1.237396e-005, 1.307183e-005, 
    1.481626e-005, 3.141492e-005, 2.947653e-005, 2.216898e-005, 
    6.727903e-006, 6.215807e-006, 8.936266e-006, 6.698356e-006, 
    -1.437918e-006, -1.46847e-006, 9.026913e-006, 5.841543e-006, 
    -3.331115e-006, -6.953091e-006, -7.793766e-006, -6.347851e-006, 
    -5.827813e-006, -1.286638e-005, -1.117211e-005, -7.598814e-006, 
    -3.278222e-006, -7.641474e-007, -4.316043e-007, 9.688556e-007, 
    -3.697642e-007, 4.103113e-007, -4.765207e-008, -5.371526e-007, 
    -3.0097e-007, -1.919426e-007, -1.561801e-007, -4.507319e-006, 
    3.686833e-006, 2.416506e-006, 4.381363e-007, -4.091824e-006, 
    -4.858233e-006, 8.226474e-006, 8.229945e-006, -9.009818e-007, 
    -7.653187e-006, -1.155109e-005, -1.075712e-005, -7.227529e-006, 
    -6.455398e-006, -3.967649e-006, -2.738998e-007, -2.083016e-008, 
    8.305251e-007,
  -1.800227e-007, -4.340864e-007, 8.625625e-007, 9.343369e-007, 
    -5.659422e-008, -8.50825e-007, -1.068878e-006, 1.963261e-006, 
    2.132141e-006, 4.319172e-007, 5.405927e-006, 1.645413e-005, 
    1.372922e-005, 1.432477e-005, 1.763407e-005, 1.334303e-005, 
    -5.470181e-006, -4.791178e-006, 9.328542e-007, -2.408735e-006, 
    -9.979029e-006, -3.119283e-006, -2.262186e-007, -4.726618e-006, 
    -5.637823e-006, -3.414571e-006, -6.446917e-007, -9.866762e-007, 
    1.662505e-006, 7.826624e-006, 1.702511e-005, 1.629471e-005, 
    1.303159e-005, 8.164626e-006, 6.872447e-006, 9.547701e-006, 
    7.643831e-006, 3.646595e-006, 4.002732e-006, 1.02796e-005, 1.038143e-005, 
    1.152633e-005, -5.8757e-007, -1.92345e-006, -9.220304e-006, 
    1.161077e-005, 2.452411e-005, 2.394322e-005, 3.907411e-005, 
    3.446716e-005, 1.532662e-005, 3.373898e-006, 1.650828e-005, 
    1.137011e-005, 4.364585e-006, 3.085566e-006, 7.006318e-006, 
    1.078028e-005, 3.051056e-006, -5.874987e-006, -7.04746e-006, 
    -9.25532e-006, -1.078344e-005, -1.032275e-005, -1.025072e-005, 
    -4.358308e-006, -7.927083e-007, -3.349942e-007, 1.306368e-006, 
    1.582348e-007, -1.412782e-007, 1.021635e-008, -9.593523e-007, 
    -2.748934e-007, -1.09396e-006, 2.968145e-007, -3.017145e-007, 
    -4.360735e-007, -4.715439e-006, 1.109717e-005, 1.023242e-005, 
    3.078378e-006, -4.077177e-006, -4.512149e-007, 1.796121e-006, 
    -3.064139e-006, -4.781741e-006, -1.146888e-005, -1.242107e-005, 
    -7.315697e-006, -5.467702e-006, -2.910413e-006, -1.343057e-006, 
    6.360651e-007, 1.458156e-007, -1.283652e-007,
  -1.971594e-007, 3.882083e-007, 8.96338e-007, 3.919287e-006, -2.875142e-006, 
    -2.00318e-006, -2.212293e-006, 3.785672e-006, 2.985231e-006, 
    -5.316942e-007, 3.003115e-006, 7.966177e-006, 8.39014e-006, 
    1.415316e-005, 1.910009e-005, 2.267811e-005, 7.834067e-006, 
    -2.815941e-007, -1.752342e-006, 1.250807e-005, -2.371482e-006, 
    3.549252e-006, 8.429488e-007, -5.977065e-006, -2.148467e-006, 
    8.140541e-006, 9.027655e-006, 5.406429e-006, 4.09612e-006, 8.656622e-006, 
    1.002155e-005, 1.418917e-005, 1.465806e-005, 8.926079e-006, 
    1.391151e-005, 1.58874e-005, 1.402402e-005, -8.823627e-007, 
    1.819137e-005, 1.271445e-005, 1.286618e-005, 4.246125e-006, 
    4.182795e-006, -3.484347e-006, -2.130913e-005, 9.991636e-007, 
    1.807142e-005, 1.359064e-005, 1.486592e-005, 3.13265e-005, 1.112501e-005, 
    -4.345638e-006, 1.248324e-005, 1.058706e-005, 4.364083e-006, 
    3.367197e-006, 3.258167e-006, 1.833621e-006, -3.901092e-006, 
    -5.280934e-006, -9.784053e-006, -1.017571e-005, -1.035677e-005, 
    -6.380398e-006, -2.463623e-006, -8.475936e-007, -3.190989e-007, 
    -2.2125e-007, -5.383954e-007, -1.767494e-006, -4.852482e-007, 
    -1.328653e-006, -1.226581e-006, -1.181132e-006, -1.334118e-006, 
    -2.922773e-007, -5.366567e-007, -1.578001e-006, -1.094487e-005, 
    5.614052e-006, 6.886112e-006, 5.513706e-006, 3.24635e-007, 4.695394e-006, 
    -4.298203e-006, -6.664013e-006, -9.28688e-006, -1.119098e-005, 
    -4.243317e-006, 1.298913e-006, 1.694541e-006, -1.106378e-006, 
    -1.669642e-006, -3.536197e-007, -6.151377e-007, 1.122889e-007,
  -7.254066e-007, -5.982483e-007, -1.83008e-006, -1.056513e-005, 
    -9.978539e-006, -5.038786e-006, 4.460453e-006, 1.049394e-005, 
    4.616415e-006, 9.072119e-006, 9.186104e-006, 9.096686e-006, 
    1.068888e-005, -9.71726e-006, 4.048685e-006, 6.12541e-006, 1.45684e-005, 
    8.057585e-006, 9.274772e-006, 1.920167e-005, 1.175682e-005, 
    2.251296e-005, 1.318632e-005, 1.667642e-005, 8.442043e-006, 
    9.928928e-006, 1.333955e-005, 7.641094e-006, 7.698218e-006, 
    7.709656e-006, 1.15539e-005, 1.019939e-005, 1.124222e-005, 4.452238e-006, 
    4.324596e-006, 2.216651e-005, 3.458191e-005, 3.634173e-006, 
    1.802026e-005, 4.053616e-005, 2.522895e-005, 1.644174e-005, 
    8.032752e-006, -1.000015e-005, -7.198469e-006, 8.714225e-006, 
    7.395225e-006, 2.129906e-006, 2.147236e-005, 1.502884e-005, 
    -1.191792e-005, -5.586422e-006, 8.84982e-006, 8.091854e-006, 
    1.582407e-005, 5.85719e-006, 5.965216e-006, 3.480432e-006, 3.891204e-006, 
    -1.212175e-006, -4.996815e-006, -7.74211e-006, -6.355314e-006, 
    -4.90841e-006, -1.855409e-006, -1.323935e-006, -1.154805e-006, 
    -1.703914e-006, -2.532668e-006, -2.787725e-006, -2.298472e-006, 
    -2.453693e-006, -2.330509e-006, -1.057452e-006, 7.180756e-008, 
    1.837594e-006, 1.00911e-005, -4.830945e-006, -3.993737e-006, 
    1.252738e-006, 8.335999e-006, 3.166933e-007, -2.540255e-007, 
    -2.351117e-006, -9.328331e-006, 4.203157e-006, 8.412979e-006, 
    6.635266e-006, 2.112774e-006, 6.433122e-006, 5.890706e-006, 
    3.702475e-006, -1.041558e-006, 8.789539e-007, 5.866432e-007, 
    -2.205043e-007,
  2.909484e-006, 1.993061e-006, 1.69166e-007, -6.824444e-006, -5.573733e-006, 
    -4.963782e-006, -2.498164e-006, 1.201857e-005, 2.413495e-005, 
    4.488804e-005, 3.224068e-005, 2.344924e-005, 1.233621e-005, 
    -2.503628e-006, 7.079812e-006, 9.034113e-006, 1.250037e-005, 
    1.420431e-005, 1.599444e-005, 2.164745e-005, 2.357566e-005, 
    1.520469e-005, 9.50673e-006, 5.143418e-006, 2.393419e-006, 
    -7.701019e-007, -4.92033e-006, -8.9901e-007, 1.131995e-005, 
    1.754492e-005, 1.171085e-005, 7.995986e-006, 9.581236e-006, 
    4.750509e-006, 2.644003e-006, 1.574212e-005, 2.35019e-005, 1.688927e-005, 
    2.900886e-005, 6.285837e-005, 3.210259e-005, 2.129255e-005, 
    7.503739e-006, 2.695655e-006, 4.287576e-006, 1.842256e-005, 
    1.331445e-005, 1.733728e-005, 6.399583e-006, 7.668423e-006, 
    2.963061e-007, 1.097948e-005, 2.631398e-005, 2.120636e-005, 
    1.716442e-005, 1.08354e-005, 2.686706e-006, 9.737996e-007, 5.158559e-006, 
    5.881266e-006, 5.908514e-007, -4.367503e-006, -4.601934e-006, 
    -5.269259e-006, -4.780512e-006, -3.541727e-006, -1.867083e-006, 
    -1.184857e-006, -1.518893e-006, -1.965431e-006, -1.783636e-006, 
    -1.45581e-006, -1.280224e-006, 3.686083e-006, 7.96172e-006, 
    1.887485e-005, 1.657582e-005, 3.685338e-006, 5.029422e-006, 
    -1.949229e-007, 4.509602e-006, 8.628267e-007, 1.269209e-005, 
    1.32971e-006, -1.647544e-005, -1.749839e-005, -1.046654e-005, 
    -1.13195e-006, -3.86899e-007, 9.576979e-007, 1.787681e-006, 
    6.412753e-006, 4.806901e-006, 7.606579e-006, 4.209361e-006, 5.577785e-006,
  5.072394e-006, 7.931925e-006, 3.304871e-006, -5.869782e-006, 
    -1.370258e-005, -1.16045e-005, -9.696902e-006, 5.985348e-006, 
    2.975095e-005, 4.546422e-005, 3.543475e-005, 1.564377e-005, 
    9.159536e-006, 6.568713e-006, 4.12493e-006, 6.665083e-006, 6.467635e-006, 
    -5.159993e-006, -1.14314e-006, 5.78566e-006, 6.722694e-006, 
    4.649955e-006, 7.501534e-006, 3.141206e-006, 6.367314e-006, 
    1.560431e-006, -4.01483e-006, 5.00086e-006, 5.035363e-006, 1.116424e-005, 
    7.223876e-006, 4.991656e-006, 7.832576e-006, 4.59305e-006, 8.780546e-006, 
    7.217408e-006, 7.07958e-006, 1.747412e-005, -1.653214e-006, 
    3.414926e-005, 9.796073e-006, 2.065924e-005, 1.826935e-006, 
    -2.506521e-005, -1.44993e-005, -2.137e-005, -2.586715e-005, 
    -2.533321e-005, -3.177374e-005, -3.410278e-005, -2.794836e-005, 
    -2.078683e-005, -1.819778e-005, -5.87129e-006, 1.342865e-006, 
    7.416238e-007, 1.040403e-005, 1.428131e-005, 1.628328e-005, 
    1.820975e-005, 1.414769e-005, 7.47868e-006, 9.531068e-006, 1.456543e-005, 
    1.288631e-005, 1.356407e-005, 1.117741e-005, 8.562984e-006, 
    9.346539e-006, 1.201608e-005, 1.002479e-005, 1.728811e-005, 
    1.581166e-005, 1.542646e-005, 1.180771e-005, 7.45161e-006, 4.272194e-006, 
    4.517329e-006, 5.197558e-006, 7.232302e-006, 1.814253e-006, 
    4.074485e-006, 5.843009e-006, 3.58923e-006, -5.820599e-006, 
    -7.653936e-006, -1.314998e-005, -8.411167e-006, -3.157016e-006, 
    1.802837e-006, -6.538685e-007, 2.846537e-007, -1.32393e-006, 
    6.085029e-007, 5.931033e-007, 3.170513e-006,
  -1.557131e-006, 1.69182e-006, -9.397299e-007, -5.582442e-006, 
    -1.233664e-005, -1.034262e-005, -1.011736e-005, -2.130838e-005, 
    1.671664e-005, 4.863643e-005, 1.728389e-005, 3.597421e-006, 
    4.469883e-006, 2.381981e-006, 5.044385e-007, 7.432238e-006, 
    1.322979e-005, 1.397832e-005, 1.097126e-005, 6.415732e-006, 
    5.651313e-006, 6.606722e-006, 8.198658e-006, 3.209134e-007, 
    -4.566755e-007, 4.754755e-006, 1.53162e-005, 7.259638e-006, 
    -7.456249e-006, 4.986716e-006, 1.061264e-005, 3.584748e-006, 
    -4.066256e-006, 9.358686e-006, 1.455274e-005, 1.766573e-006, 
    3.581525e-006, 1.922725e-005, 1.983894e-005, 2.442699e-005, 
    1.490119e-005, 2.841532e-005, -8.727322e-006, -2.9661e-005, 
    -2.291846e-005, -2.459309e-005, -3.478798e-005, -3.484982e-005, 
    -3.252771e-005, -3.431286e-005, -3.630912e-005, -3.234392e-005, 
    -2.557085e-005, -2.154977e-005, -1.495776e-005, -8.465815e-006, 
    -2.163866e-006, 8.471616e-007, 3.618033e-006, 6.040714e-006, 
    7.370641e-006, 7.310791e-006, 7.880013e-006, 9.722542e-006, 
    1.063797e-005, 1.080213e-005, 1.04907e-005, 9.792579e-006, 1.182087e-005, 
    1.739788e-005, 1.579452e-005, 2.302208e-005, 2.060486e-005, 
    2.302878e-005, 1.324295e-005, 7.2482e-006, 1.253067e-005, 3.914807e-006, 
    5.071881e-006, 1.445987e-005, 1.610447e-005, 4.117718e-006, 
    2.036832e-007, -3.721038e-006, -4.724381e-006, -3.65571e-006, 
    -1.883469e-006, 3.176719e-006, 3.433761e-006, 3.514724e-006, 
    2.398636e-006, -2.02503e-006, -1.853663e-006, -1.010008e-006, 
    -1.670382e-006, 2.485056e-006,
  -5.022404e-006, -1.86931e-006, -5.061633e-006, -1.094908e-005, 
    -8.956304e-006, -1.057946e-006, -7.605009e-006, -9.395386e-006, 
    2.730929e-006, 1.748357e-005, 1.056346e-005, 1.375411e-006, 7.64712e-007, 
    1.725338e-006, 8.024306e-006, 1.37995e-005, 1.068615e-005, 7.110615e-006, 
    7.135697e-006, 5.220903e-006, 3.1253e-006, 1.965991e-006, 2.425444e-006, 
    2.761961e-006, 4.11152e-006, 1.14635e-005, 7.689014e-006, -1.48892e-005, 
    -4.641424e-006, -1.416069e-006, 7.599876e-006, 3.930705e-006, 
    -7.963135e-006, 6.004215e-006, 1.578632e-005, 1.193661e-005, 
    7.267066e-006, 1.067123e-005, 1.634214e-005, 1.590081e-005, 
    1.471566e-005, 1.108574e-005, 3.141933e-006, 2.983739e-006, 3.46241e-007, 
    4.627145e-007, -3.151308e-006, -7.984745e-006, -1.281521e-005, 
    -1.502181e-005, -1.552473e-005, -1.682834e-005, -1.588336e-005, 
    -1.557442e-005, -1.389977e-005, -1.191444e-005, -6.325265e-006, 
    -2.287296e-006, 2.598099e-007, 1.186663e-006, 1.576825e-006, 
    3.523412e-006, 4.253569e-006, 3.657026e-006, 3.42879e-006, 4.855825e-006, 
    3.179197e-006, 5.559656e-006, 1.012562e-005, 1.567705e-005, 
    1.882219e-005, 1.990103e-005, 2.090314e-005, 2.588808e-005, 
    1.770732e-005, 1.223687e-005, 1.591472e-005, 1.198156e-005, 
    1.369148e-005, 8.577387e-006, 2.615684e-006, -9.334667e-008, 
    -1.530315e-006, -2.451455e-006, -3.471442e-006, -3.666646e-006, 
    -3.514158e-006, -3.059176e-006, -2.810328e-006, -1.048264e-006, 
    1.126558e-006, 4.839185e-006, 3.272831e-006, -2.852175e-008, 
    -1.888679e-006, -4.054069e-006,
  -1.089727e-006, 1.770277e-006, -2.145483e-006, -8.270361e-006, 
    -3.890407e-006, -4.730085e-006, -6.890503e-006, -2.052846e-006, 
    1.436507e-006, 9.340825e-006, 7.255407e-006, 5.548527e-007, 
    -4.117348e-007, -6.593423e-007, 2.663613e-006, 5.092504e-006, 
    7.891437e-006, 6.909948e-006, 8.062554e-006, 8.036476e-006, 
    4.327574e-006, 1.626491e-006, -1.902081e-007, 3.278565e-007, 
    -1.399676e-006, 2.226028e-006, -5.433423e-006, -8.15463e-006, 
    1.750668e-006, 5.332666e-006, 2.419492e-006, -3.554636e-006, 
    1.009731e-005, 1.44991e-005, 1.190781e-005, 2.38861e-005, 2.203984e-005, 
    2.234208e-005, 1.869701e-005, 1.955409e-005, 2.451319e-005, 
    2.425714e-005, 2.032497e-005, 2.108592e-005, 2.187022e-005, 
    1.977635e-005, 1.51791e-005, 1.591174e-005, 1.474672e-005, 1.385812e-005, 
    1.205383e-005, 8.636751e-006, 5.924743e-006, 1.942906e-006, 
    -1.606804e-006, -2.785735e-006, -7.784078e-006, -7.959658e-006, 
    -8.59196e-006, -5.51041e-006, -2.764125e-006, -3.088473e-006, 
    -2.957102e-006, -1.22534e-006, 9.216819e-008, 4.981244e-006, 
    5.218666e-006, 9.528085e-006, 1.332043e-005, 1.941079e-005, 
    1.313143e-005, 1.44492e-005, 1.708447e-005, 2.06893e-005, 1.367854e-005, 
    6.72444e-006, 6.248587e-006, 4.265243e-006, 5.767774e-006, 4.997196e-007, 
    -4.065198e-007, -1.392923e-007, -3.543655e-007, -2.121645e-006, 
    -2.022553e-006, -6.106675e-007, -1.25415e-006, -1.5102e-006, 
    -1.391735e-006, -1.399434e-006, -1.443392e-006, 1.386124e-007, 
    -4.691046e-007, -1.851178e-006, 2.882171e-006, 4.010693e-006,
  5.456623e-007, 3.004352e-006, 1.221927e-006, -9.988426e-007, 
    -2.184477e-006, -1.619723e-006, -2.919105e-006, -2.097305e-006, 
    -5.043712e-007, -1.446129e-006, -1.088527e-005, -4.745242e-006, 
    -7.586837e-007, -2.85572e-007, -1.359947e-006, -1.290904e-006, 
    -1.287675e-006, 1.327975e-006, 3.78617e-006, 1.317191e-005, 
    1.354171e-005, 3.875328e-006, 2.781828e-006, 4.069538e-006, 
    3.032665e-006, 4.746551e-006, -3.081283e-006, -2.670751e-006, 
    -7.874933e-007, -1.495546e-006, 1.344597e-008, 1.049822e-006, 
    2.732908e-006, 3.305357e-006, 9.957985e-006, 1.515776e-005, 
    8.803396e-006, 1.002553e-005, 1.028829e-005, 1.16736e-005, 1.184049e-005, 
    9.966674e-006, 8.438064e-006, 1.13351e-005, 8.898507e-006, 9.356967e-006, 
    8.777311e-006, 6.941489e-006, 6.674263e-006, 4.904997e-006, 
    4.078975e-006, 4.958887e-006, 3.586243e-006, -1.593149e-006, 
    -6.037668e-006, -6.32079e-006, -1.192636e-005, -1.243996e-005, 
    -1.345373e-005, -1.42045e-005, -1.375796e-005, -9.549873e-006, 
    -7.965882e-006, -8.152147e-006, -7.812892e-006, -5.972604e-006, 
    1.930039e-007, 6.826005e-006, 1.019391e-005, 9.792826e-006, 
    6.378476e-006, 8.145258e-006, 5.908591e-006, 3.635917e-006, 
    3.670932e-006, 2.717509e-006, 4.674527e-006, 3.877813e-006, 1.12786e-007, 
    -9.198643e-007, 2.883698e-007, -4.425337e-007, -1.274514e-006, 
    -1.3366e-006, -8.190345e-007, -7.259023e-007, -1.254894e-006, 
    -7.169615e-007, -1.094207e-006, -5.600017e-007, -5.751511e-007, 
    -5.806151e-007, -2.022303e-006, -4.854517e-006, -2.631265e-006, 
    -5.992424e-007,
  -5.609945e-007, 8.695747e-008, -4.450144e-007, -4.748164e-007, 
    -9.235328e-008, -6.615776e-007, -1.421537e-006, -4.69601e-007, 
    5.74722e-007, -9.320338e-007, -3.016705e-006, -1.254147e-006, 
    -1.082287e-006, -2.135497e-007, -1.724278e-006, -1.493807e-006, 
    -1.248435e-006, -6.297887e-007, 1.224718e-007, 4.178567e-006, 
    3.171745e-006, 4.468643e-006, 4.533213e-006, 7.748138e-006, 
    2.295804e-006, 2.048942e-006, 2.653183e-006, -9.789728e-007, 
    -4.582822e-006, -2.865957e-006, 1.890267e-007, 2.277923e-006, 
    1.226398e-006, 1.469038e-006, 3.954305e-006, 3.768038e-006, 
    4.422448e-006, 5.834083e-006, 3.813736e-006, 2.854847e-006, 3.70297e-006, 
    3.519935e-006, 1.861931e-006, -2.28204e-007, 3.57164e-007, 3.77795e-008, 
    9.715868e-007, 7.180197e-007, 5.980646e-007, -7.544641e-007, 
    -1.286681e-006, -2.222724e-006, -7.420458e-007, -1.459537e-006, 
    -6.047107e-006, -7.954954e-006, -7.36611e-006, -9.291092e-006, 
    -1.133478e-005, -9.832993e-006, -8.972451e-006, -7.486807e-006, 
    -3.65547e-006, -2.842611e-006, -1.417068e-006, -2.848572e-006, 
    -3.657457e-006, -9.824525e-007, 4.376758e-006, 6.308441e-006, 
    5.369666e-006, 4.320873e-006, 6.611488e-007, -7.467622e-007, 
    -6.074388e-007, 2.544904e-006, 3.174477e-006, 3.115618e-006, 
    5.344887e-007, -8.014013e-007, -1.078562e-006, -8.033885e-007, 
    -5.232441e-007, -1.482136e-006, -1.564342e-006, -1.037089e-006, 
    -5.239917e-007, -1.337096e-006, -1.072105e-006, -4.939397e-007, 
    -2.82095e-007, -1.296063e-007, -1.969099e-007, -3.439348e-007, 
    -6.042084e-007, -9.605943e-007,
  -4.753132e-007, -4.169505e-007, -9.92632e-007, -1.145121e-006, 
    -7.239141e-007, -9.359508e-008, -5.96509e-007, -4.966714e-007, 
    -3.898799e-007, -4.648825e-007, -1.133945e-006, -8.587698e-007, 
    -1.903093e-006, -2.152688e-006, -3.002245e-007, -9.186228e-007, 
    -1.123514e-006, -2.083341e-007, 1.150211e-007, 7.599932e-007, 
    2.483809e-006, 2.55757e-006, 5.319747e-006, 7.420561e-006, 2.968841e-006, 
    6.894606e-007, 1.121098e-006, 2.677028e-006, 6.310966e-007, 
    -4.897979e-006, -3.597854e-006, -2.197642e-006, -1.484122e-006, 
    -1.441156e-006, -4.681115e-007, -9.665564e-007, -5.977536e-007, 
    -4.231597e-007, -2.870629e-007, 3.246305e-007, 1.9347e-006, 
    2.865278e-006, 2.189013e-006, -7.499912e-007, -9.193682e-007, 
    -1.078316e-006, -6.258151e-007, -4.693529e-007, 5.687616e-007, 
    5.652828e-007, -4.86737e-007, -7.209337e-007, 1.567969e-008, 
    2.140583e-006, 5.404472e-007, -2.584577e-006, -4.778523e-006, 
    -3.757297e-006, -6.146698e-006, -5.281188e-006, -7.245906e-006, 
    -8.66524e-006, -6.929507e-006, -4.969255e-006, -3.395445e-006, 
    -3.107853e-006, -2.942449e-006, -5.438641e-006, -6.965018e-006, 
    -3.643053e-006, -1.548942e-006, -4.052781e-007, -2.680436e-006, 
    -1.250175e-006, 2.791821e-007, 1.438493e-006, 7.570125e-007, 
    7.80854e-007, 9.852492e-007, 9.94437e-007, 5.91408e-008, 3.79765e-007, 
    7.013814e-007, 1.368753e-007, -1.308481e-007, -1.331636e-006, 
    -1.1558e-006, -1.465496e-006, -1.233534e-006, -1.029388e-006, 
    -6.968438e-007, -3.878932e-007, -3.941018e-007, -7.052879e-007, 
    -5.756479e-007, -1.104833e-007,
  -5.982478e-007, -8.838533e-007, -6.024699e-007, -7.534682e-007, 
    -1.174675e-006, -1.394715e-006, -1.05025e-006, -5.776344e-007, 
    -3.032046e-007, -3.598292e-007, -1.373109e-006, -1.837776e-006, 
    -2.794182e-006, -2.327528e-006, -1.985049e-006, -1.256382e-006, 
    -3.484048e-007, 4.140378e-007, 1.115442e-007, 4.445851e-007, 
    8.384726e-007, 1.597439e-006, 2.3646e-006, 4.403823e-006, 5.189363e-006, 
    6.258521e-006, 5.01353e-006, 6.477317e-006, 2.819083e-006, 
    -3.821824e-007, -2.689627e-006, -2.414204e-006, -1.881735e-006, 
    -2.999074e-006, -3.142373e-006, -3.608285e-006, -2.055086e-006, 
    4.523372e-008, 7.458375e-007, 5.72486e-007, -1.541948e-007, 
    1.014802e-006, -7.981726e-007, -2.155666e-006, -2.086377e-006, 
    -1.277243e-006, -1.953509e-006, -7.308681e-007, -1.360622e-007, 
    1.251483e-006, 2.131645e-006, 1.049076e-006, 1.394073e-008, 
    -1.610038e-006, 7.083345e-007, -1.402417e-006, -3.748853e-006, 
    -5.108088e-006, -6.558963e-006, -4.875877e-006, -4.011361e-006, 
    -4.819749e-006, -5.790062e-006, -2.960578e-006, -2.714212e-006, 
    -2.486722e-006, -3.751831e-006, -4.133549e-006, -4.507817e-006, 
    -4.822728e-006, -9.591591e-006, -4.260957e-006, -2.225705e-006, 
    -1.310775e-006, -2.763387e-006, -1.209693e-006, 4.527792e-007, 
    1.014554e-006, 1.743469e-006, 1.630716e-006, 8.255583e-007, 
    2.560798e-006, 2.305739e-006, 1.041625e-006, 6.802702e-007, 
    -3.089181e-007, -9.618379e-007, -6.730029e-007, -3.590844e-007, 
    -1.03063e-006, -8.831087e-007, -9.839396e-007, -7.514816e-007, 
    -7.281365e-007, -9.988408e-007, -9.476801e-007,
  -4.482425e-007, -6.11162e-007, -9.618362e-007, -1.057949e-006, 
    -9.648164e-007, -6.677864e-007, -8.386532e-007, -8.518159e-007, 
    -4.723332e-007, -2.132447e-008, -6.171227e-007, -9.593529e-007, 
    -1.581973e-006, -3.531541e-006, -4.20855e-006, -2.778287e-006, 
    -3.365393e-006, -1.477664e-006, -6.454347e-007, -4.964232e-007, 
    -3.220796e-007, 1.433277e-006, 2.860063e-006, 2.478841e-006, 
    1.950595e-006, 3.642622e-006, 4.234694e-006, 7.106397e-006, 
    7.865114e-006, 6.128881e-006, 1.498593e-006, 1.653312e-006, 
    -8.664574e-008, -1.603086e-006, -2.48747e-006, -4.417167e-006, 
    -3.896123e-006, -3.023413e-006, -3.861551e-007, 3.670984e-007, 
    3.785217e-007, -2.344123e-007, -4.402973e-007, -2.378441e-006, 
    -2.133317e-006, -5.84743e-006, -4.262693e-006, -2.833671e-006, 
    -1.25862e-006, -3.001696e-008, 1.372678e-006, 8.983252e-007, 
    3.146952e-007, -6.685314e-007, 1.223419e-006, 3.894493e-007, 
    -6.978371e-007, -4.577603e-006, -4.317084e-006, -3.036575e-006, 
    -2.487467e-006, -1.402661e-006, -2.087123e-006, -2.558496e-006, 
    -9.648184e-007, -3.692676e-007, -1.015433e-007, -1.964933e-006, 
    -3.02987e-006, -4.374453e-006, -8.016546e-006, -3.537754e-006, 
    -5.587626e-007, -1.941095e-006, -4.226933e-006, -5.885679e-006, 
    -2.63201e-006, 6.606479e-007, 2.723466e-006, 4.647703e-006, 
    2.241914e-006, 1.017535e-006, 7.301896e-007, 3.521424e-006, 
    1.886024e-006, 6.152022e-007, -7.174604e-007, -7.244125e-007, 
    -5.7242e-007, -5.120696e-007, -2.075885e-007, -1.179642e-006, 
    -1.069373e-006, -1.183615e-006, -1.417812e-006, -8.185366e-007,
  -5.485219e-008, -1.859235e-008, -8.071124e-007, -1.448856e-006, 
    -2.109474e-006, -1.539505e-006, -1.016723e-006, -6.022212e-007, 
    -2.853233e-007, 2.250415e-007, 1.99213e-007, -3.275431e-007, 
    -1.083528e-006, -2.294249e-006, -4.238851e-006, -4.282312e-006, 
    -5.197244e-006, -5.413807e-006, -3.165221e-006, -2.35882e-006, 
    -1.527832e-006, 9.340874e-007, 2.558066e-006, 2.458476e-006, 
    1.562917e-006, 5.104174e-006, 8.606446e-006, 5.891951e-006, 
    8.562986e-006, 1.116126e-005, 7.149371e-006, 3.296918e-006, 
    -2.357818e-006, -4.172278e-006, -3.704637e-006, -2.458648e-006, 
    -1.437427e-006, -2.49492e-006, -4.212776e-006, -3.256369e-006, 
    -4.708436e-007, -7.546805e-008, 6.663631e-007, 1.469285e-006, 
    1.512781e-007, -2.375462e-006, -6.025002e-006, -5.262807e-006, 
    -3.260094e-006, -2.982682e-006, -1.066889e-006, -8.11583e-007, 
    -1.740918e-006, -7.860035e-007, -1.914468e-007, -1.641827e-006, 
    -7.072758e-007, -2.750223e-006, -2.446492e-006, -2.204843e-006, 
    -1.200257e-006, -2.775309e-006, -2.2791e-006, -1.646298e-006, 
    -1.390246e-006, -3.516334e-007, 1.317048e-006, 1.127554e-006, 
    -2.720174e-006, -2.253023e-006, -5.531529e-006, -4.637212e-006, 
    -1.767243e-006, 3.528381e-006, 1.448674e-006, -5.805708e-006, 
    -3.102134e-006, -9.807118e-007, 2.308223e-006, 3.163299e-006, 
    3.788649e-006, -3.265504e-007, -1.256882e-006, -9.53889e-007, 
    -8.259904e-007, -1.332131e-006, -1.215405e-006, 6.112714e-008, 
    -7.884873e-007, -1.406885e-006, -1.129972e-006, -1.121031e-006, 
    -5.674519e-007, -9.253285e-007, -8.326926e-007, -4.606603e-007,
  -1.022185e-006, -7.216786e-007, 3.010373e-007, 1.717035e-008, 
    -1.409865e-006, -1.703666e-006, -2.781268e-006, -3.393706e-006, 
    -2.962566e-006, -3.136662e-006, -1.83281e-006, -4.236554e-007, 
    -5.133111e-007, -2.129343e-006, -2.969519e-006, -3.548927e-006, 
    -4.098282e-006, -8.206534e-006, -1.224996e-005, -7.314202e-006, 
    -4.278339e-006, -6.900696e-006, -4.159629e-006, -1.042745e-007, 
    -2.525963e-006, -3.978825e-006, 2.675785e-006, 7.033875e-006, 
    1.048672e-005, 1.075818e-005, 1.611603e-006, 1.770299e-006, 
    -3.514149e-006, -4.711961e-006, -6.355549e-006, -4.068475e-006, 
    -6.400755e-006, -5.061378e-006, -6.397095e-007, -5.085858e-007, 
    -3.589899e-006, -2.316843e-006, -1.571287e-006, -1.715089e-006, 
    3.91134e-006, 4.834714e-006, 2.325858e-006, -9.12667e-007, -3.0557e-006, 
    -3.978332e-006, -3.464491e-006, -1.715094e-006, -3.433943e-006, 
    -2.817778e-006, -1.345046e-006, -2.01709e-006, -5.152546e-006, 
    -4.443247e-006, -3.790079e-006, -2.720177e-006, -1.713106e-006, 
    -1.25067e-006, -1.236764e-006, -3.851619e-007, 1.31954e-008, 
    -1.263775e-007, -1.099875e-007, -2.138004e-007, -4.322545e-006, 
    -1.681812e-006, -2.496408e-006, -6.622542e-006, -4.470308e-006, 
    -5.224058e-006, -3.359677e-006, -1.675347e-006, -4.173766e-006, 
    -2.059303e-006, -4.592246e-006, -7.071558e-006, -2.80088e-006, 
    -2.089353e-006, -3.435678e-006, -6.772299e-006, -4.878113e-006, 
    -4.755922e-006, -4.714198e-006, -5.889404e-006, -4.012351e-006, 
    -4.250772e-006, -4.249282e-006, -2.25948e-006, -2.091842e-006, 
    -1.602835e-006, 6.082496e-007, 6.330847e-007,
  4.026515e-008, -2.222474e-006, -3.010746e-006, -2.666779e-006, 
    -3.816858e-007, -1.318971e-006, -1.609791e-006, -5.999864e-007, 
    -2.30642e-006, -6.716913e-006, -4.059292e-006, -4.496145e-006, 
    -4.854019e-006, -8.033928e-006, -4.654594e-006, -3.544207e-006, 
    -3.203468e-006, -5.847187e-006, -1.155184e-005, -1.106433e-005, 
    -8.363742e-006, -3.050485e-006, -8.736715e-007, -1.38547e-007, 
    2.208171e-007, 2.257848e-007, -1.087504e-006, 1.933209e-006, 
    6.840908e-006, 9.051495e-006, 7.143402e-006, 6.158185e-006, 
    3.792877e-006, 2.214849e-006, 1.243545e-006, 1.946377e-006, 
    3.678142e-006, 1.095519e-006, -2.888301e-006, -9.918949e-007, 
    1.163571e-006, -1.191656e-007, -4.22413e-007, 1.426575e-006, 
    -5.952606e-007, 1.917077e-006, 4.070294e-006, 4.981746e-006, 
    8.103292e-006, 6.444046e-006, 3.490881e-006, 1.625009e-006, 
    3.050118e-007, -2.041423e-006, -2.251283e-006, -8.297138e-007, 
    -2.844103e-006, -4.510053e-006, -2.135053e-006, -1.734959e-006, 
    1.213977e-006, 3.378622e-006, 1.972448e-006, 3.151128e-006, 
    2.013178e-006, 1.88354e-006, 1.219443e-006, -7.81286e-007, 
    -3.342048e-006, -3.237739e-006, -1.367398e-006, -2.922832e-006, 
    -6.983355e-007, 4.008703e-006, 1.846045e-006, -2.641194e-006, 
    -3.068351e-006, 1.416898e-006, -2.224951e-006, -4.975707e-006, 
    -9.470634e-006, -1.559616e-006, -5.94329e-006, -7.758998e-006, 
    -1.212603e-005, -1.241511e-005, -1.069998e-005, -9.576699e-006, 
    -7.754037e-006, -6.522952e-006, -4.36849e-006, -2.293007e-006, 
    -1.302824e-006, -1.025913e-006, 9.800297e-007, 1.504553e-006,
  1.449418e-006, 6.792779e-007, 6.854843e-007, 2.768169e-006, 2.865523e-006, 
    -1.350727e-007, 6.57421e-007, 1.145931e-006, -3.499008e-008, 
    -2.294251e-006, -5.796228e-007, -1.751599e-006, -2.470081e-006, 
    -1.144128e-006, -1.822379e-006, -2.08886e-006, -8.766519e-007, 
    -7.840154e-007, 1.109671e-006, 6.358205e-007, 9.415635e-008, 
    1.947118e-006, 1.926754e-006, 3.766055e-006, 1.706465e-006, 
    2.170635e-006, 7.743956e-007, -1.101909e-006, 2.036028e-006, 
    3.186896e-006, 4.55333e-006, 4.65863e-006, 4.953175e-006, 4.950696e-006, 
    4.674275e-006, 6.823524e-006, 6.884129e-006, 6.403312e-006, 
    3.851739e-006, 3.282767e-006, 9.69573e-006, 1.023217e-005, 7.381823e-006, 
    4.87495e-006, 5.014779e-006, 4.35987e-006, 4.691668e-006, 4.718735e-006, 
    3.929723e-006, 6.76393e-006, 9.423533e-006, 8.614894e-006, 5.444184e-006, 
    4.489768e-006, 1.37815e-006, 7.152958e-007, -1.530309e-006, 
    -1.466975e-006, -4.067697e-007, 1.692024e-008, 2.628101e-006, 
    4.620886e-006, 6.224247e-006, 7.971164e-006, 7.716353e-006, 
    4.133861e-006, 5.267343e-006, 2.681496e-006, -1.53131e-006, 
    -2.902465e-006, -7.298513e-008, 3.477715e-006, 3.708188e-006, 
    8.583844e-006, 9.742169e-006, 1.099089e-005, 1.009881e-005, 
    9.566589e-006, 1.209804e-005, 9.960473e-006, 7.958501e-006, 
    3.645859e-006, -3.411988e-007, -5.736663e-006, -9.084451e-006, 
    -1.346191e-005, -1.013945e-005, -1.104396e-005, -8.716888e-006, 
    -4.82571e-006, -1.182872e-006, 2.292576e-006, 1.758615e-006, 
    2.210869e-006, 4.078231e-006, 2.302759e-006,
  2.858569e-006, 3.501061e-006, 6.023331e-006, 7.663699e-006, 4.727919e-006, 
    5.340111e-006, 5.996009e-006, 4.258036e-006, 4.938772e-006, 
    3.474983e-006, 1.700502e-006, 2.538194e-006, -1.037806e-007, 
    -3.150672e-008, 1.808339e-007, 1.220686e-006, 2.448046e-006, 
    3.093515e-006, 3.89793e-006, 5.492348e-006, 5.374633e-006, 3.934684e-006, 
    2.565765e-006, 1.580054e-006, 7.743977e-007, 9.241543e-007, 
    1.081362e-006, 5.911136e-007, 2.665163e-007, 8.00226e-007, 9.65877e-007, 
    8.998154e-007, 9.164551e-007, 6.551882e-007, 2.533525e-007, 
    1.006138e-007, 2.252589e-006, 4.309946e-006, 5.994276e-006, 
    5.039605e-006, 5.121816e-006, 9.152336e-006, 1.074502e-005, 
    1.000219e-005, 1.183652e-005, 1.170813e-005, 7.678111e-006, 
    6.950442e-006, 7.34135e-006, 6.52079e-006, 7.164519e-006, 6.625094e-006, 
    6.027807e-006, 1.031587e-005, 7.623232e-006, 6.780567e-006, 
    6.438091e-006, 5.04309e-006, 3.70944e-006, 3.455127e-006, 2.447548e-006, 
    4.649191e-006, 5.805774e-006, 8.725667e-006, 8.405783e-006, 
    6.235918e-006, 4.151746e-006, 2.569989e-006, 2.143815e-006, 
    2.704842e-006, 2.885146e-006, 4.129643e-006, 7.303586e-006, 
    6.160668e-006, 6.145767e-006, 5.57282e-006, 6.814833e-006, 5.174712e-006, 
    7.044564e-006, 1.035237e-005, 7.594666e-006, 5.229351e-006, 
    3.477475e-006, 2.692432e-006, 5.247981e-006, 3.252466e-006, 
    -1.041302e-006, -8.559437e-006, -4.982663e-006, -1.286429e-006, 
    4.922658e-007, 1.184673e-006, 4.089407e-006, 7.200275e-006, 
    9.561118e-006, 4.833972e-006,
  4.255304e-006, 3.289462e-006, 7.230819e-006, 7.67239e-006, 2.973062e-006, 
    2.68547e-006, 6.262491e-006, 4.69017e-006, 3.594938e-006, 4.301996e-006, 
    5.135468e-006, 4.911454e-006, 3.811747e-006, 1.897695e-006, 
    2.379747e-006, 3.606363e-006, 3.487899e-006, 3.118599e-006, 
    2.543414e-006, 3.099476e-006, 3.540797e-006, 4.199182e-006, 
    2.972816e-006, 2.512617e-006, 2.510879e-006, 2.285624e-006, 
    1.367712e-006, 1.087818e-006, 9.19187e-007, 6.681025e-007, 2.007023e-007, 
    1.686653e-007, 8.923644e-007, 4.13293e-007, 1.212293e-007, 
    -6.278051e-007, -9.047162e-007, -4.216727e-007, 1.627735e-006, 
    5.509733e-006, 6.999604e-006, 5.962731e-006, 4.309448e-006, 
    7.977873e-006, 9.406405e-006, 8.738334e-006, 7.190352e-006, 
    6.502163e-006, 4.577923e-006, 3.435252e-006, 3.086316e-006, 
    8.127379e-006, 7.42653e-006, 3.344598e-006, 2.713288e-006, 3.849502e-006, 
    8.219267e-006, 3.591962e-006, 1.279557e-006, 4.731402e-006, 3.96722e-006, 
    6.025402e-007, 1.914592e-006, 3.707701e-006, 6.65291e-006, 4.277406e-006, 
    2.504174e-006, 4.476838e-006, 3.376886e-006, 2.240423e-006, 
    8.275447e-007, 1.777741e-006, 4.981739e-006, 6.147258e-006, 
    7.247956e-006, 9.279976e-006, 6.120184e-006, 5.79187e-006, 6.408776e-006, 
    5.051777e-006, 5.152608e-006, 1.00161e-005, 9.463023e-006, 5.386315e-006, 
    4.826772e-006, 5.121568e-006, 5.025206e-006, 7.103263e-007, 
    -6.649108e-006, -4.561953e-006, 7.865638e-007, 5.12628e-006, 
    5.876802e-006, 6.688173e-006, 6.65936e-006, 5.624972e-006,
  1.929979e-006, 1.37069e-006, 8.570969e-007, 3.543528e-006, 2.555831e-006, 
    1.022006e-006, 1.778239e-006, 2.368572e-006, 3.706696e-006, 
    4.124673e-006, 2.210621e-006, 3.003361e-006, 3.184659e-006, 
    1.627488e-006, 2.278421e-006, 3.114129e-006, 2.826784e-006, 
    3.361985e-006, 4.287594e-006, 3.982617e-006, 3.113134e-006, 
    3.376636e-006, 3.944869e-006, 3.107175e-006, 2.512617e-006, 1.84132e-006, 
    1.532866e-006, 1.718137e-006, 2.009207e-006, 1.423591e-006, 
    8.260547e-007, 1.109674e-006, 1.504803e-006, 9.450155e-007, 
    7.140479e-007, 1.056278e-006, 1.199081e-006, -4.442154e-008, 
    1.670951e-006, 5.321483e-006, 6.564986e-006, 6.586093e-006, 
    5.051028e-006, 5.271319e-006, 4.626596e-006, 7.203998e-006, 
    9.690753e-006, 8.711995e-006, 9.367646e-006, 7.908075e-006, 
    5.557416e-006, 7.470484e-006, 5.399466e-006, 6.283106e-006, 
    2.363111e-006, 2.045221e-006, 2.666347e-006, 2.486791e-006, 
    1.288739e-006, 2.559555e-006, 2.461704e-006, 2.770917e-006, 
    3.847515e-006, 2.991448e-006, 4.03179e-006, 4.380477e-006, 2.412779e-006, 
    2.563778e-006, 2.26476e-006, 2.343241e-006, 2.647968e-006, 2.02212e-006, 
    1.462832e-006, 1.476242e-006, 3.977154e-006, 5.265355e-006, 
    4.861784e-006, 5.40791e-006, 5.056492e-006, 4.016394e-006, 7.050021e-006, 
    9.366408e-006, 5.668186e-006, 7.12353e-006, 7.206236e-006, 5.765294e-006, 
    3.258923e-006, -1.768731e-006, -6.054306e-006, -7.016173e-006, 
    -3.422261e-006, 1.786681e-006, 3.621513e-006, 3.848261e-006, 
    4.326084e-006, 3.66323e-006,
  1.539322e-006, 8.811858e-007, 1.237822e-006, 2.170884e-006, 1.57285e-006, 
    1.817478e-006, -2.48072e-007, -2.624765e-007, 1.436256e-006, 
    3.288718e-006, 1.7914e-006, 1.371934e-006, 3.284744e-006, 2.268237e-006, 
    2.085203e-006, 2.730173e-006, 1.260174e-006, 1.089059e-006, 
    2.303753e-006, 2.375029e-006, 2.43836e-006, 2.330326e-006, 3.774499e-006, 
    5.202028e-006, 3.768289e-006, 3.206265e-006, 3.558926e-006, 
    2.669824e-006, 2.205157e-006, 2.105319e-006, 1.594706e-006, 
    1.296435e-006, 9.626488e-007, 5.176007e-007, 6.387959e-007, 
    8.779598e-007, 1.043611e-006, 3.899468e-007, 2.544407e-006, 
    6.082438e-006, 9.001326e-006, 6.902001e-006, 5.446906e-006, 6.92038e-006, 
    6.244612e-006, 6.306209e-006, 4.676018e-006, 3.235569e-006, 2.65418e-006, 
    3.336903e-006, 5.799069e-006, 6.198174e-006, 5.983096e-006, 
    6.369039e-006, 5.212212e-006, 5.876307e-006, 6.921127e-006, 
    4.446543e-006, 3.144176e-006, 7.897943e-007, 1.03467e-006, 2.899069e-006, 
    6.078721e-006, 3.868125e-006, 1.999517e-006, 3.220669e-006, 
    3.158335e-006, 3.37167e-006, 1.439982e-006, 1.148167e-006, 1.945877e-006, 
    1.896455e-006, 1.12077e-008, 4.697176e-008, 7.445951e-007, 2.41402e-006, 
    3.749661e-006, 5.465529e-006, 6.589574e-006, 6.820293e-006, 
    5.975397e-006, 8.175057e-006, 8.665555e-006, 8.900748e-006, 
    8.048897e-006, 4.668565e-006, 1.683868e-006, 1.017535e-006, 
    -2.422399e-006, -4.848305e-006, -2.126111e-006, -8.190327e-007, 
    1.056023e-006, 2.532979e-006, 2.412278e-006, 1.782704e-006,
  1.758654e-007, -2.928049e-006, -1.306798e-006, 1.117371e-006, 
    3.589968e-006, 2.125187e-006, -8.838106e-008, 7.075887e-007, 
    3.224395e-006, 3.696515e-006, 2.058379e-006, 2.705587e-006, 
    2.099605e-006, 1.61507e-006, 1.658034e-006, 1.756383e-006, 2.028082e-006, 
    1.875842e-006, 2.488279e-006, 2.875462e-006, 2.921408e-006, 
    2.547883e-006, 1.662258e-006, 2.029819e-006, 1.815243e-006, 
    1.749182e-006, 1.239314e-006, 5.918578e-007, 7.453405e-007, 
    1.071676e-006, 1.093778e-006, 1.191629e-006, 1.266881e-006, 
    1.224661e-006, 6.512137e-007, 2.578226e-007, 7.99233e-007, 2.737183e-007, 
    1.184676e-006, 3.648087e-006, 2.52429e-006, 3.829928e-007, 2.567254e-006, 
    5.920011e-006, 7.924968e-006, 6.32011e-006, 6.231696e-006, 7.056973e-006, 
    9.336105e-006, 7.810972e-006, 5.630434e-006, 4.028312e-006, 
    4.155965e-006, 3.493607e-006, 3.334166e-006, 6.965081e-006, 
    7.870578e-006, 5.488131e-006, 4.192229e-006, 2.286615e-006, 2.09688e-006, 
    3.212233e-006, 4.780082e-006, 5.608828e-006, 2.918177e-006, 
    1.299663e-006, 1.461837e-006, 1.819217e-006, 1.172506e-006, 
    8.143825e-007, 2.193484e-006, 1.789413e-006, 1.204543e-006, 
    1.631213e-006, 1.940165e-006, 1.668714e-006, 1.802328e-006, 
    2.318653e-006, 7.49561e-007, -3.084206e-007, 9.415362e-007, 
    1.248996e-006, 2.999885e-006, 2.411536e-006, 4.259527e-006, 
    5.563379e-006, 6.413242e-006, 6.023081e-006, 2.683981e-006, 
    4.783578e-007, 6.643786e-007, 2.219811e-006, 3.002933e-007, 
    2.440349e-006, 2.249608e-006, 1.151642e-006,
  -3.232031e-006, -3.03906e-006, -3.779569e-007, 3.70769e-006, 4.15696e-006, 
    9.484902e-007, 5.645388e-007, 7.863182e-007, 8.404586e-007, 9.94436e-007, 
    6.944265e-007, 1.147918e-006, 1.408936e-006, 2.700869e-006, 
    2.758734e-006, 3.184411e-006, 3.274563e-006, 3.348076e-006, 2.1006e-006, 
    1.955811e-006, 2.371305e-006, 2.345972e-006, 2.387696e-006, 
    2.119476e-006, 1.284016e-006, 7.249746e-007, 6.229002e-007, 
    8.809402e-007, 5.317565e-007, 2.307529e-007, 3.315845e-007, 
    9.457608e-007, 1.012816e-006, 6.263795e-007, 3.51205e-007, 2.446614e-007, 
    1.74874e-007, 3.872156e-007, 6.690952e-007, 1.091792e-006, 2.301764e-006, 
    3.561659e-006, 4.490251e-006, 6.139313e-006, 6.91591e-006, 7.647804e-006, 
    7.093231e-006, 6.958624e-006, 7.094723e-006, 6.999356e-006, 
    6.208847e-006, 4.738104e-006, 2.640767e-006, 3.204033e-006, 
    3.532852e-006, 5.666197e-006, 5.003098e-006, 4.101334e-006, 
    3.868625e-006, 4.125166e-006, 3.890973e-006, 2.555334e-006, 
    2.437364e-006, 2.939038e-006, 2.576692e-006, 1.16282e-006, 6.541941e-007, 
    9.768037e-007, 1.136992e-006, 1.068943e-006, 1.941655e-006, 
    1.738999e-006, 1.664493e-006, 2.09762e-006, 2.153251e-006, 1.872116e-006, 
    1.361007e-006, 1.713961e-007, -2.652073e-007, -2.023753e-007, 
    1.199576e-006, 1.504553e-006, 1.360258e-006, 1.284263e-006, 3.38632e-006, 
    6.032276e-006, 6.261254e-006, 3.420846e-006, -7.254021e-007, 
    -4.658796e-007, 5.96574e-007, -9.53396e-007, -2.983927e-006, 
    -5.894124e-006, -2.790957e-006, -9.869236e-007,
  -7.600052e-006, -6.223194e-006, -3.091216e-006, -6.561158e-007, 
    1.110475e-007, -5.413767e-007, 1.810822e-007, 1.508528e-006, 
    2.445313e-006, 4.411077e-007, -3.729938e-007, -3.62279e-008, 
    5.918564e-007, 7.267117e-007, 6.397886e-007, 5.806819e-007, 
    9.037881e-007, 1.596941e-006, 1.951837e-006, 1.848275e-006, 
    1.069689e-006, 6.879704e-007, 1.058513e-006, 1.412414e-006, 
    1.207028e-006, 1.512998e-006, 1.742227e-006, 1.57459e-006, 1.330211e-006, 
    8.501454e-007, 8.004745e-007, 1.138234e-006, 1.290474e-006, 
    6.715804e-007, 3.902551e-008, 3.149453e-007, 2.983054e-007, 
    7.398764e-007, 1.615071e-006, 2.357397e-006, 4.120701e-006, 
    5.423062e-006, 5.212708e-006, 4.023843e-006, 3.188386e-006, 4.7843e-006, 
    7.08479e-006, 9.063911e-006, 7.658486e-006, 5.775723e-006, 4.138086e-006, 
    3.410661e-006, 3.108416e-006, 3.560666e-006, 3.521924e-006, 
    3.638151e-006, 2.973808e-006, 3.269348e-006, 2.511376e-006, 
    2.056145e-006, 2.046708e-006, 1.466059e-006, 1.166297e-006, 
    1.705223e-006, 1.891984e-006, 1.397017e-006, 8.277925e-007, 
    7.522931e-007, 9.276305e-007, 8.64798e-007, 1.179958e-006, 8.988222e-007, 
    1.291716e-006, 1.672689e-006, 2.001507e-006, 1.317047e-006, 
    1.144691e-006, 1.069689e-006, 8.516345e-007, 1.020763e-006, 
    1.602903e-006, 1.359515e-006, 2.692673e-006, 3.986338e-006, 
    5.013775e-006, 8.32705e-006, 7.391505e-006, 6.918144e-006, 5.689548e-006, 
    1.795372e-006, -2.246319e-006, -5.651733e-006, -5.483596e-006, 
    -5.204198e-006, -4.189927e-006, -4.904681e-006,
  -5.461494e-006, -7.965882e-006, -8.912599e-006, -6.263177e-006, 
    -2.786484e-006, -5.808643e-007, 8.046945e-007, 1.784695e-006, 
    2.128415e-006, 1.630468e-006, 1.08434e-006, 1.360012e-006, 1.820457e-006, 
    1.53982e-006, 1.357776e-006, 1.512253e-006, 1.262907e-006, 9.253959e-007, 
    8.086708e-007, 9.7159e-007, 1.318041e-006, 1.119607e-006, 7.311837e-007, 
    9.532105e-007, 8.161196e-007, 1.27458e-006, 1.738999e-006, 1.342877e-006, 
    8.441848e-007, 7.393792e-007, 1.013809e-006, 1.360261e-006, 
    1.318539e-006, 1.136247e-006, 1.098001e-006, 9.412909e-007, 
    1.437499e-006, 2.244396e-006, 3.36844e-006, 3.74991e-006, 3.953311e-006, 
    3.708187e-006, 3.402962e-006, 2.887382e-006, 2.771897e-006, 
    3.026459e-006, 4.099094e-006, 4.539673e-006, 4.7694e-006, 3.987584e-006, 
    2.573961e-006, 2.175107e-006, 2.224529e-006, 3.190372e-006, 
    3.058745e-006, 1.818969e-006, 1.379881e-006, 1.663996e-006, 
    1.731548e-006, 1.385842e-006, 1.052553e-006, 8.744837e-007, 
    8.953457e-007, 8.034549e-007, 7.085841e-007, 5.31757e-007, 5.411939e-007, 
    9.782948e-007, 1.242045e-006, 1.309349e-006, 1.814002e-006, 
    2.623382e-006, 1.890245e-006, 1.000647e-006, 7.840831e-007, 
    1.237079e-006, 1.443956e-006, 1.408938e-006, 9.313558e-007, 2.77691e-007, 
    8.133889e-007, 9.681121e-007, 1.454635e-006, 2.921903e-006, 
    3.488146e-006, 4.06954e-006, 4.593565e-006, 5.744926e-006, 6.296767e-006, 
    3.883522e-006, 1.084836e-006, -5.530474e-007, -1.440163e-006, 
    -3.552403e-006, -3.926422e-006, -3.88147e-006,
  -1.415079e-006, -2.168585e-006, -5.127455e-006, -6.531145e-006, 
    -4.671483e-006, -2.396571e-006, 1.49339e-008, 2.535464e-006, 
    4.127904e-006, 3.810756e-006, 3.153368e-006, 2.354913e-006, 
    1.460844e-006, 7.763838e-007, 4.912745e-007, 3.010364e-007, 5.53363e-007, 
    8.404581e-007, 8.176107e-007, 6.263795e-007, 4.321682e-007, 
    4.411086e-007, 7.522949e-007, 7.351578e-007, 8.332572e-007, 
    7.699273e-007, 5.809311e-007, 2.459033e-007, 1.1676e-007, 6.318428e-007, 
    7.431051e-007, 7.726587e-007, 8.332574e-007, 1.247261e-006, 
    1.684114e-006, 1.687342e-006, 1.66052e-006, 1.658285e-006, 1.746947e-006, 
    1.562173e-006, 1.374666e-006, 1.573597e-006, 1.823936e-006, 
    1.548761e-006, 1.604889e-006, 1.81872e-006, 2.182556e-006, 1.840078e-006, 
    1.724098e-006, 1.679891e-006, 1.667225e-006, 1.665984e-006, 
    1.581544e-006, 1.648847e-006, 1.304134e-006, 8.156239e-007, 9.06025e-007, 
    9.899682e-007, 9.010573e-007, 6.740627e-007, 8.498973e-007, 
    1.163814e-006, 1.195604e-006, 1.133764e-006, 9.159589e-007, 
    7.363999e-007, 7.329229e-007, 1.422846e-006, 1.499339e-006, 
    1.617307e-006, 1.698021e-006, 1.695786e-006, 1.601412e-006, 
    1.514985e-006, 1.469039e-006, 1.269116e-006, 1.313571e-006, 6.75057e-007, 
    -3.397117e-007, -3.605733e-007, 1.475555e-007, 5.498864e-007, 
    7.619797e-007, 9.154614e-007, 9.097498e-007, 7.244785e-007, 
    3.551784e-007, 7.354583e-008, -9.508585e-008, -8.887673e-008, 
    6.209148e-007, 1.954886e-007, -1.332379e-006, -1.887696e-006, 
    -2.11171e-006, -1.852181e-006,
  3.067489e-007, 1.065217e-006, 9.733249e-007, 8.983243e-007, 1.55348e-006, 
    2.445562e-006, 2.904269e-006, 2.690437e-006, 1.812262e-006, 
    1.213482e-006, 9.348323e-007, 4.152789e-007, 1.967287e-007, 8.81987e-008, 
    2.307543e-007, 6.934351e-007, 9.926994e-007, 1.222674e-006, 
    1.273338e-006, 1.047338e-006, 5.220718e-007, 2.553406e-007, 
    3.705763e-007, 4.041035e-007, 5.680172e-007, 7.170283e-007, 
    8.787056e-007, 1.021756e-006, 1.028214e-006, 1.033181e-006, 
    9.241544e-007, 5.650361e-007, 5.123857e-007, 8.228265e-007, 
    1.097505e-006, 1.092786e-006, 9.06273e-007, 8.2829e-007, 8.819345e-007, 
    1.129294e-006, 1.31978e-006, 1.358275e-006, 1.335675e-006, 1.247261e-006, 
    1.096015e-006, 8.464199e-007, 5.918585e-007, 5.329985e-007, 7.49314e-007, 
    1.109674e-006, 1.131777e-006, 7.495621e-007, 7.187662e-007, 
    1.062735e-006, 1.186167e-006, 1.170272e-006, 1.098001e-006, 
    9.181931e-007, 8.970831e-007, 7.992332e-007, 7.979913e-007, 
    6.492282e-007, 4.473172e-007, 4.530295e-007, 4.902824e-007, 
    5.210775e-007, 5.496383e-007, 5.233132e-007, 7.473268e-007, 
    1.080617e-006, 1.39975e-006, 1.63345e-006, 1.712177e-006, 1.696779e-006, 
    1.534853e-006, 9.946862e-007, 6.035309e-007, 5.081636e-007, 
    4.716558e-007, 3.914374e-007, 1.51033e-007, -2.003853e-007, 
    -3.645468e-007, -3.339997e-007, -5.435527e-008, 1.24955e-007, 
    -3.225205e-008, -3.913699e-007, -5.850848e-007, -6.938635e-007, 
    -8.153079e-007, -1.176165e-006, -1.615006e-006, -1.939602e-006, 
    -1.781153e-006, -8.987563e-007,
  2.844416e-006, 2.543661e-006, 1.897695e-006, 1.20504e-006, 7.31432e-007, 
    4.572516e-007, 2.528573e-007, 1.751232e-007, 1.27191e-007, 2.111342e-007, 
    4.565054e-007, 5.451679e-007, 5.955831e-007, 7.202561e-007, 
    8.444326e-007, 9.723353e-007, 1.101727e-006, 1.256698e-006, 
    1.174742e-006, 8.97332e-007, 6.90206e-007, 6.931862e-007, 7.940173e-007, 
    8.014681e-007, 7.530393e-007, 9.122332e-007, 1.202557e-006, 
    1.503064e-006, 1.707707e-006, 1.570367e-006, 1.268123e-006, 
    9.805301e-007, 7.691822e-007, 7.105709e-007, 7.552744e-007, 
    8.379759e-007, 9.075145e-007, 9.400489e-007, 9.137234e-007, 8.72745e-007, 
    9.375651e-007, 1.095518e-006, 1.199081e-006, 1.069689e-006, 8.56106e-007, 
    7.582546e-007, 8.409561e-007, 1.123333e-006, 1.422598e-006, 1.59421e-006, 
    1.490647e-006, 1.131281e-006, 8.101604e-007, 7.957558e-007, 
    9.671189e-007, 1.135254e-006, 1.170769e-006, 1.112654e-006, 
    8.928616e-007, 6.114783e-007, 6.149555e-007, 7.436022e-007, 
    8.255581e-007, 1.014803e-006, 1.226399e-006, 1.199081e-006, 
    1.021509e-006, 7.992328e-007, 6.596588e-007, 6.258829e-007, 
    7.885537e-007, 1.028959e-006, 1.01381e-006, 8.215848e-007, 7.81848e-007, 
    9.802823e-007, 1.164311e-006, 1.19312e-006, 1.050317e-006, 8.441843e-007, 
    6.084979e-007, 4.574995e-007, 3.653608e-007, 2.2678e-007, 8.646043e-008, 
    4.597882e-008, 3.579657e-008, -5.926722e-009, 2.064735e-008, 
    1.902722e-007, 4.185085e-007, 5.593247e-007, 9.114879e-007, 
    1.600418e-006, 2.378507e-006, 2.849136e-006,
  9.537071e-007, 1.064969e-006, 1.085086e-006, 9.430287e-007, 7.26217e-007, 
    5.928514e-007, 5.928518e-007, 6.536984e-007, 6.956702e-007, 
    6.946771e-007, 7.065983e-007, 8.287871e-007, 1.058265e-006, 
    1.289232e-006, 1.396769e-006, 1.38758e-006, 1.349085e-006, 1.336916e-006, 
    1.34238e-006, 1.346601e-006, 1.316055e-006, 1.250738e-006, 1.165801e-006, 
    1.104458e-006, 1.076394e-006, 1.077885e-006, 1.107687e-006, 
    1.147423e-006, 1.163318e-006, 1.136496e-006, 1.082106e-006, 
    1.047089e-006, 1.029456e-006, 1.053546e-006, 1.100485e-006, 
    1.151149e-006, 1.182689e-006, 1.198584e-006, 1.177226e-006, 
    1.100981e-006, 9.604137e-007, 8.054417e-007, 6.688479e-007, 
    5.863947e-007, 5.531153e-007, 5.752188e-007, 6.387968e-007, 
    7.289489e-007, 8.136371e-007, 8.551121e-007, 8.444331e-007, 
    8.002262e-007, 7.530391e-007, 7.585029e-007, 7.788678e-007, 7.64215e-007, 
    7.761359e-007, 8.258064e-007, 9.268863e-007, 1.068696e-006, 1.21572e-006, 
    1.343125e-006, 1.422846e-006, 1.457119e-006, 1.459603e-006, 
    1.407945e-006, 1.263156e-006, 1.067206e-006, 8.836732e-007, 
    8.084219e-007, 8.014681e-007, 8.054417e-007, 7.711687e-007, 
    7.272104e-007, 7.14296e-007, 7.408701e-007, 7.974945e-007, 9.022995e-007, 
    1.017286e-006, 1.081858e-006, 1.061245e-006, 1.00015e-006, 9.740731e-007, 
    9.902162e-007, 1.018032e-006, 9.840073e-007, 8.8715e-007, 7.907893e-007, 
    7.493143e-007, 7.798612e-007, 8.484071e-007, 9.090049e-007, 
    9.144683e-007, 8.968345e-007, 8.819334e-007, 9.018013e-007,
  1.173251e-006, 1.122339e-006, 1.090053e-006, 1.086328e-006, 1.109425e-006, 
    1.161332e-006, 1.225654e-006, 1.287494e-006, 1.342132e-006, 
    1.371686e-006, 1.367464e-006, 1.333688e-006, 1.276815e-006, 1.20678e-006, 
    1.128052e-006, 1.049076e-006, 9.76805e-007, 9.117366e-007, 8.561058e-007, 
    8.138857e-007, 7.820965e-007, 7.575095e-007, 7.341646e-007, 
    7.130545e-007, 6.907028e-007, 6.708347e-007, 6.529533e-007, 
    6.348237e-007, 6.221578e-007, 6.201708e-007, 6.37059e-007, 6.676064e-007, 
    7.051076e-007, 7.485692e-007, 7.93769e-007, 8.399627e-007, 8.856596e-007, 
    9.323501e-007, 9.740734e-007, 1.012568e-006, 1.051559e-006, 1.10123e-006, 
    1.158103e-006, 1.22193e-006, 1.284763e-006, 1.346602e-006, 1.398508e-006, 
    1.439238e-006, 1.470531e-006, 1.492882e-006, 1.507535e-006, 
    1.520201e-006, 1.527403e-006, 1.53088e-006, 1.531376e-006, 1.517717e-006, 
    1.488163e-006, 1.447185e-006, 1.397763e-006, 1.342877e-006, 
    1.288736e-006, 1.235837e-006, 1.185918e-006, 1.14792e-006, 1.11936e-006, 
    1.100484e-006, 1.087819e-006, 1.089309e-006, 1.103962e-006, 
    1.128548e-006, 1.155867e-006, 1.179958e-006, 1.203054e-006, 
    1.221929e-006, 1.245522e-006, 1.271351e-006, 1.302147e-006, 
    1.334433e-006, 1.36647e-006, 1.395527e-006, 1.416886e-006, 1.426323e-006, 
    1.429552e-006, 1.439734e-006, 1.455629e-006, 1.47202e-006, 1.479471e-006, 
    1.481458e-006, 1.484189e-006, 1.482451e-006, 1.476987e-006, 
    1.458857e-006, 1.421356e-006, 1.367463e-006, 1.302395e-006, 1.235588e-006,
  5.48861e-007, 5.143397e-007, 4.984452e-007, 4.994386e-007, 5.15457e-007, 
    5.437696e-007, 5.722059e-007, 6.016355e-007, 6.284577e-007, 
    6.494436e-007, 6.690632e-007, 6.837161e-007, 6.945193e-007, 
    7.032118e-007, 7.084273e-007, 7.177402e-007, 7.263084e-007, 
    7.265569e-007, 7.150084e-007, 6.925325e-007, 6.542864e-007, 6.03374e-007, 
    5.451354e-007, 4.783285e-007, 4.051885e-007, 3.28075e-007, 2.509616e-007, 
    1.768283e-007, 1.08904e-007, 4.706408e-008, -1.179524e-008, 
    -6.941309e-008, -1.312528e-007, -1.932169e-007, -2.607687e-007, 
    -3.275757e-007, -3.938862e-007, -4.567196e-007, -5.173174e-007, 
    -5.703409e-007, -6.124369e-007, -6.390103e-007, -6.551531e-007, 
    -6.624796e-007, -6.557743e-007, -6.300695e-007, -5.794063e-007, 
    -5.015468e-007, -3.989767e-007, -2.765391e-007, -1.392004e-007, 
    3.601599e-009, 1.393269e-007, 2.663592e-007, 3.771252e-007, 
    4.616891e-007, 5.148363e-007, 5.354495e-007, 5.229081e-007, 
    4.912431e-007, 4.48154e-007, 3.963723e-007, 3.345326e-007, 2.68843e-007, 
    1.994281e-007, 1.395751e-007, 1.08656e-007, 1.067924e-007, 1.342355e-007, 
    1.930953e-007, 2.682214e-007, 3.52165e-007, 4.408271e-007, 5.380577e-007, 
    6.336729e-007, 7.156293e-007, 7.739923e-007, 8.056572e-007, 
    8.123627e-007, 8.06278e-007, 7.923704e-007, 7.77221e-007, 7.650519e-007, 
    7.577255e-007, 7.542485e-007, 7.628166e-007, 7.770971e-007, 
    7.955991e-007, 8.105005e-007, 8.116178e-007, 8.016839e-007, 7.78587e-007, 
    7.46674e-007, 7.060682e-007, 6.519274e-007, 5.979107e-007,
  4.332519e-007, 5.07883e-007, 5.29986e-007, 5.071374e-007, 4.917397e-007, 
    5.085035e-007, 5.640104e-007, 6.419932e-007, 7.086755e-007, 
    7.317723e-007, 7.127736e-007, 6.586329e-007, 6.049886e-007, 
    5.705919e-007, 5.566842e-007, 5.343323e-007, 5.008048e-007, 
    4.980729e-007, 5.365675e-007, 5.905842e-007, 6.203867e-007, 
    6.188965e-007, 5.873557e-007, 5.035366e-007, 3.798569e-007, 
    2.636277e-007, 1.774495e-007, 1.315042e-007, 1.126294e-007, 
    1.164789e-007, 1.308833e-007, 1.229359e-007, 1.183415e-007, 
    1.341119e-007, 1.529867e-007, 1.825407e-007, 2.122189e-007, 
    2.107287e-007, 1.745932e-007, 8.344773e-008, -6.283176e-008, 
    -2.45868e-007, -4.606929e-007, -7.489061e-007, -1.115102e-006, 
    -1.548354e-006, -1.983716e-006, -2.385301e-006, -2.762176e-006, 
    -3.154201e-006, -3.487118e-006, -3.683192e-006, -3.627188e-006, 
    -3.273658e-006, -2.680466e-006, -1.895052e-006, -1.096225e-006, 
    -5.065122e-007, -2.061288e-007, -1.829076e-007, -3.753812e-007, 
    -6.82222e-007, -9.637297e-007, -1.084926e-006, -1.028799e-006, 
    -7.772169e-007, -4.157405e-007, -1.241597e-008, 3.520413e-007, 
    5.933152e-007, 6.747759e-007, 6.421171e-007, 5.189343e-007, 
    3.568839e-007, 2.144538e-007, 1.924743e-007, 3.576292e-007, 
    6.506853e-007, 9.042537e-007, 1.077852e-006, 1.200413e-006, 
    1.306335e-006, 1.432871e-006, 1.538049e-006, 1.530722e-006, 
    1.404435e-006, 1.176447e-006, 9.092196e-007, 7.054468e-007, 5.78787e-007, 
    4.875174e-007, 4.233179e-007, 3.643345e-007, 3.228588e-007, 
    3.085788e-007, 3.421064e-007,
  6.746513e-007, 5.508477e-007, 4.312658e-007, 3.639623e-007, 3.851965e-007, 
    4.702572e-007, 6.386404e-007, 7.646788e-007, 7.43569e-007, 6.711746e-007, 
    6.258502e-007, 6.070998e-007, 5.904601e-007, 5.956755e-007, 6.58012e-007, 
    7.287925e-007, 7.839269e-007, 8.40427e-007, 8.55204e-007, 8.29127e-007, 
    7.703917e-007, 6.753966e-007, 5.864865e-007, 6.416208e-007, 
    7.624442e-007, 7.831817e-007, 6.874417e-007, 5.758072e-007, 4.78577e-007, 
    3.863141e-007, 3.51669e-007, 3.885493e-007, 4.020845e-007, 3.829613e-007, 
    3.891702e-007, 4.619375e-007, 5.710879e-007, 5.980344e-007, 
    3.365187e-007, -7.909921e-008, -2.738079e-007, -2.831202e-007, 
    -2.056349e-007, -1.688782e-007, -7.92229e-008, -1.734716e-007, 
    -5.591619e-007, -9.087198e-007, -1.111002e-006, -1.33601e-006, 
    -1.603238e-006, -1.496074e-006, -8.476245e-007, -3.129217e-007, 
    -5.252332e-008, 2.939287e-007, 5.23034e-007, 5.113625e-007, 
    5.117345e-007, 4.762196e-007, 2.512124e-007, 1.505059e-007, 
    4.323847e-007, 1.036255e-006, 1.742693e-006, 1.83806e-006, 1.707177e-006, 
    1.628698e-006, 1.417847e-006, 1.078969e-006, 7.469212e-007, 
    6.439795e-007, 8.435309e-007, 1.078969e-006, 1.213204e-006, 1.31329e-006, 
    1.393881e-006, 1.348059e-006, 1.370659e-006, 1.52948e-006, 1.720216e-006, 
    1.552702e-006, 1.126529e-006, 7.752337e-007, 8.101279e-007, 
    1.170115e-006, 1.584741e-006, 1.592813e-006, 1.068664e-006, 
    6.077216e-007, 4.788253e-007, 6.067276e-007, 7.499025e-007, 
    7.991994e-007, 7.960948e-007, 7.546212e-007,
  2.351912e-007, 1.805533e-007, 2.733136e-007, 6.772593e-007, 1.110883e-006, 
    1.270077e-006, 1.202774e-006, 1.203394e-006, 1.131993e-006, 
    1.048049e-006, 1.164279e-006, 1.217054e-006, 1.27107e-006, 1.37364e-006, 
    1.405553e-006, 1.326329e-006, 1.037867e-006, 7.553656e-007, 
    6.813566e-007, 8.631509e-007, 1.140809e-006, 1.121686e-006, 
    8.635238e-007, 7.01722e-007, 7.369881e-007, 7.784627e-007, 7.854167e-007, 
    6.539137e-007, 6.069753e-007, 6.817297e-007, 6.900493e-007, 6.91912e-007, 
    7.074342e-007, 7.092967e-007, 6.66456e-007, 5.738204e-007, 4.282856e-007, 
    3.733995e-007, 4.856547e-007, 6.298237e-007, 7.326419e-007, 
    1.050657e-006, 1.630312e-006, 2.131737e-006, 1.942867e-006, 
    1.066308e-006, -2.160323e-008, -9.314435e-007, -3.851919e-007, 
    9.844744e-007, 6.591317e-007, -6.175469e-010, 5.935908e-008, 
    4.075491e-007, 7.012277e-007, 5.447655e-007, 2.319648e-007, 
    9.190335e-007, 2.255294e-006, 2.805642e-006, 2.516186e-006, 
    2.072258e-006, 2.577779e-006, 3.571809e-006, 4.559261e-006, 
    4.800784e-006, 4.205111e-006, 3.179041e-006, 2.121929e-006, 
    1.458702e-006, 9.546702e-007, 1.374511e-006, 2.60572e-006, 3.825505e-006, 
    4.180648e-006, 4.161525e-006, 4.146002e-006, 4.172452e-006, 
    4.171459e-006, 3.789742e-006, 2.912312e-006, 1.834585e-006, 
    1.503903e-006, 2.189107e-006, 2.701336e-006, 2.767398e-006, 
    2.546364e-006, 2.001851e-006, 1.626838e-006, 1.356133e-006, 
    1.017007e-006, 6.662094e-007, 6.095843e-007, 7.600847e-007, 
    6.510577e-007, 3.635901e-007,
  2.276654e-006, 1.899775e-006, 1.816577e-006, 2.137449e-006, 2.329922e-006, 
    2.143781e-006, 2.684073e-006, 3.538406e-006, 3.771113e-006, 
    3.937757e-006, 4.101422e-006, 3.960481e-006, 3.228958e-006, 
    2.552942e-006, 2.009299e-006, 1.407043e-006, 6.83468e-007, 3.391269e-007, 
    4.784526e-007, 7.774695e-007, 1.04805e-006, 1.636272e-006, 2.324582e-006, 
    2.060086e-006, 1.443303e-006, 1.067049e-006, 8.093821e-007, 
    8.637719e-007, 1.143665e-006, 1.040102e-006, 6.922844e-007, 
    7.056954e-007, 7.474187e-007, 5.888455e-007, 6.180269e-007, 
    7.425756e-007, 5.198033e-007, 1.610581e-007, -1.989295e-007, 
    -6.874393e-007, -1.247349e-006, -1.363827e-006, -3.700438e-007, 
    1.002106e-006, 1.357002e-006, 9.492087e-007, 4.726207e-007, 
    9.574251e-008, -2.484776e-007, 1.129509e-006, 2.702451e-006, 
    3.17681e-006, 3.802033e-006, 5.385904e-006, 5.75682e-006, 3.919258e-006, 
    2.345943e-006, 2.399713e-006, 2.697981e-006, 2.644458e-006, 
    2.627818e-006, 1.964096e-006, 1.594173e-006, 2.478564e-006, 2.93367e-006, 
    2.569337e-006, 2.821786e-006, 3.949679e-006, 4.625819e-006, 
    5.392236e-006, 5.979961e-006, 6.606432e-006, 7.096184e-006, 
    6.483125e-006, 5.054479e-006, 4.513069e-006, 4.096707e-006, 
    2.647443e-006, 2.095727e-006, 2.309063e-006, 2.670665e-006, 
    3.416096e-006, 2.839667e-006, 2.04494e-006, 1.604114e-006, 2.111871e-006, 
    2.933545e-006, 2.716112e-006, 1.454729e-006, 1.161674e-006, 
    1.899157e-006, 2.893438e-006, 4.199026e-006, 4.639853e-006, 
    4.010776e-006, 3.123536e-006,
  6.174174e-006, 5.372865e-006, 6.407008e-006, 8.038556e-006, 8.416178e-006, 
    7.857383e-006, 7.659074e-006, 7.565944e-006, 7.3274e-006, 7.022299e-006, 
    7.121017e-006, 8.948893e-006, 1.068736e-005, 1.060516e-005, 
    9.375807e-006, 7.503362e-006, 5.913282e-006, 5.143636e-006, 3.8825e-006, 
    3.072498e-006, 3.272298e-006, 3.379216e-006, 3.919011e-006, 5.08639e-006, 
    5.504741e-006, 3.640856e-006, 1.992786e-006, 2.626333e-006, 
    3.064179e-006, 1.563756e-006, 7.207218e-007, 1.67154e-006, 2.801421e-006, 
    3.816314e-006, 5.254773e-006, 6.367394e-006, 6.130838e-006, 
    4.287809e-006, 3.66072e-006, 4.329659e-006, 4.613772e-006, 3.515808e-006, 
    3.744044e-006, 5.570802e-006, 6.246446e-006, 6.475919e-006, 
    5.384905e-006, 4.192067e-006, 2.893306e-006, 1.275044e-006, 
    1.240898e-006, 1.946839e-006, 2.599008e-006, 3.45359e-006, 2.906971e-006, 
    2.248587e-006, 1.341976e-006, 6.511837e-007, 3.524146e-007, 
    2.162784e-006, 3.287199e-006, 3.625208e-006, 4.69449e-006, 6.418307e-006, 
    6.791207e-006, 4.232306e-006, 2.969184e-006, 2.772862e-006, 
    3.303592e-006, 4.921734e-006, 6.34293e-006, 6.638344e-006, 6.352489e-006, 
    5.565959e-006, 6.301952e-006, 7.393213e-006, 7.011496e-006, 
    5.607435e-006, 4.278498e-006, 5.003814e-006, 6.326663e-006, 
    6.415572e-006, 5.274022e-006, 3.039841e-006, 2.839544e-006, 
    2.881143e-006, 3.252679e-006, 3.699713e-006, 2.865371e-006, 
    2.117209e-006, 1.677625e-006, 3.000723e-006, 4.018844e-006, 
    4.856787e-006, 5.814434e-006, 6.38577e-006,
  6.254639e-006, 7.718429e-006, 1.050395e-005, 1.153809e-005, 1.050792e-005, 
    8.261195e-006, 7.607907e-006, 6.975975e-006, 5.673241e-006, 
    5.083404e-006, 4.813317e-006, 5.309399e-006, 7.805716e-006, 
    8.213265e-006, 7.460265e-006, 7.860726e-006, 1.140609e-005, 
    1.319832e-005, 1.233207e-005, 9.767333e-006, 7.947532e-006, 8.36961e-006, 
    7.60245e-006, 7.046012e-006, 6.948161e-006, 5.315242e-006, 3.227216e-006, 
    1.658249e-006, 1.040968e-006, 1.71922e-006, 2.139059e-006, 2.652776e-006, 
    3.425403e-006, 3.661213e-006, 4.929669e-006, 6.065758e-006, 
    7.830926e-006, 9.550522e-006, 9.787325e-006, 1.123721e-005, 
    1.140448e-005, 1.073293e-005, 7.642306e-006, 2.837922e-006, 
    3.319725e-006, 3.692998e-006, 2.518043e-006, 2.71114e-006, 3.3504e-006, 
    3.482772e-006, 3.548705e-006, 3.475197e-006, 4.546715e-006, 
    4.555655e-006, 3.678351e-006, 3.526606e-006, 4.207341e-006, 
    4.036721e-006, 3.799918e-006, 4.851316e-006, 4.22411e-006, 1.92896e-006, 
    3.652522e-006, 4.329035e-006, 3.727151e-006, 3.556162e-006, 
    3.364432e-006, 3.053741e-006, 4.428375e-006, 6.590781e-006, 
    7.446728e-006, 6.944192e-006, 6.755314e-006, 6.182863e-006, 
    5.530066e-006, 6.210304e-006, 6.527327e-006, 7.286539e-006, 
    6.078302e-006, 4.60533e-006, 5.017719e-006, 5.675234e-006, 5.296e-006, 
    5.422289e-006, 4.689771e-006, 5.299726e-006, 6.056827e-006, 
    4.850826e-006, 3.875048e-006, 4.433967e-006, 6.235892e-006, 
    8.254872e-006, 8.322424e-006, 5.701686e-006, 5.247943e-006, 5.576512e-006,
  7.247676e-006, 6.861113e-006, 5.913897e-006, 5.377578e-006, 5.83827e-006, 
    5.928916e-006, 5.869932e-006, 5.072225e-006, 4.72478e-006, 5.087621e-006, 
    4.404901e-006, 3.519399e-006, 3.861751e-006, 5.824855e-006, 
    6.254137e-006, 3.42416e-006, 3.364679e-006, 5.804864e-006, 8.154031e-006, 
    8.732326e-006, 8.817757e-006, 8.723508e-006, 7.458402e-006, 
    6.900724e-006, 5.965801e-006, 5.793318e-006, 5.815797e-006, 
    5.529444e-006, 2.871948e-006, 9.819832e-007, 1.20922e-006, 2.23206e-006, 
    1.091757e-006, 4.149915e-007, 2.051511e-006, 5.499765e-006, 
    6.963433e-006, 5.884591e-006, 5.301954e-006, 5.294005e-006, 
    7.766979e-006, 6.956356e-006, 4.176167e-006, 3.786499e-006, 
    5.556012e-006, 6.553153e-006, 4.402787e-006, 2.606579e-006, 
    3.684305e-006, 4.891797e-006, 7.13231e-006, 7.960318e-006, 6.862849e-006, 
    6.062406e-006, 4.122279e-006, 3.958863e-006, 3.486244e-006, 
    4.111225e-006, 6.835158e-006, 6.31995e-006, 4.756941e-006, 4.397703e-006, 
    3.983694e-006, 3.298614e-006, 4.522748e-006, 6.173175e-006, 
    6.150078e-006, 7.543336e-006, 8.634719e-006, 8.568286e-006, 
    6.122884e-006, 3.867595e-006, 2.512583e-006, 3.462525e-006, 
    5.871176e-006, 6.385266e-006, 6.6135e-006, 5.746257e-006, 5.646671e-006, 
    4.930916e-006, 4.823629e-006, 5.157166e-006, 5.378821e-006, 
    5.513431e-006, 6.733961e-006, 6.307786e-006, 3.882247e-006, 3.25466e-006, 
    4.563479e-006, 4.431482e-006, 3.981468e-006, 3.840647e-006, 
    4.402669e-006, 4.983567e-006, 5.395214e-006, 6.084514e-006,
  3.956624e-006, 4.147487e-006, 4.967667e-006, 3.178659e-006, 3.783771e-006, 
    5.523234e-006, 5.118916e-006, 2.905344e-006, 2.156685e-006, 
    2.880392e-006, 4.497913e-006, 5.324928e-006, 6.862105e-006, 
    8.442996e-006, 7.712835e-006, 4.755329e-006, 4.098063e-006, 5.90098e-006, 
    5.572285e-006, 5.521864e-006, 5.974121e-006, 4.73695e-006, 4.810714e-006, 
    5.30059e-006, 5.70478e-006, 4.985675e-006, 4.817295e-006, 5.102025e-006, 
    3.666177e-006, 3.558762e-006, 6.053844e-006, 5.728873e-006, 
    4.023554e-006, 3.547095e-006, 5.975733e-006, 6.826096e-006, 4.83865e-006, 
    3.122281e-006, 5.165606e-006, 8.871524e-006, 1.05114e-005, 8.779636e-006, 
    8.521223e-006, 9.385614e-006, 6.275124e-006, 4.217276e-006, 
    6.914132e-006, 5.858135e-006, 5.202983e-006, 6.592396e-006, 
    6.820999e-006, 5.71509e-006, 3.113964e-006, 5.494923e-006, 6.071103e-006, 
    6.019067e-006, 5.986907e-006, 6.72414e-006, 7.607281e-006, 5.633499e-006, 
    6.592638e-006, 7.883209e-006, 7.744498e-006, 5.56831e-006, 5.861737e-006, 
    5.743397e-006, 5.957105e-006, 6.503107e-006, 1.035643e-005, 
    1.154119e-005, 9.8442e-006, 7.589031e-006, 7.624547e-006, 7.759032e-006, 
    6.95623e-006, 6.586681e-006, 5.914142e-006, 4.231679e-006, 2.382563e-006, 
    1.594046e-006, 2.540517e-006, 2.44826e-006, 2.355251e-006, 2.719835e-006, 
    9.160485e-007, 8.205516e-007, 1.647693e-006, 1.815331e-006, 
    2.415971e-006, 1.024451e-006, 9.321884e-007, 1.587096e-006, 
    2.818055e-006, 4.136435e-006, 4.268311e-006, 3.943338e-006,
  7.244191e-006, 8.865441e-006, 7.195642e-006, 6.000937e-006, 3.79917e-006, 
    4.745147e-006, 4.864476e-006, 5.140642e-006, 3.608562e-006, 
    1.857425e-006, 4.634505e-006, 6.332615e-006, 8.153416e-006, 
    7.509931e-006, 5.111833e-006, 5.123136e-006, 5.532176e-006, 
    5.276743e-006, 1.869219e-006, 1.19122e-006, 2.082557e-006, 3.13334e-006, 
    4.093967e-006, 4.623576e-006, 4.764395e-006, 3.098816e-006, 
    3.346544e-006, 4.739682e-006, 3.898756e-006, 4.749862e-006, 
    4.043297e-006, 4.373236e-006, 2.927696e-006, 3.349898e-006, 
    3.876532e-006, 3.967929e-006, 3.951161e-006, 5.704038e-006, 
    7.499504e-006, 6.587175e-006, 3.50723e-006, 2.304831e-006, 7.331328e-007, 
    1.889584e-006, 2.034001e-006, 1.787143e-006, 2.046174e-006, 
    5.153564e-006, 4.726397e-006, 2.932666e-006, 1.093988e-006, 
    1.056862e-006, 1.321732e-006, 8.784191e-007, 2.097335e-006, 
    3.085031e-006, 2.530458e-006, 3.555535e-006, 3.8666e-006, 2.939378e-006, 
    3.806497e-006, 5.143753e-006, 3.671394e-006, 4.781898e-006, 
    6.134433e-006, 7.388364e-006, 7.38079e-006, 1.023486e-005, 9.889398e-006, 
    6.934748e-006, 4.553047e-006, 4.077949e-006, 3.392619e-006, 
    4.108613e-006, 2.691762e-006, 2.262117e-006, 2.067402e-006, 4.29116e-006, 
    3.853562e-006, 2.337867e-006, -1.118842e-007, -4.836729e-007, 
    5.178135e-007, 6.869377e-007, -6.593837e-008, -1.516273e-007, 
    1.335757e-006, 2.080447e-006, 2.069144e-006, 2.309051e-006, 
    2.783781e-006, 3.45545e-006, 4.071364e-006, 5.126116e-006, 5.034479e-006, 
    5.125617e-006,
  4.11272e-006, 3.002955e-006, 2.904981e-006, 3.681082e-006, 5.161015e-006, 
    3.823883e-006, 2.906461e-006, 3.389636e-006, 3.295267e-006, 
    4.955127e-006, 4.974376e-006, 6.034596e-006, 6.561349e-006, 
    5.471953e-006, 5.563466e-006, 4.861624e-006, 4.008161e-006, 3.79793e-006, 
    9.704345e-007, 7.701383e-007, 3.184374e-006, 3.791472e-006, 1.14453e-006, 
    -2.333898e-006, -3.515313e-006, -7.123999e-007, 1.488002e-006, 
    3.248202e-006, 5.893275e-006, 5.729988e-006, 3.48339e-006, 1.393131e-006, 
    8.989082e-007, 2.913293e-006, 2.384179e-006, 3.617206e-007, 
    1.664706e-006, 1.514451e-006, -8.431634e-007, -2.019151e-007, 
    1.177559e-006, 2.685436e-006, 2.185479e-007, -3.676127e-006, -2.883e-006, 
    -7.649251e-007, 2.516928e-006, 4.387268e-006, 6.94632e-007, 
    -1.045664e-007, -1.543642e-006, -1.921133e-006, 9.324394e-007, 
    1.327564e-006, 1.374257e-006, 2.69611e-006, 4.904341e-006, 7.304545e-006, 
    4.252666e-006, 1.688542e-006, 5.212551e-006, 7.274739e-006, 
    4.145004e-006, 4.702182e-006, 4.725654e-006, 7.8544e-006, 9.922183e-006, 
    9.992465e-006, 8.162977e-006, 4.466863e-006, 3.274523e-006, 
    3.931382e-007, -7.143935e-007, -4.681497e-007, 2.524466e-007, 
    -1.97726e-006, -2.224744e-006, 1.123735e-007, 2.720946e-006, 
    2.61987e-006, -7.003837e-008, -1.746417e-006, -1.315899e-006, 
    -1.960376e-006, -5.173279e-007, -1.004348e-006, -1.762441e-006, 
    -1.360106e-006, 1.959619e-006, 3.319972e-006, 2.158558e-006, 
    3.703553e-006, 3.28707e-006, 1.673772e-006, 1.07276e-006, 1.459321e-006,
  1.21817e-006, -1.267344e-006, 1.387914e-006, 2.042198e-006, 1.607208e-006, 
    2.985067e-006, 2.475448e-006, 3.040082e-006, 1.306829e-006, 1.33924e-006, 
    1.709906e-006, 2.246839e-006, 6.912815e-007, 6.033661e-007, 
    1.133973e-006, 1.15285e-006, -1.718974e-006, -1.407421e-006, 
    1.072625e-006, 2.684937e-006, 3.519897e-006, 2.877288e-006, 
    1.772609e-006, 6.77006e-007, 6.64957e-007, 1.196808e-006, 3.28806e-006, 
    1.908087e-006, 1.211709e-006, -2.444292e-006, -3.00433e-006, 
    -1.000622e-006, -3.281242e-006, -4.14054e-006, -3.208104e-006, 
    -2.90772e-006, -2.281129e-006, -1.948392e-007, 1.286211e-006, 
    -1.072764e-006, -1.819186e-006, -2.381454e-006, -2.683701e-006, 
    -2.225366e-006, 1.869346e-006, 3.089503e-006, 7.862764e-007, 
    -2.281617e-006, -4.544487e-006, -2.750759e-006, -4.218029e-006, 
    -2.084424e-006, 1.462173e-006, 1.069777e-006, 1.005901e-008, 
    -1.416229e-006, 6.972514e-007, 4.742782e-006, 5.473441e-006, 
    3.319852e-006, 1.234308e-006, 1.476325e-006, 3.242116e-006, 4.46277e-006, 
    6.771206e-006, 8.55239e-006, 7.913884e-006, 4.298116e-006, 1.16204e-006, 
    -3.558027e-006, -4.207344e-006, -6.346658e-006, -4.136687e-006, 
    -5.945585e-007, -2.654273e-006, -4.174308e-006, -8.376188e-006, 
    -7.236005e-006, -2.236167e-006, 1.612558e-006, 5.708425e-007, 
    1.30236e-006, 2.76615e-006, 4.549765e-007, -2.194203e-006, 
    -1.901022e-006, -1.282864e-006, 1.672408e-006, 2.657747e-006, 
    7.494091e-007, -3.873029e-007, -3.312405e-006, -6.521124e-006, 
    -6.197522e-006, -2.571818e-006, 6.246082e-007,
  1.407407e-006, 9.983705e-007, -2.032277e-006, -6.549126e-007, 
    -7.92872e-007, -8.543429e-008, 1.474225e-006, 2.573433e-006, 
    2.175202e-006, 1.393504e-006, 1.897406e-007, 2.132092e-007, 
    -5.935908e-008, -4.970789e-007, -2.371962e-008, 2.072502e-006, 
    4.139536e-006, 3.789484e-006, 2.235416e-006, 4.263587e-006, 
    2.073859e-006, 6.653318e-007, -2.521159e-006, -3.688663e-006, 
    -2.538414e-006, -3.20015e-006, -2.153347e-006, -4.20809e-006, 
    -4.090247e-006, -2.154709e-006, -2.982717e-006, -2.942608e-006, 
    -3.665315e-006, -3.739324e-006, -1.814591e-006, 1.208731e-006, 
    2.942481e-006, 2.498798e-006, -1.183651e-006, -1.000242e-006, 
    5.250149e-007, 2.103297e-006, 2.728524e-006, 2.844879e-006, 
    -2.379311e-007, 5.134643e-007, -8.054158e-007, -7.632003e-006, 
    -7.009879e-006, -6.091221e-006, -2.892812e-006, -6.43231e-008, 
    4.387148e-007, 4.564681e-007, -5.877264e-007, 3.442165e-006, 
    4.032248e-006, 1.626951e-006, 6.93024e-007, 3.829628e-007, 
    -2.123852e-008, 2.289315e-006, 1.518922e-006, -6.899281e-007, 
    -2.320859e-006, -8.694769e-010, -1.489127e-006, 1.784392e-007, 
    -3.917514e-006, -5.967922e-007, -2.32958e-007, 6.422379e-007, 
    6.537848e-007, -5.36094e-006, -6.830694e-006, -8.362038e-006, 
    -1.20343e-005, -1.168898e-005, -3.748009e-006, 3.034998e-006, 
    7.628776e-006, 6.001937e-006, 7.005965e-007, 2.981596e-006, 
    2.134584e-006, 2.567966e-006, 2.126762e-006, 5.129095e-006, 
    2.299985e-006, -3.012145e-006, -3.609559e-006, -3.700206e-006, 
    -2.597521e-006, 3.966161e-007, 9.519317e-007, 8.488641e-007,
  -2.110755e-006, -3.262363e-006, -2.212075e-006, -2.449871e-006, 
    -2.479053e-006, -1.713506e-006, -1.580889e-006, 3.133593e-006, 
    6.610157e-006, 6.180504e-006, 4.740978e-007, -1.913313e-006, 
    -1.987446e-006, -5.194919e-006, -2.769011e-006, -2.786528e-007, 
    1.4464e-006, 3.848098e-006, 2.714121e-006, -1.040602e-006, -1.38581e-006, 
    -1.147515e-006, -1.306462e-006, 2.26932e-006, 1.080331e-006, 
    7.798008e-008, -1.996508e-006, -2.651788e-006, -2.673891e-006, 
    -3.299614e-006, -3.430747e-006, -3.39424e-006, -4.119926e-006, 
    -1.40394e-006, 1.607212e-006, 2.093737e-006, 1.877668e-006, 
    7.985818e-007, 9.470969e-007, 2.540404e-006, 4.733607e-006, 
    6.979579e-006, 8.566551e-006, 6.444128e-006, 3.176798e-006, 
    2.614033e-006, -2.398712e-006, -5.303948e-006, -3.274781e-006, 
    -4.296384e-006, -2.357734e-006, 9.200157e-007, 2.140801e-006, 
    3.375098e-007, 1.337379e-006, 2.950175e-006, -1.695262e-006, 
    7.60705e-007, 3.074725e-006, 8.024217e-007, -9.521827e-007, 
    3.787136e-008, -3.609559e-006, -2.515695e-006, -8.18327e-008, 
    4.944704e-007, 4.567206e-006, -1.458822e-006, -4.16984e-006, 
    -2.894059e-006, -3.356981e-006, -3.996491e-006, -6.940711e-006, 
    -1.008101e-005, -1.066873e-005, -9.064004e-006, -1.151822e-005, 
    -1.195433e-005, -8.067691e-007, 8.320809e-006, 1.241031e-005, 
    1.028465e-005, 1.083823e-005, 5.73694e-006, 6.744758e-006, 3.618494e-006, 
    5.030499e-006, 3.831952e-006, 1.403814e-006, -1.958138e-006, 
    3.375062e-007, 1.643964e-006, 7.573453e-007, 1.156081e-006, 
    1.428272e-006, -1.204899e-008,
  -4.918378e-006, -6.636601e-006, -5.619597e-006, -4.374978e-006, 
    -2.617387e-006, -1.774602e-006, -3.25088e-007, 4.932299e-007, 
    1.670045e-006, -3.099449e-006, -4.497673e-006, -5.250051e-006, 
    -6.913144e-006, -5.519885e-006, -4.552679e-006, 2.41411e-006, 
    1.040188e-005, 4.484125e-006, -1.410148e-006, 3.086398e-006, 
    3.580248e-006, 1.526369e-006, -2.135215e-006, -3.244233e-006, 
    -3.888832e-006, -2.604353e-006, -7.527578e-007, -1.603988e-006, 
    -2.108758e-006, -3.511705e-006, -5.794316e-006, -5.011383e-006, 
    1.229819e-008, 3.118319e-006, 2.174704e-006, 2.411881e-006, 
    8.442785e-007, 1.878543e-006, 1.850603e-006, 2.392632e-006, 
    5.382427e-006, 1.045242e-005, 8.836509e-006, 4.165246e-006, 
    1.579274e-006, -3.971181e-007, -2.83905e-006, -1.613309e-006, 
    -3.67227e-006, 3.551813e-006, 8.676143e-007, -3.055738e-006, 
    -3.344194e-006, -1.743065e-006, -2.295772e-006, 1.849723e-006, 
    9.05864e-007, 5.693473e-007, 1.036122e-006, -5.911537e-006, 
    -6.636979e-006, -3.348661e-006, -1.718101e-006, 5.815178e-006, 
    6.972747e-006, 1.222637e-006, -3.284465e-006, -5.929665e-006, 
    -7.450584e-006, -7.832798e-006, -1.26116e-005, -1.082334e-005, 
    -1.052419e-005, -9.036812e-006, -3.502885e-006, -5.611651e-006, 
    -6.055458e-006, -5.407256e-006, 1.643227e-006, 1.408072e-005, 
    2.100157e-005, 1.360352e-005, 1.256552e-005, 1.234573e-005, 
    3.953024e-006, 3.782334e-007, -1.906605e-006, -5.465994e-006, 
    -4.08764e-006, -1.784541e-006, 3.553923e-007, -6.057344e-007, 
    -3.791725e-006, -3.775336e-006, -4.150595e-006, -5.274762e-006,
  -4.793825e-006, -3.292037e-006, -3.140046e-006, -2.688168e-006, 
    -1.158564e-006, 5.503503e-007, -6.840837e-007, -1.625465e-006, 
    -3.367677e-007, -5.774076e-006, -7.825965e-006, -4.844245e-006, 
    -3.035118e-006, -3.200776e-006, -4.265461e-006, -1.625223e-006, 
    6.556882e-006, 2.755965e-006, 7.034461e-006, 1.018121e-005, 7.66162e-007, 
    -4.836551e-006, -1.69628e-007, -1.621793e-007, 8.755687e-007, 
    -1.137581e-006, -1.308941e-006, -6.97868e-007, -1.799272e-007, 
    -9.484611e-007, -2.956388e-006, 7.778417e-007, 3.216296e-006, 
    2.677618e-006, 2.296894e-006, -2.292272e-007, -1.657254e-006, 
    2.050526e-006, 3.980102e-006, 7.796788e-006, 1.071455e-005, 
    1.275427e-005, 1.490735e-006, -1.927237e-007, -2.247349e-006, 
    2.713623e-006, 2.777568e-006, 3.513069e-006, -1.731889e-006, 
    5.790353e-007, -2.982968e-006, -4.040739e-007, 6.23129e-006, 
    6.783372e-006, 1.365343e-005, 1.169518e-005, 2.695244e-006, 
    -1.095108e-006, -4.99624e-006, -5.837159e-006, -1.710399e-006, 
    -1.031003e-008, 7.42351e-006, 9.582069e-006, 4.424532e-006, 
    -1.416476e-006, -4.689275e-006, -3.171346e-006, -6.057819e-006, 
    -7.495162e-006, -4.86287e-006, -4.975622e-006, -5.425141e-006, 
    -3.223863e-006, -2.515067e-006, -2.588827e-006, -2.548842e-006, 
    -1.008559e-006, 7.59836e-007, 1.362326e-005, 1.260526e-005, 6.22098e-006, 
    7.687997e-006, 8.138515e-006, 2.801415e-006, -1.48789e-006, 
    -5.846232e-007, -1.517064e-006, -2.571571e-006, -3.054756e-007, 
    -2.011659e-006, -1.078597e-006, -1.373272e-006, -5.852184e-006, 
    -5.528953e-006, -3.951907e-006,
  -1.791987e-006, -1.2132e-006, -1.669301e-006, -3.082041e-007, 
    -1.22028e-006, -1.411138e-006, -1.95441e-006, -5.812653e-007, 
    -3.696861e-006, -8.45964e-006, -7.683289e-006, -5.492569e-006, 
    -7.100156e-006, -1.183139e-005, -1.11257e-005, -4.339097e-006, 
    -3.116333e-006, 1.994267e-006, 8.49316e-006, 6.540984e-006, 
    1.554308e-006, -5.258917e-007, -1.60014e-006, -5.02172e-007, 
    6.305672e-007, -4.984564e-006, -2.211582e-006, 1.176451e-006, 
    2.542018e-006, 8.704956e-008, 4.570191e-006, 1.441443e-006, 3.36841e-006, 
    9.749128e-007, -1.041712e-006, -9.115761e-007, 1.277279e-006, 
    2.785277e-006, 7.284808e-006, 4.502889e-006, 5.401425e-006, 
    -8.591778e-007, 4.277863e-007, 8.15205e-006, 8.922812e-006, 
    8.106228e-006, 7.364521e-006, -3.145433e-007, 3.188798e-007, 
    3.213929e-006, 9.69656e-006, 1.439701e-005, 1.591692e-005, 2.057763e-005, 
    1.222702e-005, 9.970616e-006, -1.855318e-006, 2.955152e-006, 
    -1.875051e-007, -2.327306e-006, 3.503766e-006, 1.994522e-006, 
    2.14887e-006, 2.07809e-006, -1.906355e-006, -4.749876e-006, 
    -7.194405e-006, -8.483607e-006, -7.221599e-006, -2.768014e-006, 
    -2.746653e-006, -2.33538e-006, -2.643465e-006, -1.822658e-006, 
    -1.352278e-006, -1.132238e-006, -5.554391e-007, -3.808475e-007, 
    -6.98491e-007, 1.056405e-005, 6.320819e-006, 4.998074e-007, 
    1.516815e-006, -4.753456e-007, 3.311154e-006, 1.829729e-006, 
    -2.480672e-006, -3.897399e-006, -4.417947e-006, -5.546835e-006, 
    -4.158792e-006, -1.514829e-006, -3.826613e-006, -6.496778e-006, 
    -3.917883e-006, -1.280751e-006,
  -1.018368e-006, -4.435565e-007, -4.996843e-007, -5.750593e-007, 
    -9.767696e-007, -6.058544e-007, 1.230596e-007, -5.935619e-007, 
    -5.962934e-007, -2.046052e-006, -5.374975e-006, -2.626455e-006, 
    -1.325579e-006, -5.060432e-006, -1.821663e-006, 2.612669e-006, 
    -1.189481e-006, -4.051253e-006, -2.002467e-006, 2.739573e-006, 
    1.181903e-006, 5.301627e-008, 2.359229e-008, -6.220016e-007, 
    -2.22288e-006, -4.126256e-006, -2.538036e-006, 4.867743e-007, 
    7.55861e-007, 5.833801e-006, 8.086237e-006, 3.236536e-006, 1.362589e-006, 
    1.806146e-006, 1.316767e-006, 1.238536e-006, 1.233817e-006, 
    1.556676e-006, 2.184388e-006, 2.386299e-006, 5.648038e-006, 
    3.889574e-006, 1.055064e-005, 1.243651e-005, 9.153278e-006, 
    7.650127e-006, 5.915015e-006, 1.379996e-005, 1.0121e-005, 1.098737e-005, 
    1.956038e-005, 2.37727e-005, 1.733328e-005, 2.170615e-005, 8.949646e-006, 
    2.30869e-006, -2.552693e-006, -3.723177e-006, -6.141021e-006, 
    -3.745532e-006, -1.06691e-005, -1.269554e-005, -1.444009e-005, 
    -1.274223e-005, -1.10517e-005, -1.082097e-005, -9.727353e-006, 
    -7.158269e-006, -1.480179e-006, 4.568492e-007, -1.264608e-006, 
    -2.431343e-007, -4.785725e-007, 4.034528e-007, -2.279864e-007, 
    -4.132578e-007, 2.486028e-007, 8.965662e-008, -5.101156e-007, 
    4.301593e-006, 2.705801e-006, 7.679046e-007, -7.760982e-007, 
    -1.917155e-006, -1.041715e-006, -3.163768e-006, -5.852307e-006, 
    -4.838661e-006, -3.259134e-006, -4.71535e-006, -4.465257e-006, 
    -4.104397e-006, -6.781514e-006, -2.919011e-006, -1.02346e-006, 
    -7.491526e-007,
  -7.097906e-007, -2.974011e-007, -5.180623e-007, 1.960759e-007, 
    5.565598e-007, 5.432721e-007, -3.247201e-007, -8.165825e-007, 
    5.118559e-007, -4.215754e-007, -1.370909e-006, 1.86115e-006, 
    6.996461e-006, -1.236924e-006, -1.447897e-006, 3.787009e-006, 
    6.82101e-006, 4.015739e-006, -6.22384e-006, -2.685956e-007, 
    6.823466e-007, 1.465403e-006, -1.247976e-006, -2.037985e-006, 
    -2.572315e-006, -6.159171e-007, -6.978717e-007, 4.464015e-006, 
    2.334509e-006, 1.351547e-005, 1.567875e-005, 5.029393e-006, 
    -1.468259e-006, 3.201271e-007, -3.396212e-007, 3.376853e-006, 
    4.934273e-006, -1.045537e-007, -2.057103e-006, 2.809495e-006, 
    5.591535e-006, 8.458766e-006, 1.859031e-005, 1.173975e-005, 
    1.328364e-005, 2.336602e-005, 1.365506e-005, 1.418776e-005, 
    2.426381e-005, 2.369831e-005, 2.541332e-005, 1.888597e-005, 
    1.910378e-005, 1.019922e-005, 1.505898e-006, 6.786111e-006, 2.99501e-006, 
    -3.592795e-006, -6.888062e-006, -8.08388e-006, -1.37113e-005, 
    -1.704941e-005, -1.417485e-005, -1.176447e-005, -1.175503e-005, 
    -8.000557e-006, -4.050877e-006, -6.413675e-007, 1.000617e-006, 
    -6.258051e-008, 3.494351e-007, 1.093122e-008, 4.284448e-008, 
    1.668946e-007, -6.799883e-007, -8.778989e-008, -3.839519e-007, 
    -6.262196e-007, 2.542887e-006, 7.934614e-006, 5.131085e-006, 
    6.633491e-007, -1.811731e-006, -3.79023e-006, -9.936838e-006, 
    -1.125025e-005, -1.097346e-005, -9.99917e-006, -8.151063e-006, 
    -5.158909e-006, -2.901501e-006, -2.947197e-006, -1.034884e-006, 
    6.837181e-007, -8.802826e-007, -1.449107e-007,
  -5.671118e-007, -4.282829e-007, 4.163639e-007, -1.270198e-006, 
    -1.241733e-007, -2.232813e-006, -8.806574e-007, -1.709659e-006, 
    -1.249213e-006, 1.211993e-007, 5.093219e-006, 7.469207e-006, 
    1.594561e-005, -1.744436e-006, 1.979373e-006, 1.879911e-006, 
    9.755291e-006, 1.04451e-005, 3.279372e-006, 1.713334e-005, 5.918369e-006, 
    1.169405e-005, 1.809742e-006, 7.354218e-006, 3.54138e-006, 2.875797e-006, 
    5.04441e-006, 1.520117e-005, 7.699429e-006, 1.035146e-005, 1.400151e-005, 
    1.334436e-005, 3.361829e-006, 1.809997e-006, 2.765446e-007, 
    2.029044e-006, 4.931792e-006, 6.266058e-006, 8.464727e-006, 
    1.640655e-005, 1.033259e-005, 1.534845e-005, 1.485211e-005, 
    6.999311e-006, 2.000356e-005, 3.801472e-005, 2.567781e-005, 
    1.574978e-005, 3.230062e-005, 2.09221e-005, 2.397966e-006, 
    -2.324581e-006, 2.758949e-006, -1.173913e-005, -1.04975e-005, 
    -3.786648e-006, -5.30445e-006, -1.605971e-006, -6.30915e-006, 
    -4.963076e-006, -8.850908e-006, -7.742272e-006, -6.403154e-006, 
    -7.356578e-006, -4.514181e-006, -2.394364e-006, -1.646549e-007, 
    -8.890584e-008, -4.734811e-007, -1.568841e-006, -9.871992e-007, 
    -9.459727e-007, -1.312293e-006, -1.823029e-006, -1.299753e-006, 
    -8.016809e-007, -1.816202e-006, -8.472507e-007, 1.467068e-005, 
    5.685979e-007, 2.380828e-006, -2.25405e-006, -4.689268e-006, 
    -8.283802e-006, -6.026897e-006, -1.176968e-005, -1.533963e-005, 
    -1.448095e-005, -1.107218e-005, -5.124757e-006, -4.22202e-007, 
    1.496373e-007, 6.295886e-008, -9.520572e-007, -7.287881e-007, 
    -6.571381e-007,
  -5.846205e-007, 1.841911e-006, -4.046418e-006, -5.712231e-006, 
    -7.574818e-007, -3.040703e-006, -4.276878e-006, -2.474088e-006, 
    -3.239262e-006, -3.192694e-006, 2.312414e-006, 2.579261e-006, 
    3.706915e-006, -8.641309e-006, 1.645712e-006, 1.551954e-006, 
    1.240943e-005, 1.306148e-005, 9.318304e-006, 2.489027e-005, 
    9.711959e-006, 2.116576e-006, 2.536173e-006, 1.233121e-005, 
    9.373696e-006, 6.462258e-006, 1.177701e-005, 8.859606e-006, 
    -9.618743e-007, -5.809467e-006, -1.943234e-006, 4.305111e-007, 
    6.574766e-006, 6.487098e-006, 5.270907e-006, -3.802406e-006, 
    -7.385268e-006, 6.405142e-006, 1.199122e-005, 6.587426e-006, 
    2.020213e-006, 2.105446e-005, 1.056604e-005, -3.427391e-006, 
    6.978211e-006, 2.558381e-005, 3.734517e-005, 2.502909e-005, 
    2.457549e-005, 1.576617e-005, 1.416731e-006, 8.119969e-007, 
    6.021437e-007, -7.364513e-006, -1.351175e-005, -8.020674e-006, 
    -3.838541e-006, 4.141526e-006, 5.487229e-006, 3.556906e-006, 
    8.57679e-007, -3.430248e-006, -4.401307e-006, -2.460798e-006, 
    -1.750262e-006, -2.329793e-006, -1.267465e-006, -1.885118e-006, 
    -2.60323e-006, -2.456455e-006, -2.760686e-006, -2.373505e-006, 
    -2.453474e-006, -1.632172e-006, -7.851656e-007, 3.69487e-006, 
    2.937268e-006, 1.025214e-005, -2.590066e-006, 7.1264e-007, 8.153402e-007, 
    -6.713719e-006, -6.586686e-006, -6.806227e-006, -1.15099e-005, 
    -1.262054e-005, -2.016525e-005, -1.269926e-005, -7.667637e-006, 
    2.382571e-006, 8.513651e-006, 7.21626e-006, 4.089503e-006, 6.854571e-007, 
    1.245492e-006, 2.525785e-007,
  4.225103e-006, 2.194687e-006, -1.70742e-006, -3.927325e-006, 1.077887e-005, 
    3.656245e-006, 2.517048e-006, 8.477766e-006, 8.191659e-006, 
    3.106517e-006, -1.778457e-006, -4.649904e-006, -2.268207e-006, 
    -2.377608e-006, 5.394962e-006, 7.98727e-006, 1.574419e-005, 
    1.189845e-005, 7.16994e-006, 2.094603e-006, -1.953667e-006, 
    -3.415727e-006, 1.64027e-005, 1.693045e-005, 9.116397e-006, 3.97885e-006, 
    5.910922e-006, 2.44056e-006, 6.200135e-007, -4.153691e-006, 
    -4.717826e-006, -4.725895e-006, -5.716218e-006, -6.842492e-006, 
    -6.026647e-006, -9.760261e-006, -1.214917e-005, 7.856634e-006, 
    1.2628e-005, 7.491326e-006, 1.08473e-005, 4.510963e-006, -2.286717e-006, 
    -7.2283e-006, 1.258751e-005, 2.36803e-005, 3.473286e-005, 1.799937e-005, 
    1.153399e-005, 3.116814e-005, 2.089143e-005, 1.208262e-005, 8.16198e-006, 
    -3.816298e-006, -4.615882e-006, -1.287473e-005, -1.416603e-005, 
    -8.131552e-006, -5.421796e-006, -1.262815e-007, 1.542641e-006, 
    -2.231427e-007, -3.786259e-006, -3.133591e-006, -1.989674e-006, 
    -1.50576e-006, -1.176568e-006, -1.570083e-006, -2.456455e-006, 
    -2.389275e-006, -2.187736e-006, -2.186868e-006, -2.4572e-006, 
    1.822415e-006, 8.121135e-006, 1.280469e-005, -1.00281e-005, 
    -4.81121e-006, -1.078964e-006, 4.506357e-006, -2.220891e-006, 
    -5.093589e-006, -1.554997e-005, -1.101146e-005, -2.184907e-005, 
    -1.126615e-005, -9.353334e-006, 6.934752e-006, 6.343289e-006, 
    6.532544e-006, 1.729988e-005, 2.089652e-005, 1.404186e-005, 9.08822e-006, 
    4.853189e-006, 4.648668e-006,
  3.39908e-006, -1.760818e-006, -1.386921e-006, -6.010883e-006, 
    -8.276103e-006, 2.287074e-006, 4.559879e-006, 1.953256e-005, 
    2.883957e-005, 2.402489e-005, 8.915486e-006, 1.915421e-006, 
    2.829358e-006, 9.899304e-007, 3.447014e-006, 8.134051e-006, 
    1.052171e-005, 1.145403e-005, 1.084246e-005, 5.109974e-006, 
    9.099771e-006, 1.519857e-005, 1.128304e-005, 1.458737e-005, 
    1.300487e-005, 6.610026e-006, 3.353627e-006, 8.53675e-006, 1.383672e-005, 
    1.222963e-005, 8.532661e-006, 1.497393e-005, 1.502671e-005, 
    3.454712e-006, 2.711262e-006, -6.158902e-006, -7.398914e-006, 
    5.61538e-006, -2.75264e-006, 2.469201e-005, 2.158212e-005, 
    -3.329042e-007, -6.055212e-006, -5.469483e-006, -8.877978e-006, 
    -1.81271e-005, -6.538117e-006, -5.429218e-006, -1.265903e-005, 
    -2.381168e-005, -1.792595e-005, 3.50042e-006, 1.185885e-005, 
    1.403267e-005, 5.259732e-006, 9.677562e-006, 1.084307e-005, 
    1.572965e-005, 1.002898e-005, 4.900372e-006, 1.213238e-005, 
    1.273825e-005, 1.402671e-005, 9.585299e-006, 9.518862e-006, 
    7.348131e-006, 7.137034e-006, 9.303418e-006, 4.744781e-006, 
    5.208331e-006, 3.610307e-006, 6.287299e-006, 8.857625e-006, 9.68377e-006, 
    8.652352e-006, 1.76231e-006, -2.431247e-006, 2.484761e-006, 
    -3.346686e-006, 2.729023e-006, 3.634523e-006, 1.794586e-006, 
    -7.614435e-007, -1.573433e-006, -7.011113e-006, -6.014481e-006, 
    -5.74626e-006, 9.820484e-006, 1.449672e-005, 9.151045e-006, 
    1.280767e-005, 1.54201e-005, 1.041405e-005, 1.227731e-005, 1.01873e-005, 
    4.788737e-006,
  4.392488e-006, -2.129564e-007, -1.559281e-006, -5.538514e-006, 
    -8.958079e-006, -9.245552e-006, -2.209955e-005, 5.732218e-006, 
    5.595052e-005, 5.58919e-005, 2.224842e-005, 3.71213e-006, 3.524005e-006, 
    8.334835e-006, 1.220094e-005, 1.059832e-005, 1.202275e-005, 
    8.614235e-006, 7.930645e-006, 6.08054e-006, 1.143503e-005, 9.426225e-006, 
    8.833533e-006, 3.433106e-006, 6.438426e-006, -1.994518e-006, 
    1.012161e-005, 6.684037e-006, 3.868117e-007, 7.966912e-006, 
    5.263828e-006, 1.941733e-005, 1.69019e-006, -2.190587e-006, 
    1.165633e-005, 1.233914e-005, 2.444437e-005, 3.36719e-005, 1.699328e-005, 
    2.334888e-005, 2.939242e-005, 2.028397e-005, -1.208084e-005, 
    -3.394931e-005, -6.183073e-005, -7.244087e-005, -4.771387e-005, 
    -4.549163e-005, -3.3112e-005, -2.687797e-005, -2.808322e-005, 
    -1.65182e-005, -8.715564e-006, -1.761073e-006, 5.825601e-006, 
    1.173119e-005, 1.313301e-005, 1.373093e-005, 1.284368e-005, 
    1.165817e-005, 1.392737e-005, 1.593505e-005, 1.794807e-005, 1.892e-005, 
    1.556053e-005, 1.775337e-005, 1.952461e-005, 1.978811e-005, 
    2.100951e-005, 1.653047e-005, 1.414989e-005, 1.658574e-005, 1.28612e-005, 
    8.868054e-006, -6.68603e-006, 4.272035e-006, 3.560384e-006, 
    -2.99824e-006, -8.305666e-006, -7.07063e-007, -3.823639e-006, 
    -5.137674e-006, 1.131371e-006, 4.846603e-006, 6.325416e-006, 
    7.23017e-006, 9.06003e-006, 1.290601e-005, 1.377835e-005, 9.874137e-006, 
    8.138886e-006, 1.146831e-005, 5.955255e-006, 2.650173e-006, 
    3.302845e-006, 1.780565e-006,
  5.223723e-006, 2.897272e-006, 2.334265e-006, -2.527104e-006, 
    -4.415953e-006, -8.218121e-006, -3.063309e-006, 1.250824e-006, 
    -6.676928e-007, 1.441601e-005, 1.600831e-005, 1.031538e-006, 
    5.960737e-008, 8.33484e-006, 8.254501e-006, 7.912023e-006, 6.023794e-006, 
    1.337382e-006, 2.85655e-006, 1.457454e-006, 9.61245e-007, 3.116944e-006, 
    5.715465e-006, 1.546363e-006, 3.776695e-006, 2.675497e-006, 
    2.810482e-005, 2.590801e-006, -1.104672e-006, 1.723332e-006, 
    1.102139e-005, 1.690985e-005, -2.997491e-006, -4.821399e-006, 
    3.466004e-006, 1.220269e-005, 1.497504e-005, 7.044269e-006, 
    8.053961e-006, 1.425891e-005, 3.575435e-006, 1.234301e-006, 
    -4.311529e-006, -8.490817e-006, -1.568198e-005, -1.204137e-005, 
    -9.031224e-006, -1.030751e-005, -1.071009e-005, -1.096154e-005, 
    -1.095124e-005, -9.936841e-006, -7.266681e-006, -6.153565e-006, 
    -2.518673e-006, 2.796949e-006, 5.981952e-006, 7.704523e-006, 
    7.820008e-006, 7.244203e-006, 6.649397e-006, 5.8764e-006, 6.904829e-006, 
    7.742397e-006, 7.851301e-006, 8.417671e-006, 7.460766e-006, 
    1.279724e-005, 1.479946e-005, 1.515746e-005, 1.778739e-005, 
    1.479735e-005, 1.654352e-005, 5.299982e-006, 4.534792e-006, 
    1.237291e-006, -3.131361e-006, 5.945447e-006, -3.473178e-007, 
    -7.372437e-007, 4.130125e-007, 2.713259e-007, 8.67125e-007, 
    2.428933e-007, -1.193953e-006, -2.022084e-006, -1.979743e-006, 
    -4.3809e-007, 2.929821e-006, 5.491203e-006, 9.345011e-006, 9.455285e-006, 
    1.112918e-005, 7.561721e-006, 9.121992e-006, 6.198141e-006,
  1.773296e-007, 5.081907e-006, 3.417954e-006, -9.35619e-006, -3.502399e-006, 
    -3.634901e-006, 2.785397e-006, 2.482266e-007, -4.443151e-006, 
    1.998978e-005, 2.234193e-005, 6.02255e-006, 6.659458e-006, 5.768363e-006, 
    5.814067e-006, 6.741788e-006, 6.258864e-006, 6.006787e-006, 
    7.375704e-006, 5.461401e-006, 6.343791e-006, 2.984951e-006, 
    1.719218e-006, -2.983463e-006, -3.812962e-006, 7.96864e-006, 
    1.847086e-005, -3.987436e-006, -5.482008e-006, 6.295122e-006, 
    1.263247e-005, -4.116409e-007, 5.595502e-006, 1.534236e-005, 
    1.033136e-005, 9.993208e-006, 8.247298e-006, 1.996222e-005, 
    1.622488e-005, 1.17513e-005, 1.627381e-005, 2.144103e-005, 2.476436e-005, 
    2.660068e-005, 2.393363e-005, 2.352621e-005, 2.030904e-005, 2.13299e-005, 
    2.33675e-005, 2.034095e-005, 1.787581e-005, 1.31689e-005, 1.112099e-005, 
    7.044528e-006, 4.360205e-006, 3.789242e-006, -1.519176e-006, 
    -2.700592e-006, -4.967678e-006, -4.230715e-007, -3.784917e-007, 
    1.4541e-006, 4.942463e-006, 7.830304e-006, 1.126043e-005, 1.324154e-005, 
    1.306024e-005, 1.333418e-005, 1.181997e-005, 1.583931e-005, 
    8.855135e-006, 5.885344e-006, 7.856637e-006, 9.320647e-007, 
    -1.559255e-005, 2.985937e-006, 2.715715e-007, -5.973016e-008, 
    1.322227e-006, -1.90921e-006, -2.513315e-007, 1.285239e-007, 
    1.154876e-007, -1.789503e-006, -2.057103e-006, -1.89853e-006, 
    -1.597775e-006, -1.670045e-006, -1.319248e-006, -6.804858e-007, 
    -5.122265e-007, 6.911687e-007, 2.872195e-006, 1.46106e-006, 
    3.721652e-007, -5.295125e-006,
  -4.462643e-006, -6.635237e-006, -1.309961e-005, -1.397046e-005, 
    -1.63606e-005, -1.19999e-005, -7.007395e-006, -8.100153e-006, 
    -1.042584e-005, -6.676724e-006, -2.052064e-005, -2.597395e-006, 
    -2.367916e-006, -3.700454e-006, 3.636632e-006, 1.083192e-006, 
    -3.551436e-007, 2.991163e-006, 5.796678e-006, 9.572632e-006, 
    1.193061e-005, 4.006797e-006, 1.291686e-006, -5.919501e-007, 
    -5.760048e-006, 3.057095e-006, 1.426152e-005, 1.405549e-006, 
    -4.491583e-006, -8.925039e-006, 1.878798e-007, 8.267154e-006, 
    1.260385e-006, -7.728704e-007, -1.400454e-006, 9.027623e-006, 
    9.617819e-006, 1.788176e-005, 1.094862e-005, 1.573972e-005, 
    2.055081e-005, 1.836592e-005, 1.476382e-005, 1.729031e-005, 
    1.379326e-005, 1.40811e-005, 1.464561e-005, 1.135829e-005, 1.769625e-005, 
    1.472881e-005, 1.215898e-005, 1.250543e-005, 1.363766e-005, 
    1.104027e-005, 7.173661e-006, 5.042673e-006, -7.489107e-007, 
    -7.327772e-006, -1.180619e-005, -1.425234e-005, -1.740356e-005, 
    -1.504458e-005, -1.32593e-005, -9.572754e-006, -5.383543e-006, 
    -1.092629e-006, 7.150815e-006, 9.638563e-006, 9.470183e-006, 
    1.318219e-005, 4.559392e-006, 4.842259e-006, 3.893671e-006, 
    3.156434e-006, -3.251302e-006, 8.727075e-007, 4.799911e-006, 
    -1.369164e-006, -8.052816e-007, -4.64418e-007, 1.659037e-007, 
    -3.738915e-007, -6.921555e-007, -1.798568e-006, -2.178671e-006, 
    -2.593792e-006, -2.174201e-006, -2.42752e-006, -1.167256e-006, 
    -9.648375e-008, -3.861737e-008, 8.939471e-007, -9.136838e-007, 
    -1.270575e-006, 3.818168e-006, 3.065663e-006,
  3.006187e-006, -2.961588e-007, -2.01277e-006, -5.78115e-006, 
    -7.938593e-006, -1.084953e-005, -8.946034e-006, -6.914883e-006, 
    -4.304818e-006, -6.596244e-006, -9.105974e-006, -2.41585e-006, 
    -4.869202e-006, -2.802907e-006, -1.7222e-006, -1.460561e-006, 
    -8.519722e-007, -4.608175e-007, -8.442612e-009, 2.463163e-006, 
    1.338746e-006, 4.669034e-006, 1.472024e-005, 7.732717e-006, 
    5.352245e-006, 3.477311e-006, 6.827588e-006, 1.680019e-005, 
    2.499797e-006, -1.092963e-005, -3.603476e-006, -1.170491e-006, 
    -1.705066e-006, -1.31217e-006, 3.388148e-006, 6.199629e-006, 
    1.101742e-005, 1.442159e-005, 7.223956e-006, 7.186823e-006, 
    2.949186e-006, 4.121415e-006, 2.264733e-006, 5.57018e-006, 6.94295e-006, 
    4.164755e-006, 1.79013e-006, 2.822658e-006, 2.997621e-006, 1.873204e-006, 
    4.111516e-007, 1.776967e-006, 3.356244e-006, 6.000701e-006, 
    3.881135e-006, 2.17607e-006, -5.964175e-007, -6.805607e-006, 
    -1.014297e-005, -7.124242e-006, -6.486101e-006, -5.368638e-006, 
    -6.795673e-006, -4.198152e-006, -2.944219e-006, -3.331774e-006, 
    -4.818412e-006, -4.631165e-006, 5.274145e-006, 1.193583e-005, 
    7.862604e-006, 3.177924e-006, -1.266843e-006, -7.140106e-007, 
    -4.439262e-007, 3.056355e-006, 5.478289e-006, 4.657484e-006, 
    2.79223e-006, 1.38072e-006, 1.100234e-007, -6.674445e-007, 
    -1.437711e-006, -1.93392e-006, -1.732629e-006, -2.112486e-006, 
    -1.668928e-006, -1.586599e-006, -9.665873e-007, -5.24147e-007, 
    -4.234255e-008, -8.692211e-008, -7.351105e-008, -3.597374e-007, 
    3.390028e-007, 7.941098e-007,
  -3.432977e-006, -4.265579e-006, -2.534314e-006, -2.381949e-006, 
    -1.903995e-006, -1.002971e-006, -1.705437e-006, -1.290812e-006, 
    -1.457829e-006, -1.495455e-006, -1.496324e-006, -1.722821e-006, 
    -4.423905e-006, -2.318247e-006, -1.2774e-006, -1.56164e-006, 
    -3.933894e-007, -3.725143e-008, -6.618484e-008, 4.448007e-007, 
    9.370359e-007, 1.016012e-006, 1.113414e-005, 8.611372e-006, 
    3.972773e-006, 4.56808e-006, 6.57427e-006, 8.574753e-006, 6.605434e-006, 
    -1.107889e-005, -8.185336e-006, -8.046009e-006, -7.375209e-006, 
    -5.062175e-006, 5.435195e-007, 2.728524e-006, 4.178033e-006, 
    6.42823e-006, 5.698475e-007, 1.780196e-006, -2.188355e-006, 
    -2.315015e-006, 1.413173e-007, 4.295298e-007, 3.241378e-006, 
    2.575918e-006, 1.630314e-006, 1.353525e-006, 1.225653e-007, 
    -1.706924e-006, -3.448125e-006, -1.248714e-006, 3.572586e-007, 
    3.184382e-006, 4.275272e-006, 2.710151e-006, 1.277653e-006, 
    -3.647305e-006, -8.605419e-006, -8.379789e-006, -5.182e-006, 
    -5.934013e-006, -5.959593e-006, -3.936014e-006, -2.347304e-006, 
    -1.878911e-006, -2.788999e-006, -5.134939e-006, -7.892277e-006, 
    -3.723182e-006, 1.535063e-006, -3.326686e-006, -3.232678e-006, 
    -2.899487e-007, -7.054423e-007, 1.217055e-006, 2.052886e-006, 
    3.061695e-006, 1.508373e-006, 5.84625e-007, -1.09645e-007, 
    -7.316439e-007, -8.651341e-007, -1.17036e-006, -1.264732e-006, 
    -1.702207e-006, -2.170725e-006, -1.606219e-006, -1.201405e-006, 
    -5.7419e-007, -9.08957e-008, -1.626569e-008, -4.730981e-008, 
    8.891163e-008, 3.793599e-007, -1.216058e-006,
  -1.477324e-006, -2.394864e-006, -2.540894e-006, -2.16911e-006, 
    -1.158689e-006, -1.510232e-006, -1.350044e-006, -9.444836e-007, 
    -7.849171e-007, -1.447895e-006, -2.585226e-006, -1.649681e-006, 
    -2.842892e-006, -1.624225e-006, -1.990421e-006, -2.036367e-006, 
    -1.717109e-006, -1.842759e-007, 6.680813e-008, 5.092488e-007, 
    5.407894e-007, 3.454599e-007, 2.188981e-006, 6.92507e-006, 1.038251e-005, 
    6.903834e-006, 6.281339e-006, 1.155511e-005, 8.091823e-006, 
    -2.709405e-006, -5.122643e-006, -7.029594e-007, -1.872084e-006, 
    -8.349245e-006, -5.775941e-006, -2.619501e-006, -1.564622e-006, 
    -3.141289e-006, -2.643092e-006, -9.431133e-007, -1.574553e-006, 
    -2.757581e-006, -2.225857e-006, 3.486921e-007, 1.062456e-006, 
    2.336383e-006, 1.561025e-006, 7.763547e-007, -5.613965e-007, 
    -5.334578e-007, -3.576242e-007, 9.84599e-007, 3.861518e-006, 
    5.913776e-006, 3.796324e-006, 2.163404e-006, -9.015148e-007, 
    -1.509943e-007, -2.028168e-006, -5.279848e-006, -8.120756e-006, 
    -3.968425e-006, -3.419441e-006, -3.026797e-006, -2.296019e-006, 
    -2.950056e-006, -1.966455e-006, -1.123785e-007, -1.728036e-006, 
    -8.389728e-006, -1.110559e-005, -8.594619e-006, -4.238633e-006, 
    -5.779129e-007, -1.824768e-006, -1.948199e-006, -1.453232e-006, 
    -1.981807e-007, -5.383026e-007, -9.556597e-007, -1.022342e-006, 
    -2.318743e-006, -1.644466e-006, -1.014022e-006, -1.298758e-006, 
    -1.431502e-006, -1.742067e-006, -1.824148e-006, -1.404433e-006, 
    -8.627762e-007, -4.974492e-007, -2.498414e-007, 9.33311e-007, 
    1.8639e-007, 2.807641e-007, 1.091523e-007,
  -7.352469e-007, -2.192456e-006, -3.433101e-006, -3.125641e-006, 
    -2.266838e-006, -2.357362e-006, -2.692762e-006, -2.659483e-006, 
    -1.628819e-006, -1.470371e-006, -2.579514e-006, -3.41994e-006, 
    -4.005803e-006, -3.986556e-006, -3.091244e-006, -2.380335e-006, 
    -3.510092e-006, -2.283974e-006, -9.592609e-007, -9.375179e-008, 
    3.457083e-007, 1.341603e-006, 2.005822e-006, 2.547355e-006, 
    4.246461e-006, 7.244947e-006, 2.871952e-006, 5.718945e-006, 
    1.170113e-005, 4.261608e-006, -9.3977e-007, -2.610561e-006, 
    -1.902754e-006, -4.314392e-006, -6.481261e-006, -4.068888e-006, 
    7.696144e-009, -8.770585e-007, -2.841898e-006, -4.690137e-006, 
    -1.898155e-006, 8.456846e-008, -2.383063e-006, -2.405043e-006, 
    -7.946983e-008, -4.944668e-007, -2.397801e-007, -8.527159e-007, 
    -8.049083e-007, -3.113064e-007, 5.203019e-007, 1.015642e-006, 
    4.47507e-006, 6.639464e-006, 4.466254e-006, 1.303109e-006, 
    -7.747331e-007, -2.433978e-006, -8.648849e-007, -2.25501e-007, 
    -2.849721e-006, -4.911295e-006, -5.372736e-006, -3.522136e-006, 
    -1.73052e-006, -1.584613e-006, -1.200411e-006, -1.939508e-006, 
    -3.401437e-006, -7.962935e-006, -5.553913e-006, -4.593036e-006, 
    -5.294261e-006, -5.235152e-006, -3.933286e-006, -2.515562e-006, 
    -1.154214e-006, 7.572307e-007, -5.735656e-007, -2.955145e-006, 
    -2.455583e-006, -1.659242e-006, -1.780809e-006, -4.503854e-007, 
    -6.796154e-007, -1.004461e-006, -1.149499e-006, -1.531464e-006, 
    -1.088155e-006, -1.20364e-006, -1.113736e-006, -5.523351e-007, 
    5.230322e-007, 1.462427e-006, 1.170984e-006, 6.124391e-007,
  1.273306e-006, 2.266235e-007, -1.526995e-006, -2.637256e-006, 
    -1.860781e-006, -1.872081e-006, -1.826757e-006, -3.244478e-006, 
    -3.174815e-006, -1.961613e-006, -2.030531e-006, -2.369159e-006, 
    -3.967929e-006, -6.15815e-006, -4.379326e-006, -4.28222e-006, 
    -6.311262e-006, -6.606678e-006, -3.346179e-006, -1.564744e-006, 
    -1.527244e-006, -1.399453e-007, 1.942492e-006, 2.200406e-006, 
    2.502405e-006, 1.704246e-005, 1.683992e-005, 1.036823e-005, 
    8.665649e-006, 1.257051e-005, 1.113935e-005, 2.233683e-006, 
    3.770743e-006, 1.343215e-006, -6.348881e-006, -6.495044e-006, 
    -3.71995e-006, -2.085297e-006, -1.634908e-006, -1.124296e-006, 
    -3.561254e-006, -1.980985e-006, -1.616736e-007, -3.048526e-006, 
    -1.744798e-006, -5.987731e-007, -9.115738e-007, -5.397915e-007, 
    -1.498681e-006, 2.050183e-007, -3.676823e-007, 1.840669e-006, 
    3.575786e-006, 3.964955e-006, 2.656758e-006, 6.013897e-007, 
    -1.980983e-006, -3.304703e-006, -1.887603e-006, -2.030031e-006, 
    -6.894234e-007, -1.223383e-006, -2.699096e-006, -2.688168e-006, 
    -3.005438e-006, -9.102114e-007, -3.320463e-007, -1.092005e-006, 
    -2.919012e-006, -4.970158e-006, 4.970771e-007, -2.410512e-006, 
    -2.636889e-006, -3.861887e-006, -3.357854e-006, -7.511675e-006, 
    -7.136421e-006, -3.76838e-006, -3.955889e-006, -5.239499e-006, 
    -4.606942e-006, -2.687302e-006, -2.416096e-006, -8.533361e-007, 
    -8.139705e-007, -1.584736e-006, -6.680666e-007, -1.915417e-006, 
    -5.700922e-007, -9.365372e-007, -2.056234e-006, -7.168692e-007, 
    -4.213289e-007, 4.341219e-007, 7.1712e-007, 1.424552e-006,
  -1.241751e-007, -2.780296e-007, 3.975174e-009, -1.160551e-006, 
    -9.108321e-007, -5.044026e-007, -1.064563e-006, -2.798809e-006, 
    -3.056475e-006, -2.848231e-006, -2.919136e-006, -2.411627e-006, 
    -1.730396e-006, -3.286201e-006, -5.895393e-006, -4.947928e-006, 
    -6.249667e-006, -9.895114e-006, -1.09336e-005, -4.467118e-006, 
    -1.925974e-006, -5.254273e-006, 7.189847e-007, 4.127633e-007, 
    -7.332592e-007, 1.640373e-006, 9.99359e-006, 2.056956e-005, 
    1.773958e-005, 1.288118e-005, 1.264314e-005, 6.469585e-006, 
    4.183457e-007, 2.131863e-006, -2.420202e-007, -4.553549e-006, 
    -6.434952e-006, -7.813142e-007, -2.025565e-006, -1.442186e-006, 
    -3.673158e-007, -3.201887e-006, -3.788995e-006, -2.495206e-006, 
    -5.200633e-006, -5.002694e-006, -4.06541e-006, -1.223008e-006, 
    -3.555124e-007, -1.091383e-006, -2.172692e-008, 2.15707e-006, 
    3.904108e-006, 3.907337e-006, 3.484393e-006, 1.936907e-006, 
    -2.295272e-006, -3.076713e-006, -3.833073e-006, -3.900499e-006, 
    -2.901501e-006, -1.831599e-006, -1.872576e-006, -1.530348e-006, 
    -1.791366e-006, -1.559654e-006, -1.059968e-006, -9.347982e-007, 
    -2.019974e-006, -3.066035e-006, -2.04891e-006, -4.961592e-006, 
    -5.002075e-006, -5.731483e-006, -8.375198e-006, -7.237992e-006, 
    -1.013167e-005, -1.126913e-005, -8.843846e-006, -4.722431e-006, 
    -7.752205e-006, -7.23936e-006, -5.559377e-006, -3.957748e-006, 
    -2.438079e-006, -7.996914e-007, -4.965787e-007, -2.25181e-006, 
    -6.547798e-007, -1.12019e-006, -9.18159e-007, -9.136884e-007, 
    -1.384193e-006, -1.360351e-006, -2.1105e-006, -2.067411e-006,
  -4.028898e-006, -2.410757e-006, -2.880515e-006, -3.055978e-006, 
    -1.043326e-006, 1.610588e-007, -1.240518e-006, -1.018989e-006, 
    -2.535553e-006, -3.271049e-006, -3.506118e-006, -3.897273e-006, 
    -5.801765e-006, -1.185089e-005, -1.078099e-005, -6.140393e-006, 
    -8.788453e-006, -1.428475e-005, -1.519335e-005, -1.038773e-005, 
    -5.939844e-006, -2.950928e-006, 3.710642e-006, 1.853214e-006, 
    9.649757e-007, 1.13274e-006, -1.152352e-006, 2.086286e-006, 
    1.602061e-005, 1.881445e-005, 1.564287e-005, 1.285101e-005, 
    6.370246e-006, 5.645434e-006, 8.042407e-006, 6.953756e-006, 
    6.856033e-006, 6.698698e-006, 5.82535e-006, 2.228095e-006, 
    -4.245594e-007, -4.124646e-006, -4.654747e-006, -5.635371e-006, 
    -5.802995e-006, -8.269519e-006, -8.916108e-006, -6.417813e-006, 
    -7.737432e-006, -4.543615e-006, 3.36513e-008, 4.209323e-008, 
    -2.373385e-006, 8.707211e-007, 6.920327e-007, -4.598242e-007, 
    -3.097079e-006, -5.663431e-006, -4.651145e-006, -4.41372e-006, 
    -4.07025e-006, -2.298005e-006, -5.184329e-007, -2.868437e-007, 
    -1.634159e-006, -3.621228e-006, -2.9431e-006, -3.194062e-006, 
    -4.266944e-006, -3.789615e-006, -2.345072e-006, -4.586709e-006, 
    -1.279041e-007, 2.049655e-006, -7.025883e-007, -9.518117e-007, 
    -2.058718e-006, -8.782623e-006, -1.259285e-005, -8.016326e-006, 
    -4.477679e-006, -6.190938e-006, -8.716557e-006, -6.228565e-006, 
    -6.404145e-006, -6.771465e-006, -2.707047e-006, -1.972659e-006, 
    -3.458928e-006, -1.741443e-006, -4.27659e-007, -1.922868e-006, 
    -2.285338e-006, -3.018353e-006, -5.810208e-006, -5.148967e-006,
  -4.663318e-006, -4.462521e-006, -4.661575e-006, -6.217382e-006, 
    -2.852326e-006, -1.882387e-006, -1.483533e-006, -5.956717e-007, 
    -6.403807e-007, -9.172945e-007, -5.084985e-007, -3.922851e-006, 
    -3.89802e-006, -2.771365e-006, -3.792838e-006, -5.55403e-006, 
    -6.502863e-006, -5.882851e-006, -6.637227e-006, -6.715705e-006, 
    2.371744e-007, 4.525859e-006, 3.305948e-006, 2.449008e-006, 
    1.657634e-006, 4.26012e-006, 3.372634e-006, 1.642979e-006, 8.227549e-006, 
    1.212123e-005, 1.211724e-005, 1.364859e-005, 1.437552e-005, 
    1.143602e-005, 1.072958e-005, 9.169798e-006, 6.272272e-006, 
    4.675985e-006, 6.136546e-006, 6.629154e-006, 3.322464e-006, 
    1.695131e-006, 6.601185e-007, -9.650976e-007, -2.12602e-006, 
    -1.10182e-006, -9.597497e-007, -5.566326e-006, -7.276853e-006, 
    -8.123989e-006, -4.994872e-006, -1.151988e-006, -1.109394e-006, 
    -8.158531e-008, 2.822151e-006, -5.920738e-007, -2.20997e-006, 
    -3.906342e-006, -5.292273e-006, -4.668411e-006, -3.122166e-006, 
    -3.721561e-007, 3.777448e-006, 3.816192e-006, 8.615389e-007, 
    -2.636754e-006, 3.193854e-007, 2.274946e-007, -6.487719e-006, 
    -9.435915e-006, -3.489606e-006, -9.45729e-007, 1.162414e-006, 
    7.755676e-006, 1.023971e-005, 6.225953e-006, 4.207461e-006, 
    -3.026253e-007, -2.478311e-006, -4.485366e-006, -2.514073e-006, 
    1.927841e-006, 1.420449e-006, -4.360951e-006, -1.025969e-005, 
    -8.905427e-006, -8.676827e-006, -6.166851e-006, -3.58845e-006, 
    -5.749986e-006, -4.592415e-006, -3.283596e-006, -3.697223e-006, 
    -4.158909e-006, -2.532821e-006, -3.334007e-006,
  3.588648e-007, -8.015559e-007, -2.864497e-006, -4.616131e-006, 
    -1.12851e-006, 2.150236e-006, 1.304965e-006, 3.952555e-007, 
    9.628657e-007, 2.28124e-006, 4.331514e-006, 4.739559e-006, 2.342953e-006, 
    -1.411882e-006, -2.873809e-006, -1.51768e-006, -1.814709e-006, 
    -2.084793e-006, -1.204756e-006, -8.430325e-007, 7.799499e-007, 
    3.340472e-006, 2.358361e-006, 1.252693e-006, 6.010146e-007, 
    7.318968e-007, 1.962607e-006, 2.788133e-006, 3.316378e-006, 
    5.195044e-006, 5.402547e-006, 3.225732e-006, 1.859174e-006, 2.2733e-006, 
    2.121804e-006, 4.071493e-006, 3.847847e-006, 2.731256e-006, 3.92372e-006, 
    7.107472e-006, 5.978469e-006, 7.550414e-006, 7.498384e-006, 
    3.800298e-006, 4.988284e-006, 4.339461e-006, 4.433223e-006, 
    5.011389e-006, 3.616515e-006, -2.860979e-007, 1.522421e-007, 
    -3.439683e-006, -3.780671e-006, 6.489463e-007, 3.982204e-006, 
    3.400815e-006, 2.159046e-006, -1.065309e-006, -1.18055e-006, 
    -4.753492e-007, 4.873909e-007, 3.445519e-006, 7.35968e-006, 
    8.517376e-006, 9.34464e-006, 7.072838e-006, 3.15669e-006, 1.616656e-006, 
    -1.543522e-007, -4.023565e-006, -2.214687e-006, 2.084045e-006, 
    4.762533e-006, 5.075581e-006, 5.304062e-006, 3.070007e-006, 
    4.832567e-006, 5.398815e-006, 1.911685e-006, 2.739082e-006, 
    4.901984e-006, 3.59739e-006, 6.092589e-006, 9.681036e-006, 
    -6.576374e-007, -7.275248e-006, -5.904712e-006, -8.022784e-006, 
    -7.989383e-006, -6.781147e-006, -5.627549e-006, -3.752486e-006, 
    -2.139685e-006, -2.004952e-006, -2.510606e-006, -3.950303e-006,
  5.035474e-006, 2.686807e-006, -5.35827e-007, 1.152228e-006, 6.204971e-006, 
    8.553268e-006, 1.046483e-005, 5.065032e-006, 3.559147e-006, 
    1.955408e-006, 4.862625e-006, 1.012261e-005, 8.43853e-006, 2.133104e-006, 
    1.358245e-006, 2.690656e-006, 1.007195e-006, 7.8219e-007, -4.906169e-007, 
    1.423187e-006, 2.953661e-006, 3.518664e-006, 1.396366e-006, 
    1.543888e-006, 2.387292e-006, 2.235674e-006, 1.448025e-006, 
    1.400836e-006, 1.32012e-006, 7.479175e-007, 1.742569e-006, 1.181541e-006, 
    2.288325e-006, 3.046174e-006, 2.833831e-006, 8.499901e-007, 
    9.387768e-007, 3.949055e-006, 3.504381e-006, 9.29447e-006, 7.556122e-006, 
    5.248807e-006, 4.961956e-006, 8.907904e-006, 8.193525e-006, 
    9.767828e-006, 8.108713e-006, 6.581467e-006, 5.587684e-006, 
    6.056445e-006, 3.696347e-006, 3.548583e-006, 4.617617e-006, 
    3.755707e-006, 4.308542e-006, 4.832444e-006, 3.070003e-006, 
    3.425645e-006, 2.802899e-006, 3.651645e-006, 2.999106e-006, 
    4.648413e-006, 8.853771e-006, 1.256329e-005, 1.140609e-005, 
    7.501743e-006, 4.310287e-006, 5.02219e-006, 6.154802e-006, 4.132467e-006, 
    6.606304e-006, 1.11072e-005, 9.388346e-006, 4.408381e-006, 5.48859e-006, 
    5.749982e-006, 1.128278e-005, 9.051335e-006, 6.565326e-006, 
    4.919486e-006, 2.992649e-006, 4.040696e-006, 7.623308e-006, 
    7.302682e-006, 3.312522e-006, 2.659977e-006, 6.657028e-007, 2.42814e-006, 
    -1.64584e-006, -6.162256e-006, -5.17282e-006, -5.356478e-006, 
    -1.931072e-006, -9.612559e-007, 1.137414e-007, 2.848354e-006,
  2.960491e-006, 7.609147e-006, 8.4903e-006, 6.861983e-006, 3.496933e-006, 
    4.980468e-006, 5.95786e-006, 6.321326e-006, 4.801657e-006, 3.331159e-006, 
    3.486254e-006, 3.310049e-006, 2.317134e-006, 9.586438e-007, 
    9.128235e-007, 2.322349e-006, 2.304716e-006, 1.688055e-006, 
    1.495831e-006, 9.87081e-007, 1.187997e-006, 1.628946e-006, 3.908703e-006, 
    4.336491e-006, 3.502647e-006, 2.729771e-006, 2.618013e-006, 
    1.577043e-006, 4.592066e-007, 5.49483e-007, 1.954909e-006, 1.509989e-006, 
    8.119914e-007, 1.60821e-006, 2.223628e-006, 2.344453e-006, 2.930442e-006, 
    5.573535e-006, 2.498929e-006, 4.694737e-006, 6.370374e-006, 
    5.128604e-006, 7.166836e-006, 8.393945e-006, 1.024231e-005, 
    6.234886e-006, 5.833672e-006, 6.141505e-006, 2.645324e-006, 
    2.785395e-006, 3.022076e-006, 3.908319e-006, 4.401054e-006, 
    5.237755e-006, 4.454201e-006, 3.653764e-006, 2.587331e-006, 
    4.683056e-006, 7.530669e-006, 4.9591e-006, 5.058939e-006, 5.075206e-006, 
    6.034476e-006, 9.884807e-006, 1.002463e-005, 4.682819e-006, 
    3.853444e-006, 4.73609e-006, 5.893909e-006, 6.331634e-006, 4.583103e-006, 
    6.311515e-006, 9.592748e-006, 1.001234e-005, 7.811686e-006, 
    8.723888e-006, 9.360663e-006, 9.309006e-006, 8.101139e-006, 
    7.538116e-006, 5.255011e-006, 4.22162e-006, 3.49022e-006, 3.456818e-006, 
    4.301215e-006, 6.627779e-006, 7.572147e-006, 5.803377e-006, 1.87655e-006, 
    5.03278e-007, -8.096358e-007, -2.974648e-006, -5.891015e-007, 
    2.738831e-006, 5.380498e-007, 1.797209e-006,
  4.530453e-006, 4.238641e-006, 3.932544e-006, 5.186973e-006, 5.854921e-006, 
    3.63055e-006, 3.210831e-006, 2.983837e-006, 2.096227e-006, 1.82254e-006, 
    8.160896e-007, 2.803656e-006, 4.625696e-006, 2.811107e-006, 
    8.930792e-007, 4.799449e-007, 2.791521e-007, -1.737212e-007, 
    5.64879e-007, 9.314508e-007, 5.589191e-007, 6.318105e-007, 9.781406e-007, 
    2.546115e-006, 3.505749e-006, 3.441674e-006, 3.123286e-006, 
    3.846987e-006, 2.865745e-006, 1.71314e-006, 2.131738e-006, 3.461297e-006, 
    3.362699e-006, 1.540907e-006, 1.541777e-006, 2.005328e-006, 2.31825e-006, 
    3.339975e-006, 2.114353e-006, 2.645457e-006, 3.60683e-006, 4.714109e-006, 
    6.920103e-006, 5.937247e-006, 5.687272e-006, 6.040435e-006, 
    5.334738e-006, 4.211068e-006, 4.006051e-006, 3.492954e-006, 
    4.946191e-006, 3.816185e-006, 4.634883e-006, 3.543868e-006, 
    3.995499e-006, 4.066773e-006, 2.975135e-006, 2.855057e-006, 
    7.948527e-006, 6.746746e-006, 6.197512e-006, 5.016595e-006, 
    5.299346e-006, 6.493919e-006, 3.741188e-006, 3.178546e-006, 
    4.063922e-006, 6.894397e-006, 7.008392e-006, 3.282107e-006, 
    2.314649e-006, 2.771372e-006, 4.275643e-006, 4.292905e-006, 
    5.106382e-006, 5.27489e-006, 6.788721e-006, 7.004788e-006, 4.725161e-006, 
    2.29366e-006, -7.969666e-007, -1.341105e-006, -1.176821e-006, 
    -8.730858e-007, 1.239154e-006, 2.338238e-006, 4.056716e-006, 
    2.416966e-006, -1.395869e-006, -1.225002e-006, 7.970812e-007, 
    1.757466e-006, 1.518178e-006, 2.464774e-006, 3.722183e-006, 4.02269e-006,
  5.354485e-006, 6.47468e-006, 7.281205e-006, 8.114429e-006, 5.025917e-006, 
    1.966832e-006, 2.393998e-006, 4.300728e-006, 5.296619e-006, 
    1.396369e-006, 1.028183e-006, 1.820304e-006, 1.944357e-006, 
    2.175324e-006, 2.162907e-006, 2.824643e-006, 2.356747e-006, 
    1.580644e-006, 1.653534e-006, 1.663592e-006, 1.766039e-006, 2.18352e-006, 
    2.551827e-006, 2.670788e-006, 2.914794e-006, 2.793598e-006, 
    2.648063e-006, 2.574798e-006, 2.316014e-006, 2.275161e-006, 
    1.076861e-006, -1.344815e-007, 1.728536e-006, 2.917649e-006, 
    3.26075e-006, 2.96757e-006, 2.991535e-006, 3.294525e-006, 1.93318e-006, 
    2.067166e-006, 2.924729e-006, 3.058715e-006, 3.332648e-006, 4.15482e-006, 
    2.588458e-006, 2.910572e-006, 4.960351e-006, 5.798791e-006, 
    6.205839e-006, 6.779039e-006, 5.468853e-006, 3.045305e-006, 2.94944e-006, 
    2.85494e-006, 2.769757e-006, 2.777826e-006, 4.117188e-006, 6.768354e-006, 
    7.087609e-006, 6.078177e-006, 4.182381e-006, 4.679583e-006, 
    1.749891e-006, 2.546863e-006, 2.602987e-006, 2.485515e-006, 
    1.909212e-006, 3.409015e-006, 4.403421e-006, 2.400952e-006, 
    7.448116e-007, 1.591198e-006, 4.128495e-006, 5.927684e-006, 
    5.522374e-006, 5.25378e-006, 5.184739e-006, 4.124894e-006, 1.900521e-006, 
    2.071636e-006, -4.985632e-007, -5.879738e-007, 1.265609e-006, 
    -1.947064e-007, -1.674143e-006, -8.48624e-007, -8.790466e-007, 
    5.66366e-007, -7.445615e-007, -1.123923e-006, 1.953913e-006, 
    8.292482e-007, 2.518915e-006, 3.819661e-006, 1.791988e-006, 3.161904e-006,
  2.199789e-006, 4.03797e-006, 5.561987e-006, 6.2606e-006, 8.531286e-006, 
    7.930403e-006, 5.102287e-006, 5.059817e-006, 5.700321e-006, 
    4.123774e-006, 2.509607e-006, 2.891325e-006, 3.945211e-006, 
    4.304577e-006, 2.162534e-006, 1.430019e-006, 3.028167e-006, 
    2.762059e-006, 1.467767e-006, 2.096131e-007, 6.407527e-007, 
    2.371399e-006, 3.388155e-006, 3.817308e-006, 4.032382e-006, 
    2.969556e-006, 2.794715e-006, 2.348053e-006, 2.235921e-006, 
    2.055369e-006, 1.885744e-006, 1.212707e-006, 1.292925e-006, 
    1.179925e-006, 1.446159e-006, 2.39052e-006, 2.162656e-006, 2.964464e-006, 
    2.197427e-006, 1.79671e-006, 2.290933e-006, 2.02656e-006, 1.604983e-006, 
    2.816695e-006, 2.552323e-006, 3.055362e-006, 3.377848e-006, 
    4.377467e-006, 6.443142e-006, 4.75186e-006, 3.797069e-006, 2.869222e-006, 
    3.54052e-006, 4.011769e-006, 3.767762e-006, 4.070502e-006, 2.839162e-006, 
    1.178181e-006, 3.591122e-007, 2.625331e-006, 2.803285e-006, 
    2.558906e-006, 1.462553e-006, -1.860135e-007, 1.219428e-007, 
    3.109385e-007, 7.280469e-007, 1.675761e-006, 3.451857e-006, 
    4.506238e-006, 3.784027e-006, 3.449247e-006, 3.609062e-006, 
    3.696855e-006, 3.876662e-006, 2.910322e-006, 2.586969e-006, 
    3.386664e-006, 2.08567e-006, 2.540899e-006, 1.667071e-006, 1.160432e-006, 
    5.168258e-007, 6.49572e-007, 1.783668e-006, 4.826707e-007, 
    -1.820179e-006, -3.283276e-007, 5.575494e-007, 1.172471e-006, 
    8.435309e-007, 1.148508e-006, 1.958388e-006, 9.926644e-007, 
    1.453232e-006, 1.816703e-006,
  -1.412003e-006, 3.931455e-007, 9.813702e-007, 1.743936e-006, 2.046926e-006, 
    3.648305e-006, 4.560256e-006, 5.375598e-006, 7.030746e-006, 
    5.750736e-006, 3.209589e-006, 3.705052e-006, 3.937013e-006, 
    3.526487e-006, 2.248464e-006, 1.531842e-006, 1.566362e-006, 
    1.579526e-006, 1.958139e-006, 2.12615e-006, 1.989803e-006, 2.409022e-006, 
    2.470119e-006, 1.810494e-006, 1.9718e-006, 2.532332e-006, 2.346439e-006, 
    1.897293e-006, 1.358615e-006, 1.442061e-006, 1.425794e-006, 
    1.574185e-006, 1.728411e-006, 1.61777e-006, 1.266103e-006, 1.105419e-006, 
    1.257783e-006, 1.389906e-006, 1.661605e-006, 2.021467e-006, 
    1.798323e-006, 1.568473e-006, 1.267469e-006, 1.582877e-006, 
    1.925977e-006, 3.505997e-006, 4.844868e-006, 5.271289e-006, 
    4.494691e-006, 3.145764e-006, 2.829112e-006, 3.254665e-006, 
    3.535303e-006, 3.394613e-006, 2.374876e-006, 2.201154e-006, 
    2.518798e-006, 1.975649e-006, 6.48577e-007, 1.308845e-007, 8.3546e-007, 
    7.717572e-007, 7.296612e-007, 1.279141e-006, 1.432623e-006, 
    1.467641e-006, 1.415984e-006, 1.617026e-006, 2.130743e-006, 
    1.921878e-006, 1.59368e-006, 2.323713e-006, 2.318746e-006, 2.532951e-006, 
    2.890826e-006, 1.747163e-006, 1.053264e-006, 1.367928e-006, 1.25468e-006, 
    7.95103e-007, 1.239305e-007, 7.883982e-007, 1.176325e-006, 1.30638e-007, 
    -1.207118e-006, -2.805145e-006, -2.788382e-006, -3.437084e-006, 
    1.206743e-006, 2.657373e-006, 9.1332e-007, 1.06671e-007, -1.054213e-007, 
    4.991925e-007, 4.325102e-007, -9.256073e-007,
  -1.223257e-006, -2.923603e-006, -3.029152e-006, -3.343941e-006, 
    -2.48998e-006, 5.011789e-007, 1.631682e-006, 2.209969e-006, 
    2.382326e-006, 2.85134e-006, 3.588078e-006, 3.421185e-006, 2.436714e-006, 
    2.199786e-006, 2.347308e-006, 2.032148e-006, 1.60287e-006, 1.18663e-006, 
    9.883206e-007, 8.294992e-007, 9.597602e-007, 1.793729e-006, 
    2.069897e-006, 1.766784e-006, 2.126274e-006, 1.965838e-006, 
    2.080949e-006, 1.956399e-006, 1.415611e-006, 3.365185e-007, 
    -1.944595e-007, 1.558424e-007, 2.412762e-007, 5.631405e-007, 
    9.89065e-007, 9.249916e-007, 9.343039e-007, 1.377613e-006, 1.705687e-006, 
    2.121553e-006, 2.051145e-006, 1.374136e-006, 1.18663e-006, 1.550715e-006, 
    1.850974e-006, 2.089019e-006, 3.126761e-006, 3.308807e-006, 
    2.521528e-006, 2.703693e-006, 2.315393e-006, 1.991541e-006, 2.15595e-006, 
    2.568712e-006, 2.293911e-006, 1.349053e-006, 1.185895e-007, 
    -2.266211e-007, 2.772872e-007, 2.074989e-007, 1.528624e-007, 
    2.607749e-008, 5.175684e-007, 6.673254e-007, 6.232417e-007, 
    5.484881e-007, 1.221027e-006, 1.486764e-006, 1.129137e-006, 
    8.281331e-007, 1.484404e-006, 1.947583e-006, 1.891207e-006, 
    1.712145e-006, 1.037371e-006, 8.739548e-007, 8.398056e-007, 
    7.237009e-007, 2.923125e-007, 1.772005e-007, 3.530345e-007, 
    6.825976e-007, 6.577629e-007, 1.511253e-007, -9.742835e-007, 
    -1.941867e-006, -2.148e-006, -1.05301e-006, 1.328817e-006, 2.292672e-006, 
    2.961235e-006, 3.187484e-006, 1.777587e-006, 7.720073e-007, 
    5.684833e-007, -5.364018e-008,
  -9.680762e-007, -1.407411e-006, -2.25355e-006, -2.169605e-006, 
    -1.253307e-006, -9.970972e-008, 1.02272e-006, 2.310552e-006, 
    3.288316e-006, 3.526734e-006, 3.298125e-006, 3.294399e-006, 
    3.046419e-006, 2.264977e-006, 1.795093e-006, 1.236425e-006, 
    8.831435e-007, 1.323969e-006, 2.189478e-006, 2.425165e-006, 
    2.406662e-006, 2.153095e-006, 2.202268e-006, 2.121802e-006, 
    2.193701e-006, 2.634403e-006, 2.511095e-006, 2.111496e-006, 
    1.879534e-006, 1.210597e-006, 5.940608e-007, 2.118461e-007, 
    1.902397e-007, 2.928091e-007, 3.226116e-007, 6.566456e-007, 
    8.943198e-007, 1.002974e-006, 1.424552e-006, 1.385437e-006, 
    1.469504e-006, 1.670173e-006, 2.044814e-006, 1.954786e-006, 
    1.797951e-006, 1.750888e-006, 1.207492e-006, 1.06084e-006, 7.017213e-007, 
    6.924085e-007, 8.014354e-007, 8.724646e-007, 8.227939e-007, 
    9.809946e-007, 1.154841e-006, 9.88694e-007, 1.029424e-006, 1.149378e-006, 
    1.082944e-006, 8.590539e-007, 7.186102e-007, 8.066511e-007, 
    1.114111e-006, 1.13398e-006, 1.309069e-006, 1.142052e-006, 1.227733e-006, 
    1.62547e-006, 1.348433e-006, 8.578113e-007, 9.894379e-007, 1.487137e-006, 
    1.882514e-006, 1.609078e-006, 8.585562e-007, 2.900761e-007, 
    2.945476e-007, 8.832671e-007, 1.185389e-006, 8.126108e-007, 
    5.642585e-007, 6.519267e-007, 3.81719e-007, -7.822973e-008, 
    1.110147e-007, 4.49023e-007, 6.737821e-007, 1.363334e-006, 2.081693e-006, 
    2.263365e-006, 2.784906e-006, 2.842151e-006, 2.225616e-006, 
    9.996229e-007, -2.818524e-008, -5.602824e-007,
  9.768983e-007, 1.051901e-006, 1.111754e-006, 9.869564e-007, 1.001237e-006, 
    9.19279e-007, 1.010673e-006, 1.472857e-006, 1.66384e-006, 1.532958e-006, 
    1.754986e-006, 2.287702e-006, 2.403558e-006, 2.208974e-006, 1.8131e-006, 
    1.443799e-006, 1.270201e-006, 1.35017e-006, 1.843523e-006, 2.362829e-006, 
    2.294283e-006, 2.074988e-006, 2.069027e-006, 2.14254e-006, 1.818191e-006, 
    1.318133e-006, 9.161749e-007, 8.712232e-007, 9.423752e-007, 
    8.147224e-007, 7.227072e-007, 6.957614e-007, 6.521752e-007, 
    3.686812e-007, 2.543145e-007, 4.336255e-007, 6.172818e-007, 
    6.121909e-007, 6.17903e-007, 9.96517e-007, 1.168004e-006, 1.114608e-006, 
    8.482496e-007, 6.434832e-007, 4.269198e-007, 2.476093e-007, 
    1.485166e-007, 1.33243e-007, 2.730651e-007, 7.446868e-007, 1.011294e-006, 
    1.215315e-006, 1.357373e-006, 1.329061e-006, 1.121935e-006, 
    1.036874e-006, 9.588914e-007, 9.355458e-007, 7.645551e-007, 
    7.845479e-007, 8.352115e-007, 8.647655e-007, 1.16105e-006, 1.311552e-006, 
    1.173344e-006, 9.148087e-007, 9.504474e-007, 1.193088e-006, 
    1.372523e-006, 1.14379e-006, 1.136463e-006, 1.506012e-006, 1.745052e-006, 
    1.418965e-006, 6.400064e-007, 2.236429e-007, 1.966964e-007, 
    2.122188e-007, -2.842385e-007, -8.206807e-007, -8.188181e-007, 
    -4.140034e-007, -2.503384e-007, -3.054729e-007, -1.298872e-007, 
    5.650168e-008, 2.873453e-007, 5.199279e-007, 9.463492e-007, 
    1.470621e-006, 1.807884e-006, 1.559532e-006, 1.254182e-006, 
    9.924197e-007, 4.692647e-007, 6.239889e-007,
  1.375007e-006, 1.501543e-006, 1.389162e-006, 1.43697e-006, 1.370908e-006, 
    1.345079e-006, 1.385312e-006, 1.419957e-006, 1.368051e-006, 
    1.202525e-006, 1.063323e-006, 9.971377e-007, 9.506948e-007, 
    9.510677e-007, 9.623677e-007, 1.122307e-006, 1.349052e-006, 
    1.446408e-006, 1.565741e-006, 1.635776e-006, 1.563133e-006, 
    1.499555e-006, 1.532089e-006, 1.612059e-006, 1.631679e-006, 
    1.404436e-006, 1.060964e-006, 8.349625e-007, 7.410854e-007, 
    6.290791e-007, 4.524998e-007, 4.110252e-007, 4.187239e-007, 
    3.407415e-007, 3.551459e-007, 5.096213e-007, 5.582983e-007, 
    4.895046e-007, 4.505134e-007, 4.790741e-007, 6.511825e-007, 
    7.332631e-007, 7.02343e-007, 7.279232e-007, 8.624063e-007, 9.280955e-007, 
    8.86248e-007, 8.348388e-007, 7.418309e-007, 6.30569e-007, 6.3417e-007, 
    7.290409e-007, 9.202724e-007, 1.171605e-006, 1.268462e-006, 
    1.276783e-006, 1.303481e-006, 1.357373e-006, 1.438584e-006, 
    1.524142e-006, 1.526253e-006, 1.40754e-006, 1.337505e-006, 1.275293e-006, 
    1.085055e-006, 8.557006e-007, 7.90011e-007, 9.515645e-007, 1.039233e-006, 
    1.026071e-006, 1.01179e-006, 9.541725e-007, 7.320207e-007, 5.130978e-007, 
    2.792738e-007, 7.748736e-008, 1.401968e-007, 2.738102e-007, 
    4.142537e-007, 4.924848e-007, 4.949686e-007, 4.169854e-007, 
    4.027054e-007, 3.860655e-007, 2.55184e-007, 1.558426e-007, 1.924748e-007, 
    3.324215e-007, 5.279994e-007, 7.150088e-007, 6.049881e-007, 
    3.875562e-007, 2.652419e-007, 4.084172e-007, 6.37523e-007, 9.667156e-007,
  1.018991e-006, 1.070774e-006, 1.006326e-006, 9.082273e-007, 8.522236e-007, 
    8.484988e-007, 8.648897e-007, 8.73458e-007, 8.723403e-007, 8.5123e-007, 
    8.030497e-007, 7.845474e-007, 8.802879e-007, 1.059474e-006, 
    1.207492e-006, 1.311552e-006, 1.386928e-006, 1.429644e-006, 
    1.479314e-006, 1.522776e-006, 1.542644e-006, 1.579276e-006, 
    1.552702e-006, 1.418467e-006, 1.193088e-006, 9.261087e-007, 
    7.292892e-007, 6.693119e-007, 7.38851e-007, 8.436557e-007, 8.835159e-007, 
    8.375707e-007, 7.49654e-007, 7.270542e-007, 8.277611e-007, 9.862104e-007, 
    1.116347e-006, 1.200662e-006, 1.268587e-006, 1.376123e-006, 
    1.524018e-006, 1.692898e-006, 1.804036e-006, 1.818316e-006, 
    1.756724e-006, 1.667442e-006, 1.5455e-006, 1.370536e-006, 1.18005e-006, 
    9.97386e-007, 8.519755e-007, 7.927435e-007, 8.194413e-007, 9.689497e-007, 
    1.148757e-006, 1.320741e-006, 1.512469e-006, 1.706557e-006, 
    1.811982e-006, 1.825145e-006, 1.752751e-006, 1.633789e-006, 
    1.502907e-006, 1.438584e-006, 1.458825e-006, 1.502162e-006, 
    1.544009e-006, 1.62845e-006, 1.696126e-006, 1.694139e-006, 1.643724e-006, 
    1.507999e-006, 1.329682e-006, 1.157325e-006, 9.703151e-007, 
    8.093828e-007, 7.032118e-007, 6.719195e-007, 7.157535e-007, 
    7.268052e-007, 7.350009e-007, 7.096689e-007, 6.146743e-007, 
    5.010529e-007, 3.992284e-007, 3.211214e-007, 2.67353e-007, 2.682223e-007, 
    2.99018e-007, 3.129255e-007, 3.04854e-007, 2.534453e-007, 1.917297e-007, 
    2.135848e-007, 4.117696e-007, 7.588428e-007,
  6.145497e-007, 6.982445e-007, 7.862855e-007, 8.620332e-007, 9.175392e-007, 
    9.544196e-007, 9.869545e-007, 1.012659e-006, 1.035507e-006, 
    1.055748e-006, 1.076858e-006, 1.096976e-006, 1.112994e-006, 
    1.123425e-006, 1.126653e-006, 1.124791e-006, 1.11498e-006, 1.09474e-006, 
    1.064192e-006, 1.026071e-006, 9.843475e-007, 9.499504e-007, 
    9.253633e-007, 9.031357e-007, 8.831435e-007, 8.632753e-007, 
    8.478773e-007, 8.26519e-007, 7.937365e-007, 7.574768e-007, 7.261845e-007, 
    6.945195e-007, 6.705536e-007, 6.638479e-007, 6.75396e-007, 7.013489e-007, 
    7.350009e-007, 7.77469e-007, 8.292507e-007, 8.74575e-007, 9.077303e-007, 
    9.293367e-007, 9.424995e-007, 9.508193e-007, 9.55911e-007, 9.628648e-007, 
    9.644791e-007, 9.663418e-007, 9.757794e-007, 9.98255e-007, 1.034142e-006, 
    1.073879e-006, 1.100204e-006, 1.115974e-006, 1.121811e-006, 
    1.125784e-006, 1.132862e-006, 1.139319e-006, 1.144162e-006, 
    1.142796e-006, 1.133483e-006, 1.124294e-006, 1.124294e-006, 1.13311e-006, 
    1.158442e-006, 1.197682e-006, 1.246608e-006, 1.292181e-006, 1.32993e-006, 
    1.338126e-006, 1.316643e-006, 1.268835e-006, 1.204636e-006, 
    1.136463e-006, 1.077852e-006, 1.03377e-006, 1.001981e-006, 9.844716e-007, 
    9.755308e-007, 9.744128e-007, 9.793798e-007, 9.876997e-007, 1.00136e-006, 
    1.018992e-006, 1.033397e-006, 1.030789e-006, 1.012412e-006, 
    9.791315e-007, 9.244945e-007, 8.4974e-007, 7.619478e-007, 6.71298e-007, 
    5.895899e-007, 5.345801e-007, 5.211691e-007, 5.519646e-007,
  3.777177e-007, 3.650514e-007, 3.667901e-007, 3.748614e-007, 3.829327e-007, 
    3.93115e-007, 4.006902e-007, 3.995722e-007, 3.880239e-007, 3.671621e-007, 
    3.436927e-007, 3.141388e-007, 2.842123e-007, 2.59377e-007, 2.437308e-007, 
    2.380187e-007, 2.388878e-007, 2.433583e-007, 2.457176e-007, 
    2.478287e-007, 2.455935e-007, 2.409989e-007, 2.401296e-007, 
    2.432341e-007, 2.544099e-007, 2.7403e-007, 3.007278e-007, 3.345037e-007, 
    3.717566e-007, 4.081403e-007, 4.415438e-007, 4.672485e-007, 
    4.841365e-007, 4.886067e-007, 4.827705e-007, 4.677452e-007, 
    4.494912e-007, 4.298715e-007, 4.143496e-007, 4.107485e-007, 
    4.214278e-007, 4.534652e-007, 5.068612e-007, 5.764e-007, 6.58853e-007, 
    7.507435e-007, 8.50333e-007, 9.545165e-007, 1.054106e-006, 1.141402e-006, 
    1.209947e-006, 1.24571e-006, 1.252416e-006, 1.236893e-006, 1.212306e-006, 
    1.182504e-006, 1.145375e-006, 1.100299e-006, 1.050008e-006, 
    1.005428e-006, 9.640771e-007, 9.276937e-007, 8.940419e-007, 
    8.616316e-007, 8.417642e-007, 8.355551e-007, 8.400257e-007, 
    8.458624e-007, 8.453658e-007, 8.304651e-007, 7.997933e-007, 
    7.606775e-007, 7.151048e-007, 6.706491e-007, 6.31037e-007, 6.068233e-007, 
    6.07444e-007, 6.284299e-007, 6.663033e-007, 7.15105e-007, 7.689973e-007, 
    8.246286e-007, 8.780244e-007, 9.229761e-007, 9.545167e-007, 
    9.669341e-007, 9.608495e-007, 9.368837e-007, 8.879581e-007, 
    8.237589e-007, 7.483839e-007, 6.66055e-007, 5.890656e-007, 5.167949e-007, 
    4.544586e-007, 4.076439e-007,
  6.615937e-008, 1.61775e-007, 2.719194e-007, 3.803254e-007, 4.640199e-007, 
    5.094687e-007, 5.273498e-007, 5.160495e-007, 4.951877e-007, 
    4.669997e-007, 4.126105e-007, 3.358695e-007, 2.595009e-007, 
    2.078436e-007, 1.806491e-007, 1.681071e-007, 1.682314e-007, 
    1.727017e-007, 1.871063e-007, 2.309405e-007, 2.924075e-007, 
    3.541232e-007, 3.944806e-007, 4.174534e-007, 4.230412e-007, 
    4.044148e-007, 3.780895e-007, 3.779652e-007, 3.874027e-007, 
    3.821873e-007, 3.72129e-007, 3.716324e-007, 3.670377e-007, 3.420784e-007, 
    2.896759e-007, 2.239866e-007, 1.510949e-007, 7.298831e-008, 
    3.946184e-009, -5.044285e-008, -6.795176e-008, -6.670962e-008, 
    -8.384563e-008, -1.790888e-007, -3.047555e-007, -4.366307e-007, 
    -5.523639e-007, -5.947086e-007, -5.940879e-007, -5.79435e-007, 
    -5.084057e-007, -4.690401e-007, -5.472739e-007, -7.968674e-007, 
    -1.139592e-006, -1.494862e-006, -1.756253e-006, -1.822937e-006, 
    -1.735269e-006, -1.575204e-006, -1.333432e-006, -1.053912e-006, 
    -7.458311e-007, -4.343956e-007, -1.143935e-007, 2.381425e-007, 
    5.535503e-007, 7.107574e-007, 7.103854e-007, 6.029732e-007, 
    4.629023e-007, 3.362429e-007, 2.837164e-007, 3.074342e-007, 
    4.142257e-007, 5.831048e-007, 7.684998e-007, 9.309233e-007, 1.03548e-006, 
    1.070498e-006, 1.03548e-006, 8.978914e-007, 6.541336e-007, 4.104991e-007, 
    1.934395e-007, 1.73568e-008, -1.337644e-007, -2.275183e-007, 
    -2.565753e-007, -2.824036e-007, -3.067421e-007, -3.006576e-007, 
    -2.607967e-007, -1.66423e-007, -7.018616e-008, 1.463377e-009,
  7.517367e-007, 6.469315e-007, 4.907176e-007, 3.388499e-007, 2.455934e-007, 
    1.7146e-007, 1.471215e-007, 1.970403e-007, 2.104514e-007, 1.626437e-007, 
    1.720807e-007, 2.236141e-007, 2.428613e-007, 2.814801e-007, 
    3.266803e-007, 3.666652e-007, 4.004411e-007, 4.219237e-007, 
    4.108718e-007, 3.943564e-007, 3.703905e-007, 3.499014e-007, 
    3.126485e-007, 2.678207e-007, 2.478283e-007, 2.784998e-007, 
    2.945186e-007, 3.042046e-007, 3.138902e-007, 3.075573e-007, 
    3.246936e-007, 3.261836e-007, 3.019692e-007, 2.883098e-007, 
    3.223341e-007, 3.536267e-007, 3.89762e-007, 3.744883e-007, 3.012248e-007, 
    1.933154e-007, 1.23777e-007, 1.143401e-007, 6.927166e-009, 
    -1.389808e-007, -1.152634e-007, 7.522294e-008, 7.90742e-008, 
    -2.117476e-007, -5.943348e-007, -8.289053e-007, -9.956739e-007, 
    -1.173868e-006, -1.089673e-006, -9.554387e-007, -9.350742e-007, 
    -9.90829e-007, -1.091164e-006, -1.177963e-006, -1.337902e-006, 
    -1.545774e-006, -1.907996e-006, -2.071536e-006, -1.785683e-006, 
    -1.256692e-006, -4.932544e-007, 4.98168e-007, 1.444888e-006, 
    2.067881e-006, 2.214037e-006, 2.164366e-006, 2.06192e-006, 2.030504e-006, 
    2.173431e-006, 2.345291e-006, 2.467231e-006, 2.520504e-006, 
    2.586069e-006, 2.519014e-006, 2.298353e-006, 2.053352e-006, 
    1.793701e-006, 1.40776e-006, 1.01201e-006, 7.200715e-007, 5.328138e-007, 
    3.279224e-007, 1.040326e-007, 8.913503e-009, 1.265075e-007, 
    3.325163e-007, 5.494526e-007, 8.600182e-007, 1.096947e-006, 
    1.042185e-006, 9.177604e-007, 8.298437e-007,
  5.689494e-007, 5.602567e-007, 6.556238e-007, 6.825701e-007, 5.586423e-007, 
    4.3161e-007, 4.167089e-007, 5.321926e-007, 6.627021e-007, 7.102612e-007, 
    6.466831e-007, 4.583073e-007, 2.160392e-007, 1.314752e-007, 
    4.194396e-008, 3.94607e-009, 1.646303e-007, 4.501118e-007, 5.766476e-007, 
    6.063257e-007, 6.572379e-007, 6.514017e-007, 5.520607e-007, 
    4.927042e-007, 5.388978e-007, 6.280567e-007, 6.802106e-007, 
    6.743742e-007, 7.388218e-007, 7.616702e-007, 7.223063e-007, 
    6.089333e-007, 5.205197e-007, 4.913383e-007, 4.580589e-007, 
    4.612875e-007, 4.766854e-007, 4.539611e-007, 5.797518e-007, 
    8.009102e-007, 1.058452e-006, 1.236149e-006, 1.217274e-006, 
    8.914344e-007, 8.263655e-007, 1.127866e-006, 1.452589e-006, 
    1.187844e-006, 6.507817e-007, 2.443721e-008, -8.000952e-007, 
    -1.312695e-006, -1.66014e-006, -1.911473e-006, -1.828523e-006, 
    -1.876952e-006, -1.831503e-006, -1.786057e-006, -2.05204e-006, 
    -1.746319e-006, -4.074518e-007, 1.59961e-006, 3.422023e-006, 
    4.347141e-006, 4.76909e-006, 5.490057e-006, 6.732318e-006, 7.592487e-006, 
    7.416033e-006, 6.224558e-006, 5.083752e-006, 4.342294e-006, 
    4.271516e-006, 4.568792e-006, 4.794793e-006, 4.895005e-006, 
    5.284545e-006, 5.472176e-006, 5.41642e-006, 4.556995e-006, 3.376823e-006, 
    2.677712e-006, 2.317352e-006, 2.00803e-006, 1.758559e-006, 1.645932e-006, 
    1.673375e-006, 2.452954e-006, 3.672861e-006, 4.113934e-006, 
    3.605681e-006, 2.753956e-006, 2.093585e-006, 1.48835e-006, 9.961154e-007, 
    7.34849e-007,
  1.788609e-006, 1.290288e-006, 1.008284e-006, 1.048766e-006, 8.34686e-007, 
    7.086469e-007, 7.601798e-007, 7.391945e-007, 6.889031e-007, 
    8.151901e-007, 1.084777e-006, 1.149597e-006, 1.224724e-006, 
    8.661036e-007, 2.915394e-007, 2.598742e-007, 4.391845e-007, 
    6.952366e-007, 7.341034e-007, 8.718152e-007, 1.017226e-006, 
    1.149722e-006, 1.259618e-006, 1.282963e-006, 1.311896e-006, 
    1.357469e-006, 1.310158e-006, 1.031258e-006, 6.346384e-007, 
    5.626164e-007, 7.642786e-007, 7.872513e-007, 7.415545e-007, 
    5.936604e-007, 7.182095e-007, 1.141402e-006, 1.48475e-006, 1.329902e-006, 
    8.79018e-007, 7.000795e-007, 8.146944e-007, 8.770303e-007, 8.3332e-007, 
    7.182084e-007, 4.794174e-007, 6.92753e-007, 1.267319e-006, 1.14202e-006, 
    8.571606e-007, 1.014741e-006, 1.083165e-006, 3.307805e-007, -7.8011e-008, 
    3.265577e-007, 2.058368e-008, -5.197107e-007, -5.902402e-007, 
    -7.909093e-007, -9.478663e-007, -1.052544e-006, -2.816614e-007, 
    1.789973e-006, 2.944069e-006, 3.206331e-006, 4.569662e-006, 
    4.765488e-006, 3.719424e-006, 3.972498e-006, 5.487947e-006, 
    5.983533e-006, 5.608274e-006, 5.464972e-006, 5.402886e-006, 
    4.689616e-006, 4.416676e-006, 4.531914e-006, 4.862968e-006, 
    4.449586e-006, 4.241714e-006, 3.215396e-006, 1.92421e-006, 1.532434e-006, 
    1.497292e-006, 2.067384e-006, 3.010877e-006, 4.103628e-006, 3.83727e-006, 
    2.88521e-006, 3.952879e-006, 4.881843e-006, 4.474665e-006, 4.092201e-006, 
    3.857509e-006, 3.19205e-006, 2.785497e-006, 2.281094e-006,
  3.750844e-006, 3.492431e-006, 3.378686e-006, 3.869056e-006, 3.864092e-006, 
    3.405758e-006, 4.056812e-006, 3.106736e-006, 1.540624e-006, 
    5.796282e-007, -7.093149e-008, 1.289543e-006, 4.856511e-006, 
    6.106343e-006, 4.136162e-006, 2.405518e-006, 1.176047e-006, 
    5.329371e-007, 9.507908e-007, 1.698209e-006, 1.827477e-006, 
    2.338337e-006, 3.607294e-006, 4.468333e-006, 4.155037e-006, 
    3.531052e-006, 3.06862e-006, 3.087494e-006, 2.649028e-006, 2.033486e-006, 
    1.76812e-006, 1.06727e-006, 7.336075e-007, 6.250775e-007, 1.249063e-006, 
    1.93936e-006, 3.132692e-006, 2.850935e-006, 1.205352e-006, 3.57104e-007, 
    5.010243e-007, 1.131839e-006, 1.33201e-006, 9.819596e-007, 
    -9.278847e-008, -6.646223e-008, 1.841507e-006, 1.900735e-006, 
    1.043918e-006, 1.808476e-006, 2.591783e-006, 2.023055e-006, 
    2.351626e-006, 3.136916e-006, 3.66566e-006, 3.109721e-006, 1.917873e-006, 
    1.634751e-006, 2.326908e-006, 3.732961e-006, 3.945674e-006, 
    3.061543e-006, 2.901725e-006, 3.667521e-006, 3.252273e-006, 
    3.414698e-006, 3.982928e-006, 4.696818e-006, 5.20594e-006, 5.617587e-006, 
    5.249896e-006, 3.900597e-006, 3.317837e-006, 3.893643e-006, 
    5.457026e-006, 6.050839e-006, 5.730583e-006, 5.368487e-006, 
    5.098407e-006, 3.805731e-006, 1.666671e-006, 2.131335e-006, 
    2.778539e-006, 2.560738e-006, 2.410608e-006, 2.57303e-006, 2.697827e-006, 
    2.669143e-006, 2.956984e-006, 3.727002e-006, 4.493913e-006, 
    4.314599e-006, 2.206212e-006, 1.788731e-006, 2.501874e-006, 3.080166e-006,
  4.837015e-006, 5.687372e-006, 7.497983e-006, 7.614592e-006, 7.936336e-006, 
    7.157247e-006, 7.219583e-006, 6.865557e-006, 6.464466e-006, 
    6.737529e-006, 7.30688e-006, 6.320795e-006, 7.39083e-006, 1.0492e-005, 
    1.009911e-005, 8.975438e-006, 7.409946e-006, 6.721757e-006, 
    7.155755e-006, 6.029852e-006, 5.488073e-006, 4.896865e-006, 
    4.183474e-006, 4.094691e-006, 4.38427e-006, 5.558109e-006, 6.000051e-006, 
    5.453299e-006, 4.422509e-006, 3.199246e-006, 2.321074e-006, 
    1.067639e-006, 4.001886e-007, 1.255888e-006, 2.786863e-006, 
    5.348622e-006, 6.951243e-006, 6.611997e-006, 6.909893e-006, 
    8.388462e-006, 1.055086e-005, 9.232606e-006, 5.841106e-006, 
    4.151563e-006, 3.686524e-006, 4.311372e-006, 5.38128e-006, 4.724261e-006, 
    4.519739e-006, 4.07991e-006, 4.475287e-006, 4.61188e-006, 4.068361e-006, 
    3.638086e-006, 4.164222e-006, 3.140138e-006, 2.937244e-006, 
    4.009376e-006, 4.598593e-006, 5.851531e-006, 5.589394e-006, 
    4.557367e-006, 3.893649e-006, 4.123865e-006, 5.049478e-006, 
    6.330107e-006, 6.022025e-006, 5.335205e-006, 6.089827e-006, 
    6.587898e-006, 6.511533e-006, 4.943931e-006, 3.699928e-006, 
    4.439151e-006, 7.196735e-006, 8.08671e-006, 7.271115e-006, 7.27298e-006, 
    6.696057e-006, 5.217489e-006, 4.31063e-006, 3.22595e-006, 2.362178e-006, 
    2.756064e-006, 3.142746e-006, 3.250783e-006, 3.722902e-006, 
    3.452071e-006, 2.657342e-006, 2.701796e-006, 3.150819e-006, 
    3.979201e-006, 3.469702e-006, 3.904071e-006, 4.464231e-006, 5.372585e-006,
  5.361408e-006, 3.518007e-006, 3.881722e-006, 3.809699e-006, 4.249905e-006, 
    6.432925e-006, 5.799009e-006, 5.445851e-006, 7.264787e-006, 
    6.070704e-006, 4.807582e-006, 3.310883e-006, 4.160011e-006, 6.97732e-006, 
    7.623905e-006, 8.292096e-006, 9.449668e-006, 9.282405e-006, 
    8.357785e-006, 6.981039e-006, 6.594353e-006, 6.172651e-006, 
    7.005627e-006, 7.248265e-006, 6.906659e-006, 6.16632e-006, 5.995948e-006, 
    5.46199e-006, 3.739047e-006, 3.100409e-006, 2.620471e-006, 4.218989e-006, 
    4.659814e-006, 5.459504e-006, 5.251637e-006, 6.898459e-006, 
    8.982272e-006, 8.465202e-006, 9.839961e-006, 8.381881e-006, 9.57695e-006, 
    9.167041e-006, 7.09193e-006, 6.183582e-006, 5.272377e-006, 5.080894e-006, 
    3.277975e-006, 3.053467e-006, 3.775678e-006, 7.084109e-006, 
    8.970224e-006, 7.044993e-006, 6.370838e-006, 6.492533e-006, 
    6.434539e-006, 5.307642e-006, 3.669751e-006, 3.455301e-006, 
    3.486966e-006, 4.034089e-006, 4.21874e-006, 4.892276e-006, 7.740751e-006, 
    7.312592e-006, 7.00575e-006, 5.510916e-006, 6.187804e-006, 8.263038e-006, 
    6.423366e-006, 4.607911e-006, 4.121137e-006, 5.498001e-006, 6.64775e-006, 
    7.456885e-006, 6.587774e-006, 5.614727e-006, 3.625546e-006, 
    1.613271e-006, 1.853799e-006, 3.272515e-006, 4.56668e-006, 5.247046e-006, 
    4.999314e-006, 4.295476e-006, 4.452559e-006, 3.771453e-006, 
    3.404763e-006, 3.99125e-006, 4.886808e-006, 5.113554e-006, 5.094056e-006, 
    6.356684e-006, 8.266763e-006, 7.740131e-006, 6.695438e-006, 6.65185e-006,
  5.423868e-006, 4.200236e-006, 2.931154e-006, 3.733707e-006, 4.968017e-006, 
    4.76487e-006, 3.897869e-006, 4.425619e-006, 5.270264e-006, 4.61896e-006, 
    6.716669e-006, 6.51327e-006, 5.696063e-006, 5.723137e-006, 5.580707e-006, 
    6.150418e-006, 6.276212e-006, 5.291862e-006, 4.986898e-006, 
    6.810051e-006, 7.032822e-006, 7.901188e-006, 7.993829e-006, 
    7.444341e-006, 7.110066e-006, 6.541712e-006, 6.254118e-006, 
    6.450318e-006, 6.703016e-006, 6.840728e-006, 7.573119e-006, 
    6.897846e-006, 6.560214e-006, 7.259823e-006, 7.93708e-006, 8.991461e-006, 
    7.668241e-006, 7.055176e-006, 8.388961e-006, 7.455401e-006, 
    6.187558e-006, 7.896597e-006, 7.584793e-006, 6.554499e-006, 
    7.809547e-006, 8.634821e-006, 1.070584e-005, 8.010218e-006, 
    5.805217e-006, 6.616954e-006, 7.533134e-006, 5.439148e-006, 
    6.038668e-006, 7.213872e-006, 5.199112e-006, 2.395207e-006, 
    1.921471e-006, 5.121752e-006, 6.93833e-006, 5.079402e-006, 3.849564e-006, 
    3.30952e-006, 6.108949e-006, 6.131053e-006, 5.01409e-006, 6.398157e-006, 
    8.21076e-006, 9.472764e-006, 8.337793e-006, 7.916589e-006, 7.237715e-006, 
    9.05553e-006, 1.203415e-005, 1.008868e-005, 5.893016e-006, 3.807592e-006, 
    3.00206e-006, 2.755572e-006, 2.037708e-006, 1.16288e-006, 2.571292e-006, 
    3.996462e-006, 3.062903e-006, 1.67213e-006, 4.323574e-007, 4.633966e-007, 
    8.477255e-007, 1.258501e-006, 1.882854e-006, 2.44376e-006, 3.422025e-006, 
    5.342657e-006, 6.4333e-006, 5.114174e-006, 3.540235e-006, 5.43753e-006,
  3.998208e-006, 4.337209e-006, 5.161615e-006, 7.089329e-006, 8.009101e-006, 
    6.160364e-006, 4.955717e-006, 4.407604e-006, 4.098907e-006, 
    4.720037e-006, 5.9839e-006, 7.85747e-006, 6.156381e-006, 5.69606e-006, 
    6.747214e-006, 6.934351e-006, 8.485193e-006, 9.895339e-006, 
    1.036385e-005, 8.788549e-006, 7.023267e-006, 6.408347e-006, 
    5.643913e-006, 6.610004e-006, 9.312211e-006, 9.645002e-006, 
    8.172516e-006, 9.374049e-006, 9.217216e-006, 6.894617e-006, 
    8.011826e-006, 8.272098e-006, 8.06621e-006, 7.432416e-006, 6.410941e-006, 
    5.686124e-006, 4.44461e-006, 5.695318e-006, 6.563565e-006, 7.379156e-006, 
    8.579311e-006, 7.849159e-006, 4.874266e-006, 4.234138e-006, 
    3.684287e-006, 5.652353e-006, 5.563195e-006, 7.164206e-006, 
    6.145834e-006, 5.969499e-006, 6.030721e-006, 7.802217e-006, 
    6.779632e-006, 4.556623e-006, 9.782307e-007, -1.066452e-006, 
    1.284823e-006, 3.066263e-006, 3.656591e-006, 2.196526e-006, 
    1.698209e-006, 4.788955e-006, 5.923306e-006, 7.29881e-006, 6.927523e-006, 
    7.303279e-006, 9.001265e-006, 8.260558e-006, 7.230392e-006, 
    6.014205e-006, 9.956184e-006, 1.012718e-005, 7.679904e-006, 
    3.684283e-006, 2.891789e-006, 2.863595e-006, 2.784494e-006, 
    2.458793e-006, 3.719922e-006, 7.678773e-007, -9.822634e-007, 
    -3.524419e-007, -1.296556e-006, -1.201188e-006, -7.567578e-007, 
    7.95575e-007, 4.416725e-007, -1.329208e-006, 3.897621e-007, 
    2.587438e-006, 3.422025e-006, 3.15778e-006, 3.317469e-006, 3.239238e-006, 
    1.942215e-006, 1.59601e-006,
  3.766356e-006, 4.078785e-006, 3.650748e-006, 5.436159e-006, 3.387988e-006, 
    1.167591e-006, 1.667777e-006, 1.509452e-006, 2.500008e-006, 
    3.895006e-006, 7.783958e-006, 5.555488e-006, 3.965044e-006, 
    4.499005e-006, 4.933874e-006, 4.797774e-006, 4.158017e-006, 
    5.394693e-006, 4.615486e-006, 4.492184e-006, 4.098787e-006, 4.96467e-006, 
    5.710346e-006, 8.602281e-006, 8.946005e-006, 7.143586e-006, 
    6.783102e-006, 6.914106e-006, 7.465445e-006, 8.627489e-006, 
    9.099607e-006, 6.957442e-006, 4.680296e-006, 4.178997e-006, 
    4.044519e-006, 5.833652e-006, 4.239715e-006, 2.777793e-006, 
    1.316614e-006, 1.793574e-006, 8.470997e-007, 1.469474e-006, 
    -6.934279e-007, 4.74829e-007, 8.295327e-006, 7.925904e-006, 
    5.548298e-006, 5.22047e-006, 3.898615e-006, 1.167107e-006, 2.044162e-006, 
    3.70303e-006, 2.181372e-006, -1.044646e-007, -8.827992e-007, 
    1.169337e-006, 2.440782e-006, 1.719811e-006, 4.507274e-007, 
    1.492324e-006, 3.10798e-006, 2.870307e-006, 3.213161e-006, 1.773082e-006, 
    2.289489e-007, 1.127228e-007, 4.440768e-006, 4.185698e-006, 
    5.196616e-006, 1.114479e-005, 1.188463e-005, 8.18877e-006, 3.867062e-006, 
    3.175152e-006, 3.526078e-006, 1.570665e-006, 5.034963e-007, 
    1.195665e-006, 3.201485e-006, 6.964747e-007, -2.571353e-006, 
    -2.602395e-006, -1.356279e-006, -6.851042e-007, -4.889062e-007, 
    -1.231114e-006, 4.840149e-007, 2.349389e-006, 3.926427e-006, 
    5.030233e-006, 2.21291e-006, -1.173499e-006, -1.51759e-006, 
    -1.718137e-006, 3.162459e-007, 1.470587e-006,
  7.086419e-007, 2.659817e-006, 3.004283e-006, -6.24641e-009, 1.207456e-006, 
    2.511431e-006, 1.111093e-006, 4.786671e-007, 1.890432e-006, 
    8.366769e-007, -1.225151e-006, -9.214127e-007, 1.542616e-006, 
    2.554036e-006, 3.215273e-006, 1.86312e-006, 1.347289e-006, 2.886456e-006, 
    4.505344e-006, 3.911406e-006, 4.475292e-006, 4.849924e-006, 
    5.874623e-006, 5.078156e-006, 2.869678e-006, 5.930306e-007, 
    3.457899e-007, 2.754321e-006, 4.089463e-006, 5.096659e-006, 
    3.540728e-006, -3.036439e-007, -3.03764e-007, 2.691741e-008, 
    -1.656666e-006, -2.892968e-006, -3.633057e-006, -4.738475e-006, 
    -4.740585e-006, -5.542766e-006, -5.023086e-006, -2.412777e-006, 
    -1.434761e-006, 8.714778e-008, 2.622703e-006, 3.874276e-006, 
    -1.076514e-006, 2.352826e-007, 1.503005e-006, 4.64639e-007, 
    4.322283e-007, 1.954253e-006, 4.483227e-006, 2.01162e-006, 2.092456e-006, 
    2.569919e-006, -2.23397e-006, -5.614045e-006, -4.797083e-006, 
    -2.619407e-006, -2.224533e-006, 8.172901e-007, -4.31919e-007, 
    -1.093402e-006, -4.425929e-007, 2.008641e-006, 1.520002e-006, 
    3.856258e-006, 4.033824e-006, 3.040295e-006, 2.681798e-006, 
    9.885298e-007, 6.743649e-007, 1.266562e-006, -1.260047e-006, 
    -2.338154e-006, -1.679895e-006, -3.199686e-006, -1.910237e-006, 
    -1.270599e-006, -2.58575e-006, -3.779705e-006, -4.60362e-006, 
    -3.090652e-006, -1.048447e-006, 8.466013e-007, 3.078418e-006, 
    3.757541e-006, 1.680444e-006, 3.44553e-007, -8.423231e-007, 
    -2.004563e-007, 1.865465e-006, 1.795303e-006, 2.657212e-006, 2.178389e-006,
  1.349435e-007, -1.112407e-006, -2.52268e-006, -3.412155e-006, 
    -1.450782e-006, -1.877452e-006, -4.321555e-007, 2.194289e-006, 
    2.313374e-006, 3.69484e-006, 3.874149e-006, 4.191299e-006, 2.358331e-006, 
    2.688892e-006, 2.288914e-006, 2.049259e-006, 2.962695e-006, 
    1.989772e-006, 2.856279e-006, 2.477667e-006, 2.428122e-006, 
    1.950662e-006, 1.08379e-007, -3.169505e-006, -7.974882e-006, 
    -6.039721e-006, -1.313445e-006, -5.478796e-008, 8.358074e-007, 
    5.60256e-007, -3.709676e-006, -2.855963e-006, -3.429534e-006, 
    -2.79089e-006, -2.672554e-006, -3.31194e-006, -5.737598e-006, 
    -7.421433e-006, -7.59503e-006, -2.341625e-006, -1.014554e-006, 
    -2.477846e-006, -5.455386e-007, -7.131712e-007, 1.229091e-007, 
    -1.550619e-006, 3.399655e-007, 2.793076e-006, 2.123386e-006, 
    -4.486828e-007, 5.772563e-007, 5.376532e-007, 1.66666e-006, 
    4.601192e-006, 1.921104e-006, -1.354303e-006, 4.334652e-007, 
    -1.852968e-007, -1.248503e-006, -1.838464e-006, -5.185888e-006, 
    -4.621877e-006, -5.58524e-006, -7.965198e-006, -4.363217e-006, 
    -1.239572e-006, 1.002318e-006, -3.292447e-006, -4.897549e-006, 
    -2.516972e-006, -2.806923e-006, -2.964996e-006, -1.922635e-007, 
    -4.332676e-006, -6.767266e-006, -1.07809e-005, -1.547017e-005, 
    -1.379652e-005, -6.412616e-006, -4.751635e-006, -2.69962e-006, 
    -7.580002e-007, 1.175173e-006, 2.024921e-006, 1.467612e-006, 
    7.553353e-007, -1.653098e-007, -5.219445e-007, 1.147724e-006, 
    2.515775e-006, 2.850804e-006, 2.903333e-006, -3.928035e-007, 
    -1.150656e-006, -1.645371e-006, -1.642638e-006,
  -3.372537e-006, -6.514078e-006, -7.768007e-006, -7.785136e-006, 
    -7.141907e-006, -4.541776e-006, -1.704471e-006, 4.049089e-007, 
    3.613008e-006, 6.758019e-006, 3.403769e-006, -1.980396e-006, 
    -4.55718e-006, -4.150501e-006, -3.089035e-006, -3.088295e-006, 
    -8.125171e-007, -1.283141e-006, -3.083951e-006, -5.454785e-008, 
    1.482367e-007, -4.478947e-006, -4.754491e-006, -3.892708e-006, 
    -1.918059e-006, 1.911416e-006, 3.936982e-006, 2.706272e-006, 
    -9.226569e-007, -2.971692e-006, -4.894686e-006, -5.856935e-006, 
    -5.767153e-006, -6.320237e-006, -5.583986e-006, -4.149508e-006, 
    -3.753754e-006, -2.823675e-006, -3.164912e-006, -3.087056e-006, 
    -2.488519e-006, 1.942091e-006, 4.925303e-006, 3.330755e-006, 
    3.827954e-006, 2.997589e-006, 2.715457e-006, 6.300979e-009, 
    -6.572991e-007, -1.071185e-006, -6.738097e-006, -3.441575e-006, 
    -2.084835e-006, -8.70139e-007, -5.231701e-006, -7.516555e-006, 
    -3.01516e-006, -6.490976e-006, -5.524889e-006, -3.113135e-006, 
    2.828823e-006, -1.735407e-006, -5.06072e-006, -1.153887e-006, 
    3.016583e-006, 1.322314e-006, 7.818999e-007, -7.057351e-007, 
    -3.476089e-007, -2.857705e-007, -1.408323e-006, -3.593574e-006, 
    -4.827889e-006, -7.379836e-006, -6.062197e-006, -8.673254e-006, 
    -1.720107e-005, -1.676396e-005, -5.925722e-006, 2.091969e-006, 
    4.066991e-006, 6.57374e-006, 7.160976e-006, 6.020284e-006, 4.718542e-006, 
    4.466463e-006, 1.826978e-006, 2.254761e-006, 3.659694e-006, 
    3.142501e-006, 1.27067e-006, -1.576704e-006, -1.348588e-006, 
    -2.24253e-006, -2.56328e-006, -2.150766e-006,
  -4.097103e-006, -4.827503e-006, -6.059587e-006, -5.640119e-006, 
    -6.151224e-006, -3.974043e-006, -1.944383e-006, -7.481922e-007, 
    -1.870994e-006, -5.195943e-006, -1.288234e-005, -1.094816e-005, 
    -1.0426e-005, -6.161785e-006, -6.641225e-006, -5.311049e-006, 
    -2.814986e-006, -6.794338e-006, -2.813988e-006, -3.513269e-007, 
    8.550523e-007, 7.386934e-007, 3.417554e-006, 4.731462e-006, 
    5.596105e-006, 3.283694e-006, -9.424057e-007, -3.275305e-006, 
    -6.272303e-006, -8.981331e-006, -9.667287e-006, -9.191936e-006, 
    -6.532573e-006, -5.650425e-006, -3.084819e-006, -1.943761e-006, 
    -3.758352e-006, -2.828641e-006, 1.943063e-007, 3.730602e-006, 
    4.198995e-006, 3.426614e-006, 7.17687e-006, 1.054962e-005, 5.07183e-006, 
    8.44615e-007, -3.923633e-006, -5.238038e-006, -3.808651e-006, 
    -6.038968e-006, -3.176712e-006, 1.781664e-007, -2.13326e-006, 
    -4.789261e-006, -7.723058e-006, -1.050287e-005, -8.6699e-006, 
    -7.91491e-006, -3.744448e-006, 2.41333e-006, 3.380414e-006, 
    -1.065593e-006, 2.006778e-006, 9.538813e-006, 1.043226e-005, 
    1.087768e-005, 3.848312e-006, 3.719168e-006, 4.647256e-006, 
    2.147844e-006, 7.445233e-007, -3.612196e-006, -4.897047e-006, 
    -5.311917e-006, -6.209833e-006, -7.999719e-006, -9.973621e-006, 
    -8.156797e-006, -2.841306e-006, 3.151568e-006, 6.573247e-006, 
    8.391189e-006, 1.070646e-005, 1.190462e-005, 8.355168e-006, 
    6.102367e-006, 4.625792e-006, 2.759047e-006, -5.503807e-007, 
    -1.250115e-006, 1.058906e-007, 8.793904e-007, 1.059319e-006, 
    1.459171e-006, 1.759303e-006, -2.617415e-006,
  -4.631558e-006, -3.663357e-006, -4.494839e-006, -4.500179e-006, 
    -2.571223e-006, -2.016776e-006, -3.54874e-006, -2.391415e-006, 
    -5.25132e-006, -1.016213e-005, -1.365781e-005, -7.831579e-006, 
    -4.815334e-006, -1.413033e-006, 1.08068e-006, -3.182173e-006, 
    -1.388562e-007, -9.867326e-007, 2.001076e-006, 6.40412e-006, 
    7.622039e-006, 9.097877e-006, 5.297958e-006, 1.110606e-006, 
    -2.249855e-006, -1.366087e-006, -4.522033e-006, -7.440054e-006, 
    -7.760555e-006, -9.792569e-006, -8.644691e-006, -5.445159e-006, 
    -3.790259e-006, 1.021326e-006, -9.162031e-007, -4.673155e-006, 
    -5.485396e-006, 1.945318e-006, 8.512383e-006, 8.528527e-006, 
    6.840843e-006, 4.264806e-006, 5.551776e-006, 6.482725e-006, 
    2.174296e-006, -1.511879e-006, -5.429763e-006, -3.129393e-006, 
    2.210923e-006, 6.866547e-006, 9.536954e-006, 1.654375e-006, 
    -3.073765e-006, -2.204037e-006, -4.149755e-006, -7.32917e-006, 
    -4.960883e-006, 1.465989e-006, 6.012269e-007, 3.7262e-007, 1.125954e-008, 
    1.952511e-006, 4.526813e-006, 5.603175e-006, 6.460858e-006, 
    -5.986913e-007, -4.187132e-006, -9.152172e-007, -2.05962e-006, 
    -1.484805e-006, 1.795936e-006, -2.28265e-007, -3.905619e-006, 
    -7.290919e-006, -6.075978e-006, -5.165144e-006, -4.161426e-006, 
    -3.197195e-006, -1.765939e-006, 4.760397e-006, 8.578198e-006, 
    1.437438e-006, 2.184857e-006, 6.371583e-006, 5.198857e-006, 
    5.538735e-006, 2.558128e-006, 7.098861e-007, 1.948922e-006, 
    4.365756e-007, -1.14282e-006, -8.45419e-007, -6.205355e-007, 
    -1.62674e-006, -2.194845e-006, -4.483665e-006,
  -2.634924e-006, -2.532726e-006, -1.741228e-006, -1.225648e-006, 
    -1.802571e-006, -1.937055e-006, -3.73935e-006, -4.501796e-006, 
    -7.315011e-006, -9.329773e-006, -1.128616e-005, -5.287702e-006, 
    -2.43413e-006, -3.155845e-006, -2.054185e-007, -1.281276e-006, 
    5.790062e-007, 3.924446e-006, 3.298723e-006, 1.035032e-005, 
    5.071834e-006, 1.314729e-007, -2.583642e-006, 3.538735e-007, 
    4.272257e-006, 1.042556e-006, -5.36755e-006, -4.711652e-006, 
    -2.7596e-006, -1.339273e-006, -1.943392e-006, -1.00834e-006, 
    4.128837e-006, 2.720551e-006, -8.614388e-007, 2.769973e-006, 
    6.606899e-006, 8.701506e-006, 7.588513e-006, 2.269545e-006, 
    6.575235e-006, 5.78013e-006, 3.967281e-006, 7.201457e-006, 
    -1.083343e-006, -6.883995e-006, -6.003214e-006, 1.218636e-006, 
    1.215646e-005, 7.379516e-006, -2.618912e-006, -3.915931e-006, 
    3.688983e-007, 2.258614e-006, -1.146556e-006, -1.200693e-006, 
    1.918739e-006, 5.870403e-006, 7.487917e-006, -8.054449e-007, 
    -3.754511e-006, 5.601214e-007, 6.948994e-006, 6.280807e-006, 
    -1.961398e-006, -7.888215e-006, -6.28845e-006, -4.596541e-006, 
    -1.792883e-006, -5.43052e-007, 1.181852e-007, -1.958417e-006, 
    -4.025823e-006, -5.584113e-006, -3.015898e-006, -8.347411e-007, 
    -1.700002e-006, -2.057382e-006, -4.824519e-007, 7.441362e-006, 
    4.820002e-006, -1.177716e-006, 1.243725e-006, 2.424642e-006, 
    9.110541e-006, 5.873226e-007, -2.722101e-006, -6.333321e-007, 
    -1.234963e-006, -1.667095e-006, -2.307723e-006, -4.229349e-006, 
    -3.706069e-006, -3.209489e-006, -2.286488e-006, -2.59072e-006,
  -1.034912e-006, -4.827007e-007, -3.627461e-007, -5.017e-007, 
    -2.683723e-007, -2.116366e-006, -2.682734e-006, -1.578681e-006, 
    -9.907067e-007, -1.351315e-006, -5.851587e-006, -2.796726e-006, 
    -2.170864e-007, -1.288026e-007, -6.982718e-007, -4.315409e-006, 
    -2.89234e-006, -1.35839e-006, -7.238272e-006, -1.114511e-005, 
    -5.132737e-006, 3.546193e-007, -5.56996e-006, -1.436625e-006, 
    5.272195e-007, -1.343369e-006, -1.033301e-006, -3.799083e-006, 
    3.535893e-006, 2.886578e-006, -1.158221e-006, 1.232051e-006, 
    5.304661e-006, 4.490063e-006, 8.905528e-006, 9.436505e-006, 
    8.193128e-006, 4.994718e-006, 3.587303e-006, 5.380036e-006, 
    5.374446e-006, -1.253837e-006, 2.506822e-007, 7.270743e-006, 
    -2.669578e-006, -6.96682e-006, 3.266181e-006, 3.517263e-006, 
    7.171639e-006, -3.866397e-006, -4.798461e-006, 4.198489e-006, 
    5.383627e-006, 3.797271e-006, 1.84833e-006, 7.203311e-006, 1.193281e-005, 
    9.847769e-006, -2.43762e-006, -3.329078e-006, 5.962287e-006, 6.4128e-006, 
    3.386231e-008, -2.72036e-006, -8.764398e-006, -8.44948e-006, 
    -3.211355e-006, -1.239312e-006, -1.5839e-006, -1.822443e-006, 
    -2.136234e-006, -2.917549e-006, -2.629088e-006, -1.335294e-006, 
    -4.524022e-007, -9.430223e-007, -1.334178e-006, -1.684479e-006, 
    1.965436e-006, 1.136298e-005, -1.836344e-006, -5.878906e-006, 
    -1.709191e-006, -2.563523e-006, -2.16206e-006, -4.610944e-006, 
    -6.006565e-006, -3.385698e-006, -3.541039e-006, -2.610339e-006, 
    -2.162309e-006, -1.669084e-006, -1.3538e-006, -8.344914e-007, 
    -4.757458e-007, -5.573293e-007,
  -2.697379e-008, -1.872863e-007, -2.143552e-007, -2.419229e-007, 
    -5.425539e-007, -1.490639e-006, -8.295247e-007, -1.205406e-006, 
    -1.177964e-006, -1.130901e-006, -9.097421e-007, -8.707502e-008, 
    6.430128e-009, 5.859731e-006, 9.361411e-007, -6.426149e-006, 
    -8.92185e-006, -7.771978e-006, -9.737692e-006, -8.740926e-006, 
    -1.841689e-006, -9.85121e-007, -8.678715e-006, -3.366455e-006, 
    -3.065015e-007, -6.417085e-006, -3.170004e-006, 6.185443e-006, 
    3.979949e-006, 3.135803e-006, 4.971496e-006, 2.532674e-006, 
    2.236761e-006, 4.239477e-006, 4.041665e-006, 2.795431e-006, 
    1.145871e-006, 9.105579e-007, 1.018715e-006, 3.232407e-006, 
    6.682894e-007, 2.063516e-007, 8.813633e-006, 8.085217e-006, 
    6.563809e-006, 4.650497e-006, 5.689602e-006, 1.248179e-005, 
    2.838631e-006, -6.437658e-007, 7.368595e-006, 1.155097e-005, 
    9.78629e-006, 2.18334e-005, 1.620051e-005, 1.398297e-005, 7.162202e-006, 
    3.416793e-006, 2.263445e-006, 5.689348e-006, 3.757548e-006, 
    -2.142195e-006, -3.308956e-006, -3.952438e-006, -1.406823e-006, 
    -3.94044e-007, -2.085324e-006, -1.823557e-006, -1.043977e-006, 
    -1.532239e-006, -1.423708e-006, -1.195099e-006, -1.384717e-006, 
    -1.461956e-006, -1.009332e-006, -2.028944e-006, -2.047322e-006, 
    -2.344721e-007, 4.210296e-006, 2.670509e-006, -3.089284e-006, 
    -5.58076e-006, -2.241907e-006, -2.88117e-007, 2.084662e-007, 
    -5.247596e-006, -3.710042e-006, -4.177695e-006, -5.287086e-006, 
    -5.662223e-006, -1.697021e-006, -1.307109e-006, -4.111744e-007, 
    -4.188723e-007, -3.884497e-007, -1.426688e-006,
  -7.469471e-007, -1.118856e-006, 1.847482e-007, -7.958737e-007, 
    -7.263347e-007, -9.642565e-007, -2.424198e-007, -3.351795e-007, 
    -5.136199e-007, -1.12432e-006, -6.716964e-007, 3.743642e-006, 
    7.608005e-007, 2.610036e-006, 4.310015e-006, -1.172002e-006, 
    -8.054321e-007, -3.53928e-007, 1.65388e-006, 9.844553e-006, 4.89637e-006, 
    1.822886e-006, -4.361842e-006, 3.205711e-006, 2.757806e-006, 
    3.434689e-006, 3.6253e-006, 1.784312e-005, 1.209214e-005, 1.085436e-005, 
    9.683368e-006, 8.178722e-006, 4.208061e-006, 4.10338e-006, 8.570373e-007, 
    5.043776e-007, 1.197158e-006, 1.1943e-006, 1.556909e-007, 2.407005e-006, 
    5.247663e-006, 9.501946e-006, 1.344628e-005, 9.653933e-006, 1.15388e-005, 
    1.709433e-005, 1.980583e-005, 6.845938e-006, 3.284222e-007, 
    7.769435e-006, 9.854484e-006, 3.982808e-006, 9.011841e-006, 
    1.485097e-005, 5.589522e-006, 1.132823e-006, 2.964174e-006, 
    4.871894e-006, -1.997105e-007, -1.857989e-007, -1.943266e-006, 
    1.33611e-006, 9.676787e-007, 7.070321e-007, -1.2254e-006, -2.233213e-006, 
    -2.24737e-006, -2.633558e-006, -2.579169e-006, -3.280144e-006, 
    -2.80517e-006, -3.57643e-006, -2.006469e-006, -2.251097e-006, 
    -2.643122e-006, -2.081347e-006, -1.292951e-006, 6.10672e-007, 
    4.183352e-006, -1.736884e-006, -4.54128e-006, -2.980507e-006, 
    -1.569989e-006, -5.47398e-007, 3.769728e-007, -3.622374e-006, 
    -1.613334e-007, -4.325339e-007, -5.652782e-006, -7.130111e-006, 
    -2.645729e-006, 4.289996e-007, -1.808294e-007, -7.196304e-007, 
    -6.497175e-007, 3.253153e-007,
  -3.030182e-007, 6.181335e-008, 2.79133e-008, -1.002878e-006, -2.3746e-008, 
    -1.311081e-006, -3.641048e-008, -1.320259e-007, -9.298587e-007, 
    -1.027711e-006, -1.633692e-006, 3.239609e-006, 1.479906e-006, 
    2.379193e-006, 1.077673e-005, 1.2657e-006, 9.706215e-006, 1.169539e-005, 
    1.512538e-005, 2.670197e-005, 2.229085e-005, 1.468245e-005, 
    2.439291e-005, 2.728983e-005, 2.256752e-005, 7.581555e-006, 
    1.081659e-005, 1.779828e-005, 1.637237e-005, 1.474392e-005, 
    7.445826e-006, 7.307492e-006, 1.467314e-005, 1.107824e-005, 
    4.852785e-006, 2.588429e-006, 4.76673e-006, 3.945427e-006, 
    -5.202032e-007, 2.415323e-006, 5.630875e-006, 1.434122e-005, 
    2.462078e-005, 1.615084e-005, 1.381597e-005, 3.095864e-005, 
    2.277229e-005, 1.207377e-005, 5.698239e-007, -1.308588e-006, 
    6.530034e-006, 1.021299e-005, 1.502097e-005, 8.581934e-006, 
    -3.340378e-006, -5.875314e-006, -4.666454e-006, -3.930956e-006, 
    -3.480698e-006, 6.232112e-007, 2.503988e-006, -7.996005e-007, 
    -2.016156e-006, -2.873966e-006, -3.134982e-006, -3.148145e-006, 
    -3.163792e-006, -2.462195e-006, -2.84441e-006, -3.427543e-006, 
    -3.028812e-006, -2.815726e-006, -2.667336e-006, -2.14033e-006, 
    -9.482374e-007, 1.837411e-006, -1.346227e-006, 2.598987e-006, 
    2.139259e-007, -1.098489e-006, -5.727165e-006, -1.179082e-006, 
    -2.163553e-006, 6.576101e-007, -1.336909e-006, -1.770291e-006, 
    -1.907632e-006, 5.643451e-007, -2.055152e-006, -2.325478e-006, 
    2.071605e-006, 2.291647e-006, 3.900095e-007, -6.925575e-007, 
    2.340202e-006, 5.535512e-007,
  1.524486e-006, 2.866334e-006, 2.166562e-007, 6.954593e-006, 2.177902e-006, 
    1.056217e-006, 1.850697e-006, 1.437811e-006, 1.206595e-006, 
    1.414093e-006, -1.651696e-006, -1.231489e-006, -1.154862e-006, 
    -3.3215e-006, 2.183486e-006, 8.016505e-007, 6.562688e-006, 1.341897e-005, 
    1.454883e-005, 1.817615e-005, 2.759183e-005, 2.53672e-005, 1.601549e-005, 
    3.394048e-005, 2.957369e-005, 3.20447e-006, 4.507194e-006, 5.214133e-006, 
    6.795508e-006, 6.433162e-006, 1.65815e-005, 9.856332e-006, 1.17432e-005, 
    1.977765e-005, 1.886235e-005, 1.243064e-005, 1.14011e-005, 7.454522e-006, 
    8.07429e-006, 3.937145e-005, 4.046817e-005, 2.67904e-005, 1.852521e-005, 
    1.180877e-005, 2.375927e-005, 3.97328e-005, 2.103632e-005, 7.32737e-006, 
    6.763978e-006, -2.746561e-005, -2.881294e-006, 2.908928e-006, 
    1.155595e-005, 1.310927e-005, 3.640598e-007, -1.094345e-005, 
    -5.428898e-006, -7.685056e-006, -4.169382e-006, -5.913073e-006, 
    -2.128661e-006, -1.897812e-006, -1.966113e-006, -2.920653e-006, 
    -2.183295e-006, -1.42048e-006, -1.620403e-006, -1.591842e-006, 
    -2.290335e-006, -2.436244e-006, -2.711914e-006, -2.094013e-006, 
    -2.521676e-006, 1.21292e-007, 5.941813e-006, 2.913519e-006, 
    -7.069641e-006, -2.376391e-006, -2.218067e-007, -1.32636e-006, 
    -3.506768e-006, -2.308343e-006, -4.718106e-006, -1.243157e-006, 
    -2.240045e-006, 1.609043e-006, 1.131593e-006, -3.220339e-008, 
    1.731591e-006, 1.426997e-006, 5.166195e-006, 1.98539e-005, 9.568503e-006, 
    6.874248e-006, 4.48845e-006, 3.241596e-006,
  3.988633e-006, -4.411522e-006, -4.643858e-006, 1.975988e-006, 7.11453e-006, 
    7.40312e-006, 6.289132e-006, 6.866553e-006, 4.615856e-006, 2.623574e-007, 
    -5.933548e-006, -7.548715e-006, -6.572805e-006, -1.081555e-005, 
    -8.120296e-006, -1.412857e-005, -9.915399e-006, -9.090236e-006, 
    4.4271e-006, 1.702801e-005, 2.55557e-005, 1.581294e-005, 1.446428e-005, 
    7.186311e-006, -9.312884e-006, -1.224792e-005, 3.319001e-007, 
    4.209178e-006, 7.085218e-006, 8.539282e-007, 2.264715e-007, 
    2.168694e-006, 4.782611e-006, 3.122994e-006, 4.567919e-006, 
    -2.05588e-006, 3.279842e-006, 3.660679e-005, 4.009491e-005, 
    3.024224e-005, 3.608239e-005, 2.915967e-005, 1.472457e-005, 
    -1.19982e-006, 1.786213e-005, 1.367091e-005, -5.389928e-006, 
    -4.504298e-006, -1.132648e-006, -1.511465e-005, 3.058041e-006, 
    4.043395e-006, 1.620065e-007, 8.362884e-006, 1.568817e-005, 
    9.071184e-006, 8.695184e-006, 6.958573e-006, 5.94405e-006, 
    -3.323221e-007, 1.683802e-006, 7.258968e-007, -1.479275e-007, 
    1.746019e-006, 2.094204e-006, 2.230299e-006, 2.760904e-006, 
    2.374346e-006, 1.173812e-006, 1.843124e-006, 1.245587e-006, 
    2.072726e-006, 1.898008e-006, 4.76114e-006, 6.179853e-006, 1.448239e-006, 
    -5.994252e-007, 2.597495e-006, 6.994316e-006, -9.144678e-007, 
    -3.975163e-006, -3.370053e-006, -3.354406e-006, -9.225838e-006, 
    -3.568362e-006, -1.350567e-006, -1.952096e-006, -8.599382e-007, 
    -1.922774e-006, -5.30012e-006, 3.011621e-006, 3.315406e-005, 
    1.438305e-005, 1.06785e-005, 7.610113e-006, 6.981038e-006,
  -4.493853e-006, -5.758833e-006, -3.380868e-006, -5.743934e-006, 
    2.658577e-006, 7.818344e-006, 3.21725e-006, 1.682449e-005, 1.379919e-005, 
    9.573228e-006, -1.843055e-007, -7.75782e-006, -1.851224e-005, 
    -1.357635e-005, -9.865096e-006, -1.413118e-005, -4.407804e-006, 
    1.346772e-006, 4.244808e-006, 8.527277e-006, 8.351195e-006, 
    1.033578e-005, 9.401843e-006, -7.973722e-007, -7.901122e-006, 
    -4.94386e-006, -6.002352e-006, -4.064605e-007, 6.05578e-007, 
    5.655093e-006, -8.454172e-007, -5.591937e-007, -7.805873e-006, 
    -7.043054e-006, -1.607856e-006, 3.875626e-006, 6.303773e-006, 
    1.675981e-005, 1.948261e-005, 1.940551e-005, 2.184781e-005, 
    1.595539e-005, -2.207758e-006, -2.732007e-005, -1.857136e-005, 
    -1.556182e-005, -1.903303e-005, -1.254617e-005, -1.070177e-006, 
    -2.67553e-006, 2.736073e-006, 8.392301e-006, 4.088968e-006, 
    5.551523e-006, 8.38597e-006, 8.157243e-006, 8.922292e-006, 1.046617e-005, 
    1.181386e-005, 9.021132e-006, 8.423225e-006, 6.677305e-006, 
    5.808195e-006, 6.307384e-006, 5.39655e-006, 4.054828e-006, 4.316711e-006, 
    4.295851e-006, 7.271859e-006, 6.413558e-006, 3.963929e-006, 
    2.348643e-006, 2.471326e-006, 5.664551e-007, -3.581776e-006, 
    5.628011e-006, 4.925922e-006, 6.120252e-006, 6.407208e-007, 
    1.776054e-006, 2.240231e-006, -3.0025e-006, -5.2219e-006, -3.852605e-006, 
    -1.01293e-006, -1.439218e-005, -1.562292e-005, 1.030312e-005, 
    1.523604e-005, -1.502063e-006, -4.373025e-006, 1.247783e-005, 
    -4.273898e-008, 4.369213e-008, 2.803987e-006, -1.770917e-006,
  2.283574e-006, 3.986039e-006, -6.769129e-006, -1.317116e-005, 
    -7.935152e-006, -3.528367e-006, -1.469307e-007, 8.387964e-006, 
    9.771291e-006, 2.33276e-005, 1.701933e-005, 6.081837e-008, 
    -8.133453e-006, -5.777467e-006, -2.42508e-006, 1.184362e-006, 
    1.782268e-006, 7.497485e-006, 8.611594e-006, 1.051423e-005, 
    1.093828e-005, 1.582076e-005, 1.903358e-005, 1.244728e-005, 
    9.038507e-006, -1.418382e-006, 5.564809e-006, -4.276542e-006, 
    -2.720481e-006, -4.928705e-006, 3.108724e-006, 5.625778e-006, 
    1.132968e-006, -6.296512e-006, -2.578912e-006, 4.76835e-006, 
    4.430709e-006, -1.379252e-006, -2.54254e-006, -1.903776e-005, 
    -2.789462e-005, -2.039513e-005, -1.501408e-005, -2.250825e-005, 
    -2.805407e-005, -3.159558e-005, -2.226907e-005, -7.432107e-006, 
    -1.458095e-006, -5.408394e-006, -3.813235e-006, -1.37206e-006, 
    2.188899e-007, -2.678753e-007, 1.54261e-006, 3.32082e-006, 5.170305e-006, 
    5.094805e-006, 5.285166e-006, 5.3593e-006, 5.867554e-006, 5.011358e-006, 
    5.886304e-006, 4.159509e-006, 2.212796e-006, 3.662059e-006, 
    2.713353e-006, 2.662437e-006, 4.665153e-006, 6.282424e-006, 
    8.716408e-006, 9.303763e-006, 1.024949e-005, 4.076304e-006, 
    5.560956e-006, -9.258474e-006, -5.625952e-006, 2.701418e-006, 
    1.942346e-006, 1.181259e-006, 3.46126e-006, -1.065338e-006, 
    -6.800425e-006, -9.400181e-006, -7.352515e-006, -4.901034e-006, 
    -9.219184e-007, 1.534282e-005, 2.177206e-005, 4.439145e-006, 
    3.844711e-006, -1.458597e-006, 8.050331e-006, 2.064648e-006, 
    6.321541e-006, 5.727976e-006,
  3.257861e-006, 4.120375e-006, 1.405278e-006, -1.133633e-005, 
    -1.033163e-005, 5.583679e-006, 3.815047e-006, -1.42495e-005, 
    -1.173556e-005, 1.064512e-005, 4.245524e-005, 6.608265e-006, 
    -3.031048e-006, 4.857488e-006, 1.781646e-006, 5.509046e-006, 
    1.061766e-005, 1.183894e-005, 1.28213e-005, 1.071552e-005, 1.446762e-005, 
    1.683057e-005, 1.724085e-005, 1.101055e-005, 7.762734e-006, 
    -2.725585e-006, 7.307997e-006, 1.18177e-005, -1.19726e-005, 
    -1.373926e-005, -4.902642e-006, -9.559444e-007, -9.750656e-007, 
    -2.660869e-006, -4.183523e-006, 1.210203e-006, 7.242561e-006, 
    3.645539e-006, -5.175709e-006, -6.989649e-006, -3.379231e-006, 
    -5.132752e-007, 1.8766e-005, 1.3659e-005, 1.656612e-006, 5.110327e-006, 
    2.832239e-007, 8.067509e-007, 5.848437e-006, 5.580463e-006, 
    7.232884e-006, 6.368362e-006, 7.073315e-006, 7.004637e-006, 
    6.639319e-006, 5.637572e-006, 4.908521e-006, 3.675203e-006, 2.46759e-006, 
    3.653859e-006, 3.31051e-006, 2.005676e-006, 1.959477e-006, 3.411096e-006, 
    6.040156e-006, 4.690484e-006, 7.303155e-006, 7.490038e-006, 
    1.026575e-005, 1.724806e-005, 1.18249e-005, 1.514501e-005, 1.668655e-005, 
    1.42559e-005, 3.100024e-006, -2.329938e-005, -9.869676e-006, 
    -1.477856e-006, -1.071633e-005, -4.197314e-006, -2.136107e-007, 
    3.429477e-007, -1.566263e-006, -4.206374e-006, -3.732271e-006, 
    -1.447177e-006, -1.729307e-006, -1.578557e-006, -5.841534e-007, 
    -1.906133e-006, 4.491194e-007, -3.264384e-006, 1.845721e-006, 
    1.410233e-006, -7.828494e-007, -4.070898e-007,
  -1.045369e-005, -1.35381e-005, -1.025265e-005, -1.518718e-006, 
    -2.979024e-006, -1.216227e-006, -3.865396e-006, -4.162306e-006, 
    -1.316471e-005, -1.253277e-005, -3.474383e-005, -2.298531e-006, 
    -3.017389e-006, 4.399037e-006, 9.539937e-006, 9.875836e-006, 
    1.614636e-005, 1.401562e-005, 1.481781e-005, 1.096201e-005, 
    1.200671e-005, 1.040719e-005, 2.264736e-005, 2.101595e-005, 
    8.628725e-006, -8.835414e-007, 6.89349e-006, 7.69406e-006, -2.4498e-006, 
    -8.381176e-006, -1.192604e-005, -1.089203e-005, 1.357104e-006, 
    -7.280738e-006, 1.137875e-005, 1.445957e-005, 1.282168e-005, 
    1.426349e-005, 2.048423e-005, 2.898658e-005, 1.853293e-005, 
    1.658635e-005, 2.285325e-005, 1.677607e-005, 1.904153e-005, 
    1.042195e-005, 9.742835e-006, 7.980398e-006, 1.074419e-005, 
    1.165863e-005, 1.174059e-005, 1.472566e-005, 1.29857e-005, 1.217918e-005, 
    1.111188e-005, 8.734281e-006, 5.400889e-006, 1.686778e-006, 
    -2.187026e-006, -5.440816e-006, -7.200149e-006, -1.010984e-005, 
    -7.724044e-006, -3.702226e-006, 2.365232e-007, 3.717552e-006, 
    9.184914e-006, 1.577148e-005, 1.657205e-005, 1.658012e-005, 
    2.009891e-005, 1.642887e-005, 4.863759e-007, 4.452573e-006, 
    -8.591043e-006, -1.020844e-005, -1.84314e-005, -1.798127e-005, 
    -5.693516e-006, 2.593774e-007, 6.934988e-007, 7.589397e-007, 
    -7.869321e-007, -3.43498e-007, -7.643312e-007, -1.713288e-006, 
    -9.974119e-007, -1.348086e-006, -7.753847e-007, -7.829594e-007, 
    1.010533e-007, -1.208387e-006, -9.519757e-006, -5.898652e-006, 
    -7.78502e-006, -6.726536e-006,
  3.738915e-006, 9.28485e-008, -1.008972e-006, -2.559424e-006, 
    -5.156824e-006, -6.143035e-006, -6.146012e-006, -6.611798e-006, 
    -6.785645e-006, -1.156706e-005, -8.995237e-006, -1.046461e-006, 
    -3.853715e-006, -4.818303e-007, 7.945884e-006, 7.803588e-006, 
    7.294961e-006, 1.01345e-005, 7.332834e-006, 5.698799e-006, 4.927787e-006, 
    1.064871e-005, 3.544759e-005, 1.720846e-005, 2.003806e-005, 
    -8.444877e-006, -1.098441e-005, 5.331101e-006, 1.609595e-005, 
    -6.680217e-006, -1.024159e-005, -1.789979e-005, -5.700844e-006, 
    -3.946625e-007, -4.543646e-006, -1.342989e-006, 1.855639e-005, 
    2.787398e-005, 2.729467e-005, 2.235519e-005, 1.499835e-005, 
    7.575087e-006, 1.022104e-005, 1.915541e-005, 1.444714e-005, 
    6.450931e-006, 9.440231e-006, 1.188303e-005, 8.89982e-006, 4.755308e-006, 
    3.215522e-006, 3.471072e-006, 1.919736e-006, 2.889055e-006, 
    3.386759e-006, 2.487598e-006, 1.537152e-006, 1.165754e-007, 
    -1.124054e-007, -1.005235e-006, -9.770474e-007, -1.97741e-006, 
    -3.476467e-006, -3.730159e-006, -4.939389e-006, -6.088518e-006, 
    -3.654786e-007, 7.910858e-006, 1.603003e-005, 1.35917e-005, 
    1.420239e-005, 7.055176e-006, -6.281371e-006, -2.381606e-006, 
    -5.89692e-006, -1.374585e-005, -1.493112e-005, -1.168838e-005, 
    -5.803533e-006, -4.247104e-007, -5.553375e-008, 2.251036e-007, 
    -5.877528e-007, -4.901513e-007, -8.24185e-007, -7.355229e-007, 
    -8.782017e-007, -1.417501e-006, -2.610464e-007, -2.403085e-007, 
    3.511434e-007, 2.814803e-007, -3.517696e-006, -4.520171e-006, 
    1.261105e-006, 7.736653e-006,
  -6.111804e-009, 1.256014e-006, -1.549004e-006, -2.211979e-006, 
    -7.254584e-008, -6.396594e-007, -1.382482e-006, -3.177948e-006, 
    -3.386068e-006, -3.452998e-006, -3.703587e-006, -1.75824e-006, 
    -7.050886e-006, -1.801701e-006, -2.722213e-007, 4.341669e-006, 
    5.375814e-006, 4.810811e-006, 4.225074e-006, 2.450594e-006, 2.35684e-006, 
    5.308015e-006, 2.019564e-005, 1.77557e-005, 2.048869e-005, 1.231887e-005, 
    3.55191e-006, 7.906778e-006, 9.404586e-006, 5.956339e-006, 
    -1.833292e-005, -2.438665e-005, -2.013386e-005, -1.236476e-005, 
    -1.660191e-005, -1.357064e-005, 3.178131e-006, 7.865416e-006, 
    1.16934e-005, 1.122227e-005, 9.617106e-007, 2.234527e-006, 5.952488e-006, 
    8.598687e-006, 9.516472e-006, 4.899721e-006, 4.028128e-006, 
    4.406002e-006, 2.318595e-006, 2.514422e-006, 2.765155e-007, 
    -1.11774e-006, -4.670546e-007, -2.047321e-006, -7.398676e-007, 
    9.391197e-007, -2.575653e-007, -1.858452e-006, -2.470268e-006, 
    -1.843052e-006, -1.81387e-006, -3.565129e-006, -3.001494e-006, 
    -1.544905e-006, -3.347077e-006, -1.915074e-006, -5.42616e-006, 
    -9.175539e-006, -3.762332e-006, 6.83227e-006, 2.661312e-006, 
    4.002166e-006, 3.570789e-006, 1.245063e-005, 6.403534e-007, 
    -9.422771e-006, -1.103707e-005, -9.333497e-006, -8.563602e-006, 
    -3.819444e-006, -1.190132e-006, 7.634208e-008, -2.122433e-007, 
    -6.458686e-007, -8.305169e-007, -7.54646e-007, -1.220556e-006, 
    -1.187153e-006, -9.17194e-007, -2.481318e-007, -9.353221e-008, 
    -1.593458e-007, -3.285237e-006, -4.975027e-006, 1.320836e-006, 
    2.425755e-006,
  5.790071e-007, -3.367923e-007, -1.076637e-006, -1.067944e-006, 
    -1.69491e-006, -1.343616e-006, -7.385031e-007, -1.843301e-006, 
    -1.481451e-006, -2.826405e-006, -7.365672e-006, -2.355404e-006, 
    -3.005964e-006, -2.119593e-006, -9.353221e-008, 2.088619e-006, 
    1.135441e-006, 7.126209e-007, 1.104149e-006, 1.111476e-006, 
    2.296987e-007, 1.774701e-006, 1.000349e-005, 1.001964e-005, 7.91435e-006, 
    5.09579e-007, 5.023867e-007, 1.055e-005, 9.969721e-006, -2.421715e-006, 
    -3.034653e-006, -4.839185e-006, -1.453399e-005, -1.15221e-005, 
    -1.914418e-005, -6.049406e-006, 1.661323e-006, 6.782138e-007, 
    7.978542e-006, 4.976704e-006, -9.437645e-007, 2.83093e-007, 
    5.295844e-006, 6.337808e-006, 5.626899e-006, 3.593515e-006, 
    2.402288e-006, 3.397189e-006, 3.904327e-006, 4.359557e-006, 
    1.469974e-006, 5.063657e-007, 1.000461e-006, 3.32021e-007, 6.640685e-007, 
    1.065034e-006, -2.101333e-007, -9.55938e-007, -1.051179e-006, 
    -2.866885e-006, -9.907062e-007, -2.209247e-006, -1.332935e-006, 
    -1.358393e-006, -5.175943e-007, -9.928181e-007, 2.403776e-007, 
    -1.347589e-006, -5.744549e-006, -1.775268e-006, -5.361351e-006, 
    -3.60002e-006, -2.216839e-007, 2.608169e-006, 2.545239e-007, 
    -7.173698e-006, -1.085913e-005, -1.190755e-005, -1.011233e-005, 
    -6.345811e-006, -4.115855e-006, -2.574699e-006, 2.494444e-007, 
    1.248955e-007, 2.79133e-008, -7.270792e-007, -1.344732e-006, 
    -9.085006e-007, -8.363554e-007, -6.906839e-008, 2.443539e-008, 
    -2.706079e-007, -1.44246e-006, -1.624006e-006, 7.332342e-007, 
    8.951597e-007,
  2.395091e-007, -2.747061e-007, 7.398103e-008, 1.329649e-007, 7.497601e-008, 
    -3.18787e-007, -3.857183e-007, -1.311329e-006, -1.894834e-006, 
    -1.784938e-006, -2.530865e-006, -2.577059e-006, -2.592705e-006, 
    -4.238911e-006, -3.328326e-006, -1.271469e-006, -1.402971e-006, 
    -1.560303e-006, -1.929976e-007, -3.492114e-007, 8.714414e-008, 
    2.039817e-006, 6.865805e-006, 7.289121e-006, 1.096574e-005, 1.27961e-005, 
    5.565431e-006, 4.646898e-006, 8.590108e-006, 7.620401e-007, 
    -1.234621e-007, 1.59911e-007, -5.214564e-006, -1.045816e-005, 
    -1.562477e-005, -2.066782e-005, -9.727388e-006, -1.596072e-006, 
    -4.04942e-006, -5.186999e-006, 1.245957e-006, 6.95607e-007, 
    1.295875e-006, 2.043043e-006, 5.155523e-006, 5.135781e-006, 
    2.238996e-006, 1.103404e-006, 3.333871e-007, 1.610306e-007, 
    2.540392e-007, -1.566263e-006, -1.016162e-006, -1.130405e-006, 
    1.1907e-006, 1.160152e-006, -3.371651e-007, -6.636246e-007, 
    -5.257889e-007, -2.878669e-007, 7.877497e-007, -1.373789e-006, 
    -1.537826e-006, -1.159833e-006, -8.218249e-007, 1.848712e-007, 
    8.361758e-007, 1.08279e-006, -2.022984e-006, -7.192648e-008, 
    6.559949e-006, 7.111303e-007, 2.55192e-006, -9.332125e-007, 
    -2.765191e-006, -9.670392e-006, -1.364527e-005, -1.15976e-005, 
    -1.07229e-005, -1.050907e-005, -8.814065e-006, -4.677255e-006, 
    -1.639401e-006, -1.645603e-007, 1.606577e-007, -4.021094e-007, 
    -1.52515e-007, -7.157796e-007, -9.576752e-007, -1.373542e-006, 
    -3.67962e-007, -3.882028e-007, -6.972776e-007, -4.227239e-007, 
    -1.194604e-006, -4.748777e-007,
  7.860092e-007, 4.758169e-007, 9.936316e-007, 3.403393e-007, 1.980338e-007, 
    -1.455001e-006, -1.977163e-006, -2.160323e-006, -1.802571e-006, 
    -1.895331e-006, -1.969961e-006, -2.155107e-006, -2.731286e-006, 
    -3.324104e-006, -3.349188e-006, -4.36582e-006, -2.866886e-006, 
    -1.571479e-006, -1.154991e-006, -9.189325e-007, 1.096698e-006, 
    4.564075e-006, 2.911039e-006, 2.438051e-006, 9.365229e-006, 
    2.296342e-005, 2.367073e-005, 1.105079e-005, 5.350219e-006, 
    7.260191e-006, 6.059396e-006, 8.630093e-006, 7.525054e-006, 
    1.370376e-006, -8.896277e-007, -7.464274e-006, -7.653023e-006, 
    -1.925138e-006, -1.388074e-006, -2.775119e-006, 2.977598e-006, 
    3.523844e-006, 1.951279e-006, 2.824985e-006, 1.4773e-006, 2.513052e-006, 
    1.83654e-006, 2.019081e-006, 5.293359e-007, -1.023986e-006, 
    -1.128666e-006, -1.454379e-006, -2.21558e-006, -2.723463e-006, 
    -9.736941e-007, -1.779717e-007, 2.823508e-007, 2.271531e-006, 
    -1.640628e-007, -3.46603e-007, -2.138586e-007, -1.088309e-006, 
    -7.97861e-007, -1.421723e-006, 1.736953e-007, -2.465169e-007, 
    -4.788508e-007, 1.603089e-006, 7.855115e-007, 6.494156e-007, 
    6.161603e-006, 6.224809e-006, 5.466214e-006, 3.451206e-006, 
    -2.239549e-006, -5.943983e-006, -1.350521e-005, -1.344249e-005, 
    -9.906438e-006, -6.797312e-006, -7.31265e-006, -6.193321e-006, 
    -3.396994e-006, -8.287798e-007, -1.968465e-007, -3.755349e-007, 
    -4.044687e-007, -1.173617e-006, -8.757193e-007, -1.263522e-006, 
    -1.205532e-006, -4.114231e-007, -5.070387e-007, -2.403089e-007, 
    -2.750782e-007, -1.371555e-006,
  -1.352804e-006, -1.467419e-006, -1.152509e-006, 2.26969e-008, 
    -9.800351e-008, -5.870088e-007, -1.815736e-006, -2.784062e-006, 
    -2.238555e-006, -2.553093e-006, -3.888486e-006, -3.492363e-006, 
    -1.605627e-006, -2.879676e-006, -5.5147e-006, -5.46031e-006, 
    -5.129006e-006, -3.857442e-006, -5.635397e-006, -1.142946e-006, 
    4.262699e-007, -2.809156e-008, 7.808012e-008, 4.758163e-007, 
    -2.313682e-007, 4.737426e-006, 1.4334e-005, 1.030524e-005, 1.379957e-005, 
    1.104372e-005, 1.396721e-005, 1.776068e-005, 1.053932e-005, 
    6.676673e-006, 1.659952e-006, 3.406862e-006, -4.411646e-006, 
    -1.068764e-005, -5.929945e-006, -1.842938e-006, 2.236047e-007, 
    2.389741e-006, 4.699552e-006, 5.757038e-006, 2.490331e-006, 
    1.316117e-006, -1.590357e-006, -2.891969e-006, 2.313118e-007, 
    -1.997901e-006, -3.051164e-006, -3.479075e-006, -5.549343e-006, 
    -5.830479e-006, -4.597904e-006, -3.894196e-006, -4.038986e-006, 
    -1.362738e-006, -4.167623e-007, -1.87869e-006, -1.559309e-006, 
    -1.338897e-006, -9.132204e-007, -1.332936e-006, -8.619352e-007, 
    8.813822e-008, -8.436814e-007, -3.180059e-006, -2.672179e-006, 
    3.943063e-006, 7.496994e-006, 7.760742e-006, 5.602433e-006, 
    4.797526e-006, 2.975235e-006, -2.675042e-007, -6.873441e-006, 
    -1.190109e-005, -1.010848e-005, -6.717097e-006, -7.625322e-006, 
    -5.789128e-006, -4.691903e-006, -3.070778e-006, -2.371919e-006, 
    -9.967898e-007, -3.62621e-007, -1.663619e-006, -1.460466e-006, 
    -1.172128e-006, -1.067448e-006, -8.926067e-007, -3.140694e-007, 
    -2.915933e-007, -1.134998e-006, -2.026709e-006,
  -3.118964e-006, -2.974671e-006, -3.937906e-006, -3.872962e-006, 
    -1.716392e-006, -2.039498e-006, -2.450026e-006, -2.160819e-006, 
    -1.652319e-006, -2.09662e-006, -3.217933e-006, -3.228488e-006, 
    -5.46838e-006, -1.134142e-005, -9.642446e-006, -4.493969e-006, 
    -4.654281e-006, -9.888066e-006, -1.103968e-005, -5.699349e-006, 
    -1.661133e-006, 6.71891e-007, 2.641447e-006, 5.500488e-006, 
    6.806942e-006, 3.164235e-006, 3.849562e-006, 1.264868e-005, 
    1.741943e-005, 1.868529e-005, 1.123173e-005, 9.797601e-006, 
    1.283595e-005, 1.242752e-005, 7.67281e-006, 2.849934e-006, 
    -1.213979e-006, -8.561248e-006, -6.132483e-006, -6.720205e-006, 
    -7.858158e-006, -8.196665e-006, -6.155453e-006, -7.102666e-006, 
    -7.100803e-006, -3.615052e-006, -1.323628e-006, -3.704408e-007, 
    -5.538539e-006, -5.195192e-006, -4.031039e-006, -6.871072e-006, 
    -1.03988e-005, -9.899367e-006, -9.359571e-006, -6.676741e-006, 
    -6.529219e-006, -5.977628e-006, -3.922015e-006, -4.647077e-006, 
    -3.997884e-006, -2.730168e-006, -1.824302e-006, -6.772843e-007, 
    -1.649213e-006, -1.851248e-006, -1.994672e-006, -3.627094e-006, 
    -5.99638e-006, -2.731163e-006, 4.380541e-006, 8.231244e-006, 
    7.425973e-006, 5.387112e-006, 7.754159e-006, 5.672602e-006, 
    8.813731e-008, -6.233309e-006, -1.195597e-005, -1.002367e-005, 
    -9.684918e-006, -5.351905e-006, -4.208488e-006, -6.465765e-006, 
    -6.506121e-006, -4.860166e-006, -2.373037e-006, -1.501442e-006, 
    -2.072405e-006, -1.590602e-006, -1.981385e-006, -3.129146e-006, 
    -3.119212e-006, -3.195953e-006, -5.493589e-006, -3.173477e-006,
  -6.916523e-006, -5.819057e-006, -2.731782e-006, -3.929341e-006, 
    -3.242396e-006, -3.617532e-006, -5.55816e-006, -3.064077e-006, 
    -3.018131e-006, -4.226993e-006, -2.166285e-006, -4.266352e-006, 
    -6.520901e-006, -7.217528e-006, -4.794725e-006, -3.688684e-006, 
    -4.747412e-006, -4.048548e-006, -3.498943e-006, -5.573809e-006, 
    -5.178059e-006, 1.398075e-006, 8.356787e-007, 2.927054e-006, 
    7.644891e-006, 5.812291e-006, 6.079767e-006, 7.057659e-006, 
    7.735041e-006, 1.296397e-005, 1.642923e-005, 1.620733e-005, 
    1.836912e-005, 1.833857e-005, 1.883429e-005, 1.915007e-005, 
    1.650325e-005, 1.014145e-005, 1.028147e-006, -4.920221e-007, 
    3.269903e-006, 4.700778e-006, 4.066875e-006, 6.518894e-007, 
    -3.142435e-006, -3.075889e-006, -9.232826e-007, 4.134708e-007, 
    4.453868e-007, -2.431403e-006, -4.672787e-006, -7.876664e-006, 
    -7.327677e-006, -7.42478e-006, -8.22895e-006, -9.007897e-006, 
    -8.109986e-006, -7.335128e-006, -5.687429e-006, -4.479562e-006, 
    -6.602355e-006, -2.132383e-006, -5.497559e-007, -3.004224e-006, 
    -4.03576e-006, -5.131365e-006, -4.410895e-006, -3.441945e-006, 
    -6.715361e-006, -1.008067e-005, -2.520064e-006, 2.272762e-006, 
    6.356306e-006, 7.850391e-006, 8.446437e-006, 8.990082e-006, 
    5.457267e-006, 4.142239e-007, -2.609475e-006, -5.896298e-006, 
    -6.739952e-006, -6.030408e-006, -4.199675e-006, -4.301124e-006, 
    -6.461296e-006, -8.679086e-006, -7.027415e-006, -4.257165e-006, 
    -3.927724e-006, -3.043341e-006, -3.955663e-006, -3.097853e-006, 
    -1.983868e-006, -4.120448e-006, -4.755982e-006, -4.237049e-006,
  -1.010587e-005, -2.427798e-006, -4.388793e-006, -6.148992e-006, 
    -3.388301e-006, -4.369793e-006, -5.324961e-006, -2.263763e-006, 
    -1.205408e-006, 2.145738e-006, 4.640569e-006, 7.653871e-007, 
    -2.030691e-006, -7.589824e-008, -1.731914e-006, -2.309085e-006, 
    -3.06296e-006, -2.63331e-006, -1.443205e-006, 3.181131e-007, 
    -2.264009e-006, 1.060063e-006, 2.486855e-006, 1.411859e-006, 
    1.501141e-006, 1.330523e-006, 2.793568e-006, 5.10027e-006, 2.127859e-006, 
    2.538012e-006, 3.609282e-006, 6.152664e-006, 9.269615e-006, 
    9.899561e-006, 9.666721e-006, 1.062363e-005, 1.305041e-005, 
    9.816984e-006, 7.764094e-006, 3.366764e-006, 1.880122e-006, 
    7.803337e-006, 1.016293e-005, 1.125767e-005, 8.295945e-006, 
    7.942781e-006, 4.169182e-006, 4.822356e-006, 9.242911e-006, 9.95916e-006, 
    8.315808e-006, 4.839494e-006, 2.796922e-006, 1.565604e-007, 
    -2.133875e-006, -7.652401e-006, -4.734498e-006, -4.680731e-006, 
    -3.986588e-006, -5.625219e-006, -4.575797e-006, -2.249608e-006, 
    -1.04398e-006, -3.061972e-006, -6.37015e-006, -4.956151e-006, 
    -1.674793e-006, -4.398607e-007, 7.427916e-007, -6.836679e-006, 
    -3.533842e-006, -4.432139e-006, 1.646662e-006, 4.737794e-006, 
    5.663158e-006, 9.118612e-006, 7.220569e-006, 6.503451e-006, 5.89413e-006, 
    2.01572e-006, -1.191132e-006, -3.539804e-006, 1.185232e-006, 
    2.076569e-006, -1.063603e-006, -2.591834e-006, -2.861547e-006, 
    -7.425648e-006, -4.86588e-006, -4.205758e-006, -2.593451e-006, 
    -2.972933e-006, -3.480318e-006, -3.639387e-006, -5.369284e-006, 
    -1.273096e-005,
  -2.146046e-006, -1.870128e-006, -3.339883e-006, 7.160888e-007, 
    3.173916e-006, 2.299475e-007, 8.605093e-007, 1.076081e-006, 
    -1.961052e-007, 2.89001e-008, 3.187457e-006, 2.572537e-006, 
    4.815302e-007, -9.849919e-008, 1.838403e-006, 2.24148e-006, 1.32332e-006, 
    1.395094e-006, 1.004063e-006, 6.530163e-007, 8.792667e-007, 
    2.394964e-006, 2.663552e-006, 3.428107e-006, 2.618604e-006, 
    2.799653e-006, 2.978964e-006, 2.717323e-006, 2.674486e-006, 
    1.794318e-006, 1.242977e-006, 3.780024e-006, 5.736298e-006, 
    4.286045e-006, 5.750082e-006, 7.65495e-006, 5.870908e-006, 5.252881e-006, 
    4.977333e-006, 5.330612e-006, 3.554524e-006, 6.775655e-006, 
    8.356667e-006, 6.890019e-006, 7.914598e-006, 9.849766e-006, 
    1.118453e-005, 1.061208e-005, 1.044916e-005, 1.18788e-005, 1.137341e-005, 
    9.863801e-006, 6.501105e-006, 4.280831e-006, 1.881494e-006, 
    -2.905756e-006, -2.585259e-006, 1.022312e-006, 1.576886e-006, 
    -2.851393e-007, -9.469659e-009, 2.173427e-006, -6.845039e-008, 
    -1.168402e-006, 2.675715e-007, -8.334791e-008, 3.179879e-006, 
    5.947151e-006, 3.242594e-006, 2.956349e-007, 2.280842e-006, 
    5.109956e-006, 6.516504e-006, 4.953868e-006, 5.837013e-006, 
    1.081263e-005, 1.564196e-005, 7.382499e-006, 6.037171e-006, 
    6.232007e-006, 3.54409e-006, 4.554884e-006, 3.874895e-006, 4.480753e-006, 
    5.289636e-006, 6.839606e-006, 6.427837e-006, 4.134781e-007, 
    -4.795722e-006, -6.524504e-006, -4.05526e-006, -1.686096e-006, 
    -2.663861e-006, -1.261416e-006, 2.017532e-007, -1.803688e-006,
  -8.297757e-007, -2.376393e-006, 1.526965e-006, 3.944559e-006, 
    3.500374e-006, 1.98865e-006, 2.229806e-006, 3.567311e-006, 1.769735e-006, 
    5.616221e-007, 2.471454e-006, 3.268169e-006, 1.71547e-006, 2.419425e-006, 
    1.882734e-006, 1.847468e-006, 2.395335e-006, 1.714601e-006, 
    2.298229e-006, 2.133695e-006, 2.408374e-006, 1.749741e-006, 
    2.166354e-006, 2.789218e-006, 2.2349e-006, 1.397455e-006, 3.410722e-006, 
    2.45593e-006, 1.694234e-006, 3.140638e-006, 2.596373e-006, 3.909539e-006, 
    5.818501e-006, 4.019932e-006, 4.881344e-006, 4.584683e-006, 3.98454e-006, 
    2.773448e-006, 1.765386e-006, 3.252026e-006, 3.075942e-006, 
    3.473064e-006, 6.565548e-006, 7.691577e-006, 7.621915e-006, 
    7.553741e-006, 1.042209e-005, 1.079053e-005, 9.055035e-006, 
    6.817134e-006, 5.773552e-006, 6.764109e-006, 7.892246e-006, 
    5.537115e-006, 2.808965e-006, 9.863015e-007, 1.238255e-006, 2.15269e-006, 
    1.880122e-006, 1.99275e-006, 1.110602e-006, 2.688887e-006, 2.622703e-006, 
    2.197394e-006, 3.689132e-006, 3.935869e-006, 4.217867e-006, 
    5.337568e-006, 6.505566e-006, 2.685161e-006, 4.202351e-006, 
    8.489043e-006, 9.293577e-006, 7.429813e-006, 7.184321e-006, 
    7.771179e-006, 9.955436e-006, 8.672323e-006, 7.11565e-006, 8.686471e-006, 
    9.224037e-006, 9.543917e-006, 6.78596e-006, 3.387629e-006, 3.390731e-006, 
    5.886177e-006, 5.054198e-006, 7.06784e-006, 9.259511e-007, 
    -2.239178e-006, -3.196328e-006, -2.950832e-006, -3.728053e-006, 
    -2.987341e-006, -4.167632e-007, -2.096367e-007,
  1.022318e-006, 1.575397e-006, 2.572534e-006, 3.059804e-006, 1.565568e-007, 
    7.213112e-007, 2.719931e-006, 4.29399e-006, 3.805728e-006, 3.011126e-006, 
    3.517764e-006, 2.901724e-006, 4.212161e-006, 2.999453e-006, 
    3.203847e-006, 3.519996e-006, 4.125358e-006, 3.911777e-006, 
    4.921455e-006, 2.887321e-006, 2.151825e-006, 2.739304e-006, 3.39284e-006, 
    3.520619e-006, 3.43258e-006, 2.616365e-006, 2.0387e-006, 2.438921e-006, 
    3.813302e-006, 2.517027e-006, 8.205279e-008, -3.473506e-007, 
    2.670877e-006, 1.95724e-006, 3.248919e-006, 4.803112e-006, 4.550908e-006, 
    1.924954e-006, 1.266696e-006, 3.016592e-006, 3.99398e-006, 4.946289e-006, 
    5.403877e-006, 1.002734e-005, 9.518959e-006, 8.608748e-006, 
    7.709961e-006, 6.862827e-006, 6.17427e-006, 6.346501e-006, 7.844066e-006, 
    7.926892e-006, 7.320785e-006, 5.489184e-006, 5.605789e-006, 
    3.242463e-006, 3.058931e-006, 5.209295e-006, 2.619345e-006, 
    8.374136e-007, 3.440777e-006, 4.71557e-006, 5.738777e-006, 3.967658e-006, 
    4.68179e-006, 8.211749e-006, 9.272713e-006, 6.408961e-006, 7.072189e-006, 
    4.587666e-006, 4.387246e-006, 6.395923e-006, 7.133529e-006, 
    6.939194e-006, 2.852799e-006, 3.94257e-006, 7.384861e-006, 8.417266e-006, 
    8.438996e-006, 5.895863e-006, 5.13516e-006, 5.417163e-006, 3.782134e-006, 
    2.091845e-006, 4.715814e-006, 7.19003e-006, 5.127957e-006, 2.741162e-006, 
    6.299178e-007, -2.056888e-006, 1.599981e-006, 1.855164e-006, 
    -4.065823e-007, -2.035558e-007, -1.505048e-006, 1.468688e-007,
  2.863604e-006, 2.506968e-006, 3.610151e-006, 3.014105e-006, 7.24167e-007, 
    1.086517e-006, 3.016838e-006, 5.273368e-006, 7.828918e-006, 
    5.175643e-006, 2.941835e-006, 3.418174e-006, 3.229301e-006, 
    3.290151e-006, 4.025894e-006, 4.726995e-006, 3.415817e-006, 
    1.333502e-006, 1.973508e-006, 3.444626e-006, 3.46437e-006, 1.947927e-006, 
    1.606939e-006, 2.129598e-006, 3.140641e-006, 2.058073e-006, 
    4.335961e-007, 1.017474e-006, 1.44042e-006, 1.915391e-006, 3.299954e-006, 
    4.92791e-006, 2.591037e-006, 1.520884e-006, 9.795967e-007, 1.875527e-006, 
    2.217514e-006, 1.351136e-006, 9.751302e-007, 1.792708e-006, 2.37795e-006, 
    2.900857e-006, 5.303295e-006, 9.343991e-006, 8.919185e-006, 
    6.724496e-006, 5.760019e-006, 3.640454e-006, 3.475548e-006, 
    4.487333e-006, 4.720907e-006, 4.723515e-006, 5.110574e-006, 
    5.145097e-006, 5.85178e-006, 7.491903e-006, 8.062118e-006, 6.688355e-006, 
    2.527831e-006, 4.997944e-006, 9.03107e-006, 8.985251e-006, 5.752318e-006, 
    1.261227e-006, 1.662074e-006, 4.131941e-006, 3.750968e-006, 
    3.843231e-006, 4.11257e-006, 1.846598e-006, 1.989772e-006, 3.331746e-006, 
    3.939962e-006, 3.227438e-006, 2.539503e-006, 2.319834e-006, 
    3.023044e-006, 3.176526e-006, 3.110837e-006, 4.142992e-006, 
    3.912148e-006, 3.361425e-006, 8.042643e-007, -9.396699e-007, 
    8.235093e-007, 1.815679e-006, 1.639599e-006, 7.04551e-007, 1.73956e-006, 
    -1.112876e-007, -3.158093e-007, -1.455381e-006, -5.954571e-007, 
    4.488684e-007, 2.223349e-006, 1.093345e-006,
  1.694111e-006, 2.33126e-006, 3.200244e-006, 1.400058e-006, -5.677794e-008, 
    1.821512e-006, 1.824247e-006, 2.479402e-006, 4.102014e-006, 4.66975e-006, 
    2.042798e-006, 8.084844e-007, 2.323807e-006, 2.751598e-006, 
    3.034099e-006, 2.68417e-006, 1.909061e-006, 7.286408e-007, 1.502508e-006, 
    1.842873e-006, 2.04553e-006, 1.675485e-006, -2.594306e-007, 
    -2.153483e-007, 7.278941e-007, 2.441777e-006, 3.189071e-006, 
    1.833437e-006, 1.031258e-006, 1.193307e-006, 3.341062e-006, 
    3.835161e-006, 1.824372e-006, 1.649656e-006, 1.853676e-006, 
    1.575026e-006, 9.428441e-007, 1.061928e-006, 1.719318e-006, 
    2.326168e-006, 2.260604e-006, 9.047217e-007, 1.685542e-006, 
    3.709119e-006, 4.222714e-006, 4.877e-006, 3.797285e-006, 2.489957e-006, 
    1.856532e-006, 1.84424e-006, 3.316477e-006, 4.71818e-006, 4.511548e-006, 
    5.263559e-006, 6.655329e-006, 8.393052e-006, 1.238557e-005, 
    1.044954e-005, 6.621425e-006, 4.622807e-006, 4.750955e-006, 
    2.789468e-006, 9.692958e-007, 2.24607e-007, 7.404369e-007, 1.011388e-006, 
    1.475808e-006, 1.761539e-006, 2.899866e-006, 1.808974e-006, 
    2.127859e-006, 3.397686e-006, 3.700552e-006, 1.644689e-006, 
    1.790473e-006, 2.896139e-006, 1.765141e-006, 1.584959e-006, 
    1.673124e-006, 1.987787e-006, 2.611649e-006, 1.494683e-006, 
    5.165439e-007, 1.305192e-006, 3.106617e-006, 7.069206e-006, 
    4.189562e-006, 1.63637e-006, 2.209437e-006, 2.395707e-006, 2.005199e-007, 
    1.170582e-006, 2.659084e-006, 4.414193e-006, 5.052332e-006, 4.095803e-006,
  1.699822e-006, 1.262474e-006, 1.463392e-006, 1.769983e-006, 9.339037e-007, 
    1.224227e-006, 1.836417e-006, 3.269289e-006, 4.799012e-006, 
    3.897492e-006, 2.51591e-006, 4.473804e-007, -5.270304e-007, 
    5.997463e-007, 1.999709e-006, 2.457672e-006, 2.103894e-006, 
    1.562111e-006, 1.228698e-006, 1.750487e-006, 1.474443e-006, 
    9.346477e-007, 1.960593e-006, 2.736697e-006, 2.544595e-006, 
    1.928184e-006, 2.471332e-006, 2.848703e-006, 2.624192e-006, 2.06366e-006, 
    1.616873e-006, 1.914647e-006, 1.245834e-006, 6.204814e-007, 
    -3.299647e-007, -2.114994e-007, -9.303494e-008, -7.675617e-007, 
    -5.634147e-007, 5.577731e-007, 5.859602e-007, -2.251595e-007, 
    3.896375e-007, 1.533674e-006, 1.222985e-006, 9.896576e-007, 1.6016e-006, 
    2.277119e-006, 2.873164e-006, 3.124746e-006, 2.428615e-006, 
    1.820647e-006, 1.92781e-006, 2.314248e-006, 1.940105e-006, 1.237391e-006, 
    1.760918e-006, 3.062286e-006, 2.595879e-006, 1.487978e-006, 
    1.008037e-006, 5.52558e-007, 1.365661e-007, -2.473917e-008, 
    -3.926743e-008, 7.843955e-007, 1.782898e-006, 1.729377e-006, 
    2.571423e-007, 5.631127e-007, 1.525356e-006, 1.527591e-006, 
    7.416784e-007, 1.138424e-007, -2.773122e-007, 1.184988e-006, 
    2.011506e-006, 2.14512e-006, 3.831308e-006, 4.478143e-006, 2.555274e-006, 
    1.601724e-006, 2.127857e-006, 3.405632e-006, 4.880967e-006, 4.01844e-006, 
    8.375391e-007, 5.283382e-007, 2.066761e-006, 2.59737e-006, 1.928554e-006, 
    1.398821e-006, 1.442407e-006, 1.017723e-006, 2.000826e-006, 1.822632e-006,
  1.165989e-006, 1.519657e-007, -5.298871e-007, -6.310802e-008, 
    7.406861e-007, 9.16767e-007, 1.318725e-006, 6.187447e-007, 
    -1.082935e-008, 1.306071e-007, 6.361279e-007, 4.297472e-007, 
    1.967919e-007, -4.456961e-007, 6.392384e-008, 2.675724e-007, 
    4.062786e-007, 6.540104e-007, 2.01312e-006, 2.404276e-006, 3.120028e-006, 
    2.392603e-006, 2.773204e-006, 3.125368e-006, 2.966545e-006, 
    1.902602e-006, 2.030255e-006, 1.770478e-006, 9.122978e-007, 
    5.422498e-007, 2.49318e-007, 1.694725e-007, 1.08254e-007, 2.234901e-007, 
    1.327171e-007, 2.850816e-007, 5.736674e-007, 7.082745e-007, 
    2.598731e-007, 1.29985e-007, 1.846238e-007, 4.145977e-007, 1.234043e-007, 
    1.530821e-007, 2.408751e-007, 5.428719e-007, 1.150342e-006, 
    8.797615e-007, 1.046159e-006, 1.793453e-006, 1.743656e-006, 
    1.301962e-006, 6.269393e-007, 9.306741e-007, 9.48929e-007, 1.171453e-006, 
    1.56832e-006, 1.66853e-006, 2.336848e-006, 2.351127e-006, 1.393355e-006, 
    1.363677e-006, 1.567948e-006, 1.154689e-006, 9.090672e-007, 
    1.272159e-006, 1.453705e-006, 7.862568e-007, 1.780418e-007, 
    3.510195e-007, 5.410093e-007, 6.143973e-007, 7.817871e-007, 6.66555e-008, 
    1.610283e-007, 5.372835e-007, 1.533551e-006, 2.232539e-006, 
    2.363794e-006, 1.223978e-006, 9.578685e-007, 4.640196e-007, 3.60953e-007, 
    1.772963e-006, 2.34231e-006, 1.514551e-006, 1.171578e-006, 1.046405e-006, 
    9.995947e-007, 2.326045e-006, 2.396703e-006, 2.650391e-006, 
    2.719436e-006, 1.719319e-006, 2.007036e-006, 1.684052e-006,
  9.637051e-007, 4.32975e-007, -8.117668e-007, -7.801018e-007, 1.650033e-007, 
    3.34132e-007, 9.058394e-007, 1.365293e-006, 8.240077e-007, 4.343401e-007, 
    8.277329e-007, 1.547334e-006, 1.948921e-006, 1.700692e-006, 
    1.385781e-006, 1.754211e-006, 2.13059e-006, 1.931287e-006, 2.330017e-006, 
    2.335978e-006, 1.58943e-006, 9.635814e-007, 5.165462e-007, 9.319156e-007, 
    1.174556e-006, 9.597316e-007, 3.056939e-007, 1.114768e-008, 6.34886e-007, 
    1.045289e-006, 1.013376e-006, 3.070616e-007, 2.56025e-007, 5.21514e-007, 
    4.213034e-007, 3.431969e-007, 3.572281e-007, 5.709358e-007, 
    6.988378e-007, 8.037664e-007, 7.305025e-007, 5.067366e-007, 
    5.474669e-007, 7.560827e-007, 6.474281e-007, 5.289644e-007, 
    4.944436e-007, 3.643065e-007, 3.337618e-008, 1.859917e-008, 
    7.013205e-008, 4.679937e-007, 1.082791e-006, 1.199516e-006, 
    1.225842e-006, 1.375846e-006, 1.752225e-006, 2.166601e-006, 
    2.143505e-006, 1.658969e-006, 1.01201e-006, 5.85713e-007, 5.840989e-007, 
    4.956851e-007, -1.393437e-008, -6.014134e-007, -5.374632e-007, 
    7.870085e-008, 3.412097e-007, 5.788829e-007, 6.247037e-007, 
    -5.987658e-009, 3.824357e-007, 9.131659e-007, 1.052616e-006, 
    1.273028e-006, 2.371617e-006, 2.857395e-006, 1.681569e-006, 
    3.032114e-007, -1.331364e-008, 3.983428e-008, -4.494209e-007, 
    -4.208614e-007, 7.059152e-007, 1.033492e-006, 1.09198e-006, 
    1.094214e-006, 1.745271e-006, 2.990264e-006, 3.112576e-006, 
    2.280347e-006, 1.828718e-006, 2.155675e-006, 1.904466e-006, 1.346292e-006,
  5.429956e-007, 4.666272e-007, 4.74327e-007, 6.486707e-007, 9.810892e-007, 
    1.161021e-006, 6.559958e-007, 2.53789e-007, 1.820154e-007, 1.465005e-007, 
    -1.194894e-008, 4.69111e-007, 1.202248e-006, 1.799785e-006, 
    2.158406e-006, 2.195535e-006, 2.36516e-006, 2.750976e-006, 2.717074e-006, 
    2.366773e-006, 1.644813e-006, 9.982255e-007, 7.039275e-007, 
    7.467684e-007, 7.589383e-007, 4.520984e-007, 2.366523e-007, 
    3.402147e-007, 1.033368e-006, 1.062673e-006, 2.905449e-007, 
    -3.32323e-007, -3.046312e-007, 1.646308e-007, 4.144731e-007, 
    3.407122e-007, 1.994008e-007, 2.573906e-007, 4.13108e-007, 2.070994e-007, 
    -1.697756e-007, -8.359712e-008, -4.249432e-008, -3.280911e-008, 
    2.439797e-007, 4.836402e-007, 4.193168e-007, 1.37064e-007, 1.549456e-007, 
    4.114936e-007, 8.041384e-007, 1.158662e-006, 1.61501e-006, 2.115938e-006, 
    2.345416e-006, 2.28072e-006, 2.10203e-006, 1.794445e-006, 1.640467e-006, 
    1.941346e-006, 2.171445e-006, 2.112833e-006, 1.667661e-006, 1.11756e-006, 
    4.723402e-007, -8.570805e-008, -2.509873e-007, 7.572044e-008, 
    -1.332683e-007, -6.493456e-007, -6.8486e-007, -8.061807e-008, 
    2.901734e-007, 5.567797e-007, 9.70784e-007, 1.073975e-006, 1.416204e-006, 
    1.6694e-006, 1.594522e-006, 1.663688e-006, 1.538393e-006, 6.840605e-007, 
    -1.938674e-007, -4.57369e-007, -2.085187e-007, 2.500644e-007, 
    8.466072e-007, 1.308295e-006, 1.687778e-006, 1.989526e-006, 
    2.150459e-006, 2.169955e-006, 1.980833e-006, 1.561613e-006, 8.31953e-007, 
    6.022269e-007,
  8.437505e-007, 9.216092e-007, 1.085522e-006, 1.397576e-006, 1.623951e-006, 
    1.753963e-006, 1.70156e-006, 1.494187e-006, 1.086764e-006, 6.983405e-007, 
    6.301675e-007, 7.468939e-007, 7.611739e-007, 6.312853e-007, 
    6.369974e-007, 8.920551e-007, 1.252291e-006, 1.655492e-006, 
    1.913033e-006, 1.868703e-006, 1.705162e-006, 1.317236e-006, 
    8.467314e-007, 5.134425e-007, 3.686528e-007, 2.316851e-007, 
    -7.813424e-008, -2.313682e-007, -1.910107e-007, -9.837549e-008, 
    -5.454058e-008, -1.061976e-007, -1.620767e-007, -1.57358e-007, 
    -1.975911e-007, -2.447782e-007, -1.784679e-007, 4.567937e-009, 
    7.410654e-008, 3.014839e-008, 8.056395e-008, 2.175298e-007, 
    2.608676e-007, 2.171578e-007, 2.731613e-007, 4.857513e-007, 
    5.917975e-007, 5.802492e-007, 6.492912e-007, 6.260702e-007, 
    4.307412e-007, 3.361188e-007, 5.108348e-007, 9.922667e-007, 
    1.423655e-006, 1.382304e-006, 1.153075e-006, 1.100548e-006, 
    1.232672e-006, 1.526473e-006, 1.592783e-006, 1.447993e-006, 
    1.186478e-006, 8.233869e-007, 6.443245e-007, 6.958576e-007, 
    7.827807e-007, 7.419264e-007, 6.817008e-007, 5.077295e-007, 
    1.538269e-007, -1.969706e-007, -2.804168e-007, -1.815724e-007, 
    -1.65802e-007, -1.670439e-007, -1.465546e-007, -1.03093e-007, 
    4.778076e-008, 1.8127e-007, 3.256873e-007, 5.196516e-007, 7.226797e-007, 
    7.240455e-007, 6.148944e-007, 5.29212e-007, 5.231275e-007, 5.631127e-007, 
    4.792939e-007, 2.70554e-007, 9.410996e-009, -1.186149e-007, 
    1.282469e-007, 5.165457e-007, 7.739641e-007, 7.90852e-007,
  1.051498e-006, 1.100547e-006, 1.09856e-006, 1.055596e-006, 9.650712e-007, 
    8.754164e-007, 7.876242e-007, 6.735063e-007, 5.708121e-007, 
    4.619096e-007, 2.408751e-007, -5.391985e-008, -3.400219e-007, 
    -5.185875e-007, -5.106399e-007, -3.980117e-007, -2.379488e-007, 
    -8.670168e-008, 4.790536e-008, 1.463764e-007, 2.467114e-007, 
    4.170811e-007, 6.496634e-007, 8.721877e-007, 1.000214e-006, 
    1.013624e-006, 9.747569e-007, 8.740503e-007, 6.896489e-007, 
    4.909671e-007, 3.033363e-007, 1.527101e-007, 4.045478e-008, 
    -7.601557e-009, 1.512285e-008, 2.369097e-008, -1.418289e-008, 
    -8.34732e-008, -1.219678e-007, -1.577307e-007, -1.754875e-007, 
    -1.378626e-007, -8.086545e-008, -3.130936e-009, 1.063922e-007, 
    2.31686e-007, 3.682803e-007, 5.523093e-007, 7.63037e-007, 8.890761e-007, 
    8.591496e-007, 7.642789e-007, 7.303786e-007, 8.138252e-007, 
    9.407333e-007, 1.071615e-006, 1.151957e-006, 1.175302e-006, 
    1.168721e-006, 1.218516e-006, 1.300844e-006, 1.384167e-006, 
    1.436073e-006, 1.41012e-006, 1.370508e-006, 1.381931e-006, 1.397205e-006, 
    1.380565e-006, 1.316118e-006, 1.226091e-006, 1.124763e-006, 
    9.928874e-007, 8.570385e-007, 8.025249e-007, 8.046359e-007, 
    8.213997e-007, 8.509537e-007, 9.078265e-007, 9.182572e-007, 
    8.472284e-007, 7.713568e-007, 8.048844e-007, 8.883305e-007, 
    9.792277e-007, 9.665619e-007, 8.196612e-007, 6.091825e-007, 4.41172e-007, 
    3.604573e-007, 3.400924e-007, 3.431969e-007, 3.148848e-007, 
    2.524239e-007, 3.767232e-007, 6.526434e-007, 9.113028e-007,
  1.892172e-007, 1.469975e-007, 1.265084e-007, 1.411613e-007, 1.831331e-007, 
    2.542861e-007, 3.433206e-007, 4.453927e-007, 5.546681e-007, 
    6.710216e-007, 7.987992e-007, 9.375044e-007, 1.08279e-006, 1.23677e-006, 
    1.384291e-006, 1.519271e-006, 1.634258e-006, 1.724782e-006, 
    1.776688e-006, 1.786001e-006, 1.756323e-006, 1.688523e-006, 
    1.591665e-006, 1.473201e-006, 1.342816e-006, 1.210941e-006, 
    1.084654e-006, 9.618429e-007, 8.550514e-007, 7.640306e-007, 
    6.823223e-007, 6.081889e-007, 5.359184e-007, 4.60916e-007, 3.815674e-007, 
    2.974998e-007, 2.195172e-007, 1.592916e-007, 1.160781e-007, 
    8.640018e-008, 6.690402e-008, 5.746665e-008, 5.436254e-008, 
    6.417235e-008, 9.024916e-008, 1.335868e-007, 1.956751e-007, 
    2.778797e-007, 3.662933e-007, 4.466353e-007, 5.24494e-007, 5.92046e-007, 
    6.424616e-007, 6.656826e-007, 6.663035e-007, 6.489188e-007, 
    6.232144e-007, 5.950262e-007, 5.752822e-007, 5.690736e-007, 
    5.804977e-007, 6.088101e-007, 6.473047e-007, 6.815771e-007, 
    7.041774e-007, 7.083993e-007, 7.019423e-007, 7.002038e-007, 
    7.129941e-007, 7.277711e-007, 7.324895e-007, 7.281435e-007, 
    7.086478e-007, 6.814532e-007, 6.550033e-007, 6.440762e-007, 
    6.507814e-007, 6.761134e-007, 7.194512e-007, 7.825329e-007, 
    8.590252e-007, 9.445828e-007, 1.035603e-006, 1.117933e-006, 
    1.177538e-006, 1.199392e-006, 1.167231e-006, 1.084033e-006, 
    9.650719e-007, 8.278569e-007, 6.860478e-007, 5.509437e-007, 
    4.329763e-007, 3.456803e-007, 2.857032e-007, 2.351626e-007,
  6.838118e-007, 7.206922e-007, 7.540957e-007, 7.812904e-007, 8.036423e-007, 
    8.201575e-007, 8.277325e-007, 8.289742e-007, 8.179223e-007, 
    8.024005e-007, 7.811662e-007, 7.612979e-007, 7.430442e-007, 7.26156e-007, 
    7.067845e-007, 6.840603e-007, 6.609636e-007, 6.348864e-007, 6.04215e-007, 
    5.713082e-007, 5.333103e-007, 4.981683e-007, 4.653857e-007, 
    4.353352e-007, 4.14225e-007, 4.037944e-007, 4.030493e-007, 4.093823e-007, 
    4.272636e-007, 4.462627e-007, 4.631506e-007, 4.792936e-007, 
    4.948156e-007, 5.14808e-007, 5.376564e-007, 5.618707e-007, 5.891895e-007, 
    6.189919e-007, 6.510294e-007, 6.905175e-007, 7.355934e-007, 
    7.868783e-007, 8.433788e-007, 9.026107e-007, 9.622152e-007, 1.02182e-006, 
    1.082542e-006, 1.142147e-006, 1.190824e-006, 1.229567e-006, 
    1.253533e-006, 1.257134e-006, 1.240619e-006, 1.207588e-006, 
    1.157048e-006, 1.086392e-006, 9.978539e-007, 8.960292e-007, 
    7.924662e-007, 6.8791e-007, 5.95895e-007, 5.171673e-007, 4.568178e-007, 
    4.210547e-007, 4.123626e-007, 4.383151e-007, 4.939466e-007, 5.72426e-007, 
    6.60094e-007, 7.454037e-007, 8.23386e-007, 8.941665e-007, 9.530261e-007, 
    1.000834e-006, 1.036224e-006, 1.054851e-006, 1.047028e-006, 1.01884e-006, 
    9.728944e-007, 9.185051e-007, 8.59894e-007, 7.975575e-007, 7.341032e-007, 
    6.631988e-007, 5.919214e-007, 5.325653e-007, 4.882343e-007, 
    4.650133e-007, 4.537133e-007, 4.540857e-007, 4.678693e-007, 4.89476e-007, 
    5.210168e-007, 5.581455e-007, 5.991237e-007, 6.410953e-007,
  1.228077e-006, 1.264336e-006, 1.290413e-006, 1.28259e-006, 1.225345e-006, 
    1.139167e-006, 1.023062e-006, 8.929247e-007, 7.62788e-007, 6.453171e-007, 
    5.401399e-007, 4.569417e-007, 4.050359e-007, 3.834293e-007, 
    3.893897e-007, 4.014348e-007, 4.217997e-007, 4.53713e-007, 4.878615e-007, 
    5.092199e-007, 5.182848e-007, 5.190299e-007, 5.083507e-007, 
    4.892275e-007, 4.676208e-007, 4.488701e-007, 4.333481e-007, 
    4.227932e-007, 4.18447e-007, 4.077678e-007, 3.934875e-007, 3.836777e-007, 
    3.785864e-007, 3.732467e-007, 3.770963e-007, 4.005656e-007, 
    4.168327e-007, 4.2627e-007, 4.614121e-007, 5.369113e-007, 6.206061e-007, 
    6.92256e-007, 7.307507e-007, 7.241691e-007, 6.872888e-007, 6.533887e-007, 
    6.589767e-007, 7.441618e-007, 9.24093e-007, 1.187347e-006, 1.444765e-006, 
    1.665426e-006, 1.849703e-006, 1.947555e-006, 1.904341e-006, 
    1.780165e-006, 1.558883e-006, 1.214666e-006, 8.355555e-007, 4.76934e-007, 
    2.49443e-007, 2.239867e-007, 3.160017e-007, 4.549552e-007, 6.157634e-007, 
    7.843946e-007, 9.171395e-007, 1.012383e-006, 1.05659e-006, 1.012382e-006, 
    9.208645e-007, 8.878335e-007, 9.291844e-007, 9.860571e-007, 
    1.025918e-006, 1.035479e-006, 1.019585e-006, 1.055099e-006, 1.1455e-006, 
    1.23143e-006, 1.302086e-006, 1.379572e-006, 1.446627e-006, 1.451967e-006, 
    1.427628e-006, 1.390872e-006, 1.350515e-006, 1.309288e-006, 
    1.279982e-006, 1.289668e-006, 1.319471e-006, 1.332261e-006, 
    1.299975e-006, 1.25403e-006, 1.215783e-006, 1.209078e-006,
  1.095705e-006, 8.589006e-007, 7.446583e-007, 7.121241e-007, 7.214375e-007, 
    7.128692e-007, 6.548788e-007, 5.582696e-007, 4.725878e-007, 
    4.031733e-007, 3.409609e-007, 2.753959e-007, 1.965438e-007, 
    1.623953e-007, 2.084648e-007, 2.633507e-007, 3.228312e-007, 
    3.813182e-007, 4.588043e-007, 5.083507e-007, 5.095924e-007, 
    4.667516e-007, 3.814424e-007, 3.217136e-007, 3.141389e-007, 3.4034e-007, 
    4.010623e-007, 4.73333e-007, 5.19154e-007, 5.271013e-007, 5.3182e-007, 
    5.388981e-007, 5.06488e-007, 4.338448e-007, 3.795798e-007, 3.618226e-007, 
    3.674105e-007, 3.815666e-007, 4.046634e-007, 3.984546e-007, 
    3.313995e-007, 2.700564e-007, 2.727882e-007, 2.455938e-007, 
    2.133079e-007, 1.977855e-007, 1.652515e-007, 2.664551e-007, 
    5.505708e-007, 1.073974e-006, 1.769858e-006, 2.326788e-006, 
    2.390491e-006, 2.070365e-006, 1.511819e-006, 1.127121e-006, 
    8.972711e-007, 6.088094e-007, 4.342173e-007, 3.388495e-007, 
    4.287522e-007, 6.651844e-007, 9.081987e-007, 1.198647e-006, 
    1.394846e-006, 1.332509e-006, 1.19368e-006, 1.132337e-006, 1.103031e-006, 
    8.546785e-007, 5.089719e-007, 3.297851e-007, 3.888931e-007, 
    7.164704e-007, 1.144879e-006, 1.589057e-006, 2.068006e-006, 
    2.463135e-006, 2.577129e-006, 2.546084e-006, 2.35299e-006, 2.069247e-006, 
    1.975493e-006, 2.10501e-006, 2.321946e-006, 2.592775e-006, 2.779784e-006, 
    2.805613e-006, 2.797541e-006, 2.696959e-006, 2.42849e-006, 2.051242e-006, 
    1.810712e-006, 1.766381e-006, 1.692124e-006, 1.438804e-006,
  1.240991e-006, 1.087882e-006, 8.247521e-007, 5.678312e-007, 5.403883e-007, 
    5.391464e-007, 4.636472e-007, 4.49988e-007, 4.328515e-007, 4.304922e-007, 
    4.442758e-007, 3.854161e-007, 2.69808e-007, 2.552794e-007, 2.869444e-007, 
    2.880619e-007, 3.011005e-007, 2.400056e-007, 2.264705e-007, 2.57763e-007, 
    2.99362e-007, 3.732468e-007, 5.087232e-007, 6.198612e-007, 6.46559e-007, 
    5.90928e-007, 5.427477e-007, 5.603806e-007, 6.484217e-007, 7.204439e-007, 
    7.328616e-007, 7.497496e-007, 7.49998e-007, 7.152286e-007, 6.412195e-007, 
    6.23959e-007, 7.277703e-007, 6.569899e-007, 5.06364e-007, 4.057812e-007, 
    5.551652e-007, 7.355936e-007, 8.163081e-007, 8.493391e-007, 
    1.100299e-006, 1.646676e-006, 2.062418e-006, 2.314e-006, 2.487721e-006, 
    2.030504e-006, 1.403786e-006, 1.043178e-006, 1.046034e-006, 1.33884e-006, 
    1.54249e-006, 1.327539e-006, 1.044294e-006, 8.472261e-007, 8.092293e-007, 
    1.412602e-006, 2.149091e-006, 2.315859e-006, 1.682063e-006, 
    3.854148e-007, -9.740688e-007, -1.370192e-006, -5.161055e-007, 
    1.078939e-006, 2.744391e-006, 3.831929e-006, 3.80523e-006, 3.574636e-006, 
    4.113312e-006, 4.612004e-006, 4.922445e-006, 5.212893e-006, 
    5.062144e-006, 4.725626e-006, 4.392461e-006, 3.988639e-006, 
    3.545701e-006, 3.13443e-006, 2.73421e-006, 2.658462e-006, 3.161749e-006, 
    3.491809e-006, 3.399671e-006, 2.957852e-006, 2.320828e-006, 
    1.938987e-006, 1.81332e-006, 2.009767e-006, 2.086508e-006, 1.837162e-006, 
    1.638231e-006, 1.422413e-006,
  4.540605e-006, 2.844728e-006, 1.643571e-006, 1.273526e-006, 1.281721e-006, 
    1.357593e-006, 1.421419e-006, 1.513806e-006, 1.261232e-006, 
    9.433404e-007, 1.013997e-006, 1.226587e-006, 1.120043e-006, 
    7.640299e-007, 5.646025e-007, 4.930771e-007, 3.731228e-007, 
    4.097548e-007, 5.203959e-007, 7.590629e-007, 9.824562e-007, 
    1.323941e-006, 1.652139e-006, 1.617246e-006, 1.475188e-006, 
    1.344554e-006, 1.079438e-006, 1.091234e-006, 1.25018e-006, 1.379821e-006, 
    1.371749e-006, 1.145003e-006, 1.110606e-006, 1.51629e-006, 1.863984e-006, 
    2.248806e-006, 2.443018e-006, 2.154557e-006, 1.7824e-006, 1.501141e-006, 
    1.43334e-006, 1.62718e-006, 1.677844e-006, 1.322078e-006, 1.292897e-006, 
    1.788111e-006, 3.181617e-006, 4.115673e-006, 4.256861e-006, 
    3.807094e-006, 2.079303e-006, 4.955591e-007, -3.385321e-007, 
    2.840716e-008, 1.100299e-006, 9.480573e-007, 1.176668e-006, 1.71584e-006, 
    1.388014e-006, 1.093096e-006, 1.869943e-006, 3.023666e-006, 
    2.670011e-006, 1.152452e-006, 4.194226e-008, 3.803234e-007, 
    2.005791e-006, 3.706511e-006, 3.476038e-006, 3.041545e-006, 
    2.582094e-006, 1.77768e-006, 3.457537e-006, 5.80596e-006, 6.173397e-006, 
    6.322658e-006, 6.587278e-006, 5.902569e-006, 4.39097e-006, 3.073584e-006, 
    2.44997e-006, 2.528822e-006, 2.791579e-006, 3.674597e-006, 4.829065e-006, 
    6.059032e-006, 5.499369e-006, 4.539237e-006, 3.961693e-006, 
    3.810322e-006, 3.937851e-006, 4.030238e-006, 4.212529e-006, 
    4.214764e-006, 4.633612e-006, 5.137147e-006,
  3.838137e-006, 2.519881e-006, 2.490948e-006, 2.684911e-006, 3.021181e-006, 
    3.405383e-006, 3.620456e-006, 4.469947e-006, 4.255991e-006, 
    3.710112e-006, 3.599471e-006, 3.922826e-006, 5.192031e-006, 5.25114e-006, 
    3.917238e-006, 2.732225e-006, 2.175666e-006, 1.591541e-006, 
    1.599488e-006, 1.892917e-006, 2.371989e-006, 2.718813e-006, 
    2.667527e-006, 3.096059e-006, 3.592765e-006, 2.35212e-006, 1.745393e-006, 
    1.494433e-006, 2.356217e-006, 3.366888e-006, 3.458655e-006, 
    3.356953e-006, 3.987521e-006, 4.162735e-006, 4.837881e-006, 
    6.147817e-006, 5.435666e-006, 3.713836e-006, 3.109099e-006, 
    3.390729e-006, 4.00888e-006, 3.960575e-006, 2.865589e-006, 1.871307e-006, 
    1.618733e-006, 2.604695e-006, 2.596003e-006, 1.764271e-006, 
    2.329271e-006, 2.106499e-006, 2.01225e-006, 2.751223e-006, 3.400664e-006, 
    3.718431e-006, 2.702172e-006, 1.283706e-006, 8.320776e-007, 
    7.281424e-007, 2.220866e-006, 3.379306e-006, 3.199624e-006, 
    1.922223e-006, 3.569175e-006, 4.432571e-006, 3.835281e-006, 
    3.468715e-006, 3.024783e-006, 2.608418e-006, 1.970277e-006, 
    3.183108e-006, 4.11741e-006, 3.971627e-006, 4.534269e-006, 4.390475e-006, 
    4.24705e-006, 5.227547e-006, 5.818752e-006, 4.718549e-006, 3.232655e-006, 
    2.881112e-006, 2.870433e-006, 3.185467e-006, 2.968778e-006, 
    3.236752e-006, 3.67733e-006, 4.120887e-006, 3.732836e-006, 3.036331e-006, 
    2.856524e-006, 2.581473e-006, 2.98815e-006, 3.928663e-006, 4.627155e-006, 
    4.310382e-006, 3.872783e-006, 4.577609e-006,
  4.815529e-006, 4.599462e-006, 3.211542e-006, 3.584075e-006, 5.696436e-006, 
    5.742257e-006, 5.420021e-006, 5.491422e-006, 5.210908e-006, 
    4.614116e-006, 4.387246e-006, 6.410326e-006, 8.830277e-006, 
    9.944762e-006, 9.464695e-006, 8.454394e-006, 7.19214e-006, 7.666495e-006, 
    8.078139e-006, 7.616203e-006, 6.05332e-006, 4.789702e-006, 4.576739e-006, 
    4.86694e-006, 4.594622e-006, 4.87228e-006, 4.07134e-006, 3.38775e-006, 
    3.851052e-006, 4.522844e-006, 6.108205e-006, 6.273111e-006, 
    5.570273e-006, 6.300557e-006, 8.049956e-006, 9.285639e-006, 
    8.462095e-006, 8.488423e-006, 7.094794e-006, 6.811548e-006, 
    5.815902e-006, 2.399309e-006, 1.281845e-006, 3.150824e-006, 
    3.721538e-006, 4.602944e-006, 4.045763e-006, 2.492689e-006, 
    2.637977e-006, 3.865085e-006, 3.458656e-006, 2.702422e-006, 
    3.663794e-006, 5.361037e-006, 5.631244e-006, 3.970261e-006, 
    3.248921e-006, 3.698564e-006, 5.70277e-006, 5.292366e-006, 3.403273e-006, 
    1.880993e-006, 3.89352e-006, 4.775295e-006, 5.138139e-006, 5.964161e-006, 
    5.428215e-006, 5.744119e-006, 5.781498e-006, 4.687876e-006, 
    5.037806e-006, 6.071201e-006, 6.55226e-006, 4.572392e-006, 3.214771e-006, 
    4.047126e-006, 4.307276e-006, 3.679688e-006, 4.182602e-006, 
    2.727629e-006, 1.09533e-006, 2.389123e-006, 4.301315e-006, 3.271025e-006, 
    2.422652e-006, 1.808847e-006, 1.401177e-006, 1.515667e-006, 
    7.282651e-007, 3.957202e-007, 6.238342e-007, 1.218018e-006, 
    1.797797e-006, 2.917493e-006, 3.500999e-006, 4.302311e-006,
  2.898869e-006, 2.928173e-006, 4.333724e-006, 5.140624e-006, 4.402644e-006, 
    4.184714e-006, 5.988872e-006, 7.978302e-006, 7.905906e-006, 
    7.266523e-006, 7.828545e-006, 7.929002e-006, 6.824461e-006, 
    6.495264e-006, 7.43553e-006, 9.925883e-006, 1.051001e-005, 1.060637e-005, 
    1.195927e-005, 1.19173e-005, 1.002448e-005, 7.858844e-006, 6.826442e-006, 
    6.450437e-006, 4.810563e-006, 6.450437e-006, 5.598338e-006, 
    5.271011e-006, 6.218601e-006, 7.990226e-006, 9.988842e-006, 
    8.367226e-006, 3.704648e-006, 3.652003e-006, 5.262198e-006, 
    5.939826e-006, 6.04165e-006, 6.06785e-006, 5.36464e-006, 6.164335e-006, 
    5.924676e-006, 6.016564e-006, 5.175019e-006, 4.663043e-006, 
    6.984645e-006, 7.99072e-006, 6.270257e-006, 2.496414e-006, 1.491579e-006, 
    1.897759e-006, 2.62233e-006, 2.308039e-006, 3.520867e-006, 4.496023e-006, 
    4.958207e-006, 3.299958e-006, 3.139894e-006, 5.61448e-006, 5.77504e-006, 
    2.915134e-006, 1.774079e-006, 1.95103e-006, 4.994095e-006, 3.541232e-006, 
    2.914016e-006, 4.011486e-006, 4.534766e-006, 4.141377e-006, 
    5.447839e-006, 7.409453e-006, 6.25461e-006, 5.083626e-006, 6.575854e-006, 
    7.364746e-006, 4.616104e-006, 3.27624e-006, 2.986289e-006, 2.139903e-006, 
    2.348768e-006, 1.697712e-006, 8.063726e-007, 8.552979e-007, 
    1.285322e-006, 8.356783e-007, 1.872104e-008, 7.749568e-007, 1.5035e-006, 
    1.838154e-006, 1.919861e-006, 1.797176e-006, 1.798913e-006, 
    1.940847e-006, 2.262464e-006, 1.832441e-006, 2.211924e-006, 2.893157e-006,
  6.426595e-006, 6.25635e-006, 5.649252e-006, 5.792803e-006, 5.459262e-006, 
    5.092323e-006, 4.995964e-006, 5.208301e-006, 3.878373e-006, 
    5.140875e-006, 5.182472e-006, 5.696438e-006, 7.311974e-006, 
    7.558585e-006, 7.541326e-006, 7.870643e-006, 8.438627e-006, 
    9.211126e-006, 8.512387e-006, 6.377051e-006, 6.379287e-006, 
    5.025766e-006, 4.574878e-006, 5.960685e-006, 5.672226e-006, 
    6.443486e-006, 6.914735e-006, 6.135402e-006, 5.312364e-006, 
    3.738922e-006, 3.100908e-006, 4.841115e-006, 6.129691e-006, 
    5.893631e-006, 2.470337e-006, 1.977856e-006, 4.511796e-006, 
    4.578604e-006, 4.299825e-006, 4.890411e-006, 5.014586e-006, 
    6.188919e-006, 6.939072e-006, 7.787319e-006, 7.770062e-006, 
    8.853873e-006, 9.497227e-006, 7.965762e-006, 5.575241e-006, 
    4.765488e-006, 4.812053e-006, 4.680176e-006, 4.904812e-006, 
    5.598089e-006, 7.036548e-006, 3.96691e-006, 2.371242e-006, 2.690873e-006, 
    4.007392e-006, 3.146102e-006, 2.259236e-006, 6.428831e-006, 
    7.552748e-006, 5.153413e-006, 5.054568e-006, 8.230008e-006, 
    8.999283e-006, 6.369599e-006, 4.922571e-006, 4.190924e-006, 
    4.988759e-006, 4.361043e-006, 5.414064e-006, 5.083999e-006, 
    6.041151e-006, 4.15777e-006, 2.472574e-006, 2.07049e-006, 1.53355e-006, 
    7.097624e-007, 1.234906e-006, 3.79741e-006, 3.718556e-006, 2.256627e-006, 
    1.179396e-007, -3.262394e-007, 1.021694e-006, 2.823368e-006, 3.8251e-006, 
    4.881593e-006, 2.640583e-006, 6.609644e-007, 2.597866e-006, 
    4.568421e-006, 4.996333e-006, 5.825084e-006,
  5.832037e-006, 5.339185e-006, 2.901976e-006, 2.2118e-006, 4.607533e-006, 
    5.520356e-006, 4.593134e-006, 5.631744e-006, 7.278319e-006, 
    8.800474e-006, 7.927891e-006, 7.882569e-006, 9.036532e-006, 8.22057e-006, 
    5.91487e-006, 5.682286e-006, 7.160976e-006, 6.988994e-006, 5.424616e-006, 
    3.873527e-006, 3.693847e-006, 4.088106e-006, 3.604437e-006, 
    3.735448e-006, 4.352351e-006, 5.18719e-006, 6.797018e-006, 5.472793e-006, 
    3.880854e-006, 3.736692e-006, 7.082373e-006, 8.391686e-006, 
    5.360045e-006, 3.838886e-006, 4.334353e-006, 5.461497e-006, 
    6.104357e-006, 5.845453e-006, 4.371479e-006, 4.838876e-006, 
    4.114558e-006, 4.479014e-006, 6.788816e-006, 8.120609e-006, 
    1.034026e-005, 8.680772e-006, 6.059407e-006, 6.502962e-006, 
    3.222847e-006, 3.298219e-006, 4.364523e-006, 6.673336e-006, 
    4.926173e-006, 4.671116e-006, 5.833159e-006, 3.716945e-006, 
    5.218484e-006, 6.139127e-006, 3.202729e-006, 3.056201e-006, 
    7.037792e-006, 8.676299e-006, 6.818622e-006, 4.362162e-006, 
    6.245424e-006, 6.262682e-006, 6.250635e-006, 5.462864e-006, 
    3.843848e-006, 4.710728e-006, 5.087855e-006, 2.975114e-006, 
    5.414186e-006, 9.501946e-006, 8.325009e-006, 4.720292e-006, 
    2.924084e-006, 2.692861e-006, 2.481762e-006, 1.43905e-006, 1.370257e-006, 
    4.853773e-007, 1.140283e-006, 2.342436e-006, 3.587551e-006, 
    3.843106e-006, 1.712117e-006, 9.291816e-007, 1.159657e-006, 
    9.658143e-007, 1.446999e-006, 3.456418e-006, 4.670866e-006, 
    4.582207e-006, 4.862346e-006, 4.724634e-006,
  2.961704e-006, 3.528196e-006, 5.413691e-006, 8.562554e-006, 9.591604e-006, 
    5.244314e-006, 3.69559e-006, 5.883077e-006, 6.80385e-006, 5.993097e-006, 
    7.105344e-006, 6.833397e-006, 8.286883e-006, 1.042867e-005, 
    1.140023e-005, 7.816507e-006, 6.099643e-006, 5.776656e-006, 
    5.296592e-006, 6.056551e-006, 7.214992e-006, 6.797014e-006, 5.15491e-006, 
    4.666021e-006, 4.501242e-006, 4.420031e-006, 6.023645e-006, 
    7.557966e-006, 9.493255e-006, 1.020987e-005, 8.805815e-006, 
    8.185554e-006, 5.774422e-006, 7.044993e-006, 7.970975e-006, 
    8.122224e-006, 4.774305e-006, 3.043166e-006, 2.47543e-006, 8.621282e-007, 
    1.815679e-006, 2.71422e-006, 3.003674e-006, 1.439796e-006, 4.223457e-006, 
    4.872529e-006, 4.725005e-006, 5.8267e-006, 4.19465e-006, 2.228193e-006, 
    1.736953e-006, 3.804238e-006, 2.441653e-006, 1.716711e-006, 
    3.019941e-006, 3.391971e-006, 3.740413e-006, 5.175396e-006, 
    3.789217e-006, 3.362424e-006, 6.064372e-006, 9.950225e-006, 
    8.657798e-006, 9.036285e-006, 8.169784e-006, 5.686503e-006, 
    5.212398e-006, 8.473271e-006, 7.150171e-006, 4.736678e-006, 
    3.502617e-006, 4.787467e-006, 7.531642e-006, 4.884329e-006, 
    2.199879e-006, 2.514793e-006, 1.592041e-006, 3.025281e-006, 
    3.644052e-006, 2.840132e-006, 1.41049e-006, 1.089124e-006, 1.399192e-006, 
    7.349718e-007, 1.226563e-007, -7.686795e-007, -7.093222e-007, 
    4.667527e-007, 1.245462e-006, 1.916884e-006, 4.835772e-006, 
    4.090714e-006, 3.148834e-006, 4.924314e-006, 4.753321e-006, 3.963927e-006,
  4.014099e-006, 6.28168e-006, 7.529652e-006, 4.31982e-006, 1.610042e-006, 
    4.799269e-006, 4.054211e-006, 7.120743e-006, 5.305781e-006, 
    2.315737e-006, 3.851552e-006, 8.066221e-006, 1.061693e-005, 
    7.395047e-006, 4.857753e-006, 4.542591e-006, 4.620699e-006, 
    2.639714e-006, 6.140253e-007, -2.837696e-007, 2.462017e-006, 
    4.327892e-006, 3.081539e-006, 1.324563e-006, 2.478781e-006, 
    4.621939e-006, 4.191545e-006, 3.765123e-006, 3.011497e-006, -1.1874e-007, 
    -1.110537e-006, -8.402021e-007, 1.963323e-006, 3.330133e-006, 
    1.195047e-006, 6.188202e-009, -1.783446e-007, -5.555921e-007, 
    -4.295507e-007, -1.271837e-007, 1.473445e-006, 4.477273e-006, 
    3.653739e-006, -2.399611e-008, 2.184606e-006, 7.394428e-006, 
    7.705738e-006, 3.243707e-006, -8.025781e-007, -3.195457e-006, 
    -1.581911e-006, 2.331763e-007, 2.07136e-006, 7.413037e-007, 
    -1.256922e-008, -1.123324e-006, 1.563229e-006, 4.57004e-006, 
    3.720423e-006, 3.313122e-006, 2.422526e-006, 3.743397e-006, 
    3.039688e-006, 2.401794e-006, 7.875024e-007, 4.835772e-006, 
    6.582064e-006, 6.04289e-006, 6.865412e-007, 2.107008e-007, 2.91688e-006, 
    4.074078e-006, 4.229169e-006, 3.996589e-006, 3.443383e-006, 
    1.577013e-006, 2.336819e-007, -1.132139e-006, 1.394348e-006, 
    2.62717e-006, 2.920598e-006, 2.04826e-006, 1.018714e-006, -7.623476e-007, 
    -4.041347e-006, -4.53644e-006, -2.643617e-006, 2.773453e-006, 
    4.830436e-006, 4.477402e-006, 4.539863e-006, 2.988403e-006, 
    3.837275e-006, 5.931379e-006, 4.649133e-006, 2.751596e-006,
  6.585789e-006, 8.560317e-006, 5.164842e-006, 1.256143e-006, 1.63848e-006, 
    2.653e-006, 4.759157e-006, 7.230141e-006, 7.633966e-006, 9.823561e-006, 
    1.006223e-005, 9.178095e-006, 7.010973e-006, 3.487961e-006, 
    2.242226e-006, 7.538456e-007, 1.950521e-007, -6.14953e-007, 
    5.457259e-007, 3.486222e-006, 2.337219e-006, -3.105924e-007, 
    -1.41179e-006, -3.608715e-006, -4.962363e-006, -7.50897e-006, 
    -6.706792e-006, -6.178918e-006, -6.067781e-006, -4.014149e-006, 
    -2.74209e-006, -1.692177e-006, -1.317414e-006, -2.198176e-007, 
    -4.726426e-007, 4.312387e-007, 1.371747e-006, -4.350186e-007, 
    -3.397727e-007, 2.328405e-006, 5.412574e-006, 6.300557e-006, 
    4.457284e-006, 3.327772e-006, 4.21092e-006, 3.478155e-006, 3.750847e-006, 
    -2.625384e-007, -1.254208e-006, -1.207765e-006, -1.379998e-006, 
    1.358203e-007, -6.499613e-007, 3.561581e-008, 1.304321e-006, 
    1.370383e-006, 3.224093e-006, 9.630894e-007, -9.782852e-007, 
    1.427881e-006, 2.049383e-006, 3.117857e-007, -2.328823e-006, 
    1.164553e-007, -3.509449e-007, 3.12164e-006, 4.765243e-006, 
    6.616217e-006, 4.72178e-006, 5.533399e-006, 4.632748e-006, 2.959223e-006, 
    -7.496783e-007, -6.68093e-007, -3.984838e-006, -7.386774e-006, 
    -6.402432e-006, -1.368695e-006, 1.768865e-006, 2.104885e-006, 
    2.418681e-006, 1.461403e-006, 6.922564e-007, -1.06981e-006, 
    1.994616e-006, 1.902725e-006, 4.167086e-007, 1.054232e-006, 
    -3.57406e-007, -1.034419e-006, -8.991847e-007, 4.307403e-007, 
    2.381053e-006, 1.96134e-006, 2.52758e-006, 5.413069e-006,
  3.455571e-007, -1.966979e-006, -3.834593e-006, -2.483306e-006, 
    -1.085824e-006, 6.786031e-007, 1.441909e-006, 3.160263e-006, 
    5.921325e-006, 9.425577e-006, 5.571768e-006, 8.166862e-007, 
    5.580223e-007, 7.524832e-007, -2.210862e-006, -1.772401e-006, 
    -4.069661e-006, -8.189709e-007, -8.158677e-007, -1.450904e-006, 
    -3.193843e-006, -3.680616e-006, -4.646956e-006, -7.720691e-006, 
    -9.300093e-006, -9.032739e-006, -5.538664e-006, -5.771e-006, 
    -4.705318e-006, -2.009077e-006, -2.540302e-006, -5.036865e-006, 
    -5.387541e-006, -6.131482e-006, -3.244757e-006, -4.093126e-007, 
    -3.797577e-007, -7.216149e-007, -7.412345e-007, 4.593021e-007, 
    3.493424e-006, 6.322412e-006, 5.992726e-006, 6.190912e-006, 
    4.122754e-006, 5.020545e-006, 3.122143e-006, 8.323295e-007, 
    -1.516095e-006, -3.433997e-006, -4.422567e-006, -5.224498e-006, 
    -7.858278e-006, -1.286611e-006, -1.207445e-008, -7.162012e-006, 
    -3.142428e-006, 6.574919e-007, 8.164352e-007, 1.476928e-006, 
    5.963957e-007, -2.212473e-006, -2.322242e-006, -1.344233e-006, 
    2.394518e-008, -6.148257e-007, 5.752197e-006, 5.242706e-006, 
    6.836879e-006, 3.049743e-006, 2.204106e-006, -6.294154e-006, 
    -3.936908e-006, -5.767521e-006, -6.160666e-006, -3.655157e-006, 
    -2.064207e-006, -5.501282e-006, -3.161313e-006, 4.943176e-007, 
    1.023187e-006, -1.428307e-007, 2.466611e-006, 5.129701e-006, 
    7.248145e-006, 4.658326e-006, 5.267037e-006, 4.141377e-006, 
    1.263834e-007, -1.88639e-006, -3.081714e-006, -3.009191e-006, 
    9.476935e-007, 1.477427e-006, 1.032131e-006, 1.032e-006,
  -9.580604e-006, -8.2323e-006, -5.826629e-006, -4.75834e-006, 
    -3.647086e-006, -1.967477e-006, -1.764325e-006, -1.94289e-006, 
    7.647723e-007, -1.926273e-007, -6.77869e-006, -5.649184e-006, 
    -4.448275e-006, -8.012508e-006, -9.305431e-006, -9.027401e-006, 
    -8.226589e-006, -6.069271e-006, -2.823921e-006, -1.768531e-007, 
    -1.040129e-006, -3.135719e-007, -3.996021e-006, -4.226866e-006, 
    -1.191005e-006, -7.45953e-007, -1.580916e-006, -1.164677e-006, 
    2.084653e-007, -1.8664e-006, -7.55976e-006, -7.758688e-006, 
    -5.490114e-006, -2.356895e-006, 6.859227e-007, 1.240742e-006, 
    2.803608e-008, 2.137296e-006, 4.624049e-006, 3.984913e-006, 
    4.819999e-006, 8.729319e-006, 1.103527e-005, 1.211014e-005, 
    1.165665e-005, 4.88371e-006, -2.006713e-006, -5.826125e-006, 
    -6.95651e-006, -1.172227e-005, -1.479949e-005, -1.20188e-005, 
    -1.102936e-005, -8.034727e-006, -6.649916e-006, -1.741722e-006, 
    2.051616e-006, -1.406079e-008, -8.195857e-007, -5.072874e-006, 
    -8.447125e-006, -9.144002e-006, -9.69012e-006, -5.397349e-006, 
    -6.591428e-006, 6.976188e-008, 3.097928e-006, -1.694789e-006, 
    -3.027686e-006, -2.713277e-006, -2.174846e-006, -1.194723e-006, 
    3.136411e-007, -4.286718e-006, -3.342857e-006, -3.701227e-006, 
    -4.315156e-006, -3.186145e-006, 9.817086e-007, 1.274642e-006, 
    -1.515236e-007, 6.485443e-007, 1.150216e-006, 6.9007e-006, 9.534357e-006, 
    6.721268e-006, 1.904591e-006, -3.824898e-007, 6.193659e-007, 
    1.502383e-006, 8.74672e-007, -1.412162e-006, -3.496709e-006, 
    -4.163907e-006, -3.012545e-006, -5.485146e-006,
  -7.444771e-006, -5.410267e-006, -4.181295e-006, -5.127767e-006, 
    -3.430896e-006, -7.798553e-007, -4.617159e-007, 4.509793e-007, 
    4.156936e-008, -1.648716e-006, -5.941125e-006, -4.223763e-006, 
    -3.546755e-006, -5.762682e-006, -8.90459e-006, -1.064604e-005, 
    -8.097568e-006, -5.715989e-006, -2.030558e-006, -1.328954e-007, 
    6.728842e-007, 2.307042e-006, 8.447441e-007, 3.138901e-006, 
    3.476534e-006, 3.441022e-006, 4.3978e-006, 7.384497e-007, -2.555827e-006, 
    -5.291182e-006, -5.230584e-006, -2.220922e-006, 1.320957e-006, 
    4.337947e-006, 3.392096e-006, 5.941562e-006, 6.559586e-006, 
    4.071093e-006, 3.993357e-006, 5.062517e-006, 9.417879e-006, 
    1.054789e-005, 8.842446e-006, 4.3084e-006, 3.206333e-006, -1.2665e-006, 
    -2.024968e-006, -7.079194e-006, -1.042513e-005, -1.436114e-005, 
    -1.123165e-005, -3.237794e-006, -3.758843e-006, 2.913031e-006, 
    4.921334e-006, 3.6561e-006, 2.040317e-006, -1.261033e-006, 
    -3.826648e-006, -4.574926e-006, -5.276401e-006, -5.504142e-006, 
    -1.941393e-006, 9.118012e-007, 2.050256e-006, -3.568974e-006, 
    -1.259945e-005, -1.011754e-005, -8.861494e-006, -1.216185e-005, 
    -1.144164e-005, -7.468241e-006, -5.43945e-006, -6.220393e-006, 
    -4.015645e-006, -2.02845e-006, -2.791264e-006, 1.065137e-007, 
    4.605796e-006, 4.237863e-007, 3.164232e-006, 2.0428e-006, 3.285553e-006, 
    4.828322e-006, 4.023037e-006, -4.819558e-007, -3.667948e-006, 
    -1.70137e-006, 7.445324e-007, -1.607614e-006, -1.010078e-006, 
    -2.685216e-006, -4.975031e-006, -6.663331e-006, -8.040821e-006, 
    -9.728625e-006,
  -4.695012e-006, -3.902146e-006, -3.482057e-006, -1.770286e-006, 
    -7.19629e-007, 7.00079e-008, -2.798466e-006, -8.970783e-007, 
    1.556895e-006, -3.888734e-006, -8.307674e-006, -3.295298e-006, 
    -4.079468e-006, -4.792742e-006, -4.518557e-006, -6.59491e-006, 
    -4.921385e-006, -4.861158e-006, -5.654148e-006, 4.920839e-007, 
    4.020554e-006, 6.840583e-007, -4.681715e-007, 7.810413e-007, 
    -2.294684e-006, -4.026078e-007, -2.322251e-006, -4.338874e-006, 
    -3.085563e-006, -1.396389e-006, -8.549832e-007, 2.653496e-006, 
    5.252756e-006, 5.704509e-006, 6.675569e-006, 4.76524e-006, 4.702777e-006, 
    6.468813e-006, 5.243069e-006, 3.888057e-006, 3.087118e-006, 4.22023e-006, 
    1.71423e-006, -3.489507e-006, -5.015139e-006, -4.64683e-006, 
    -5.501286e-006, -3.99565e-006, -1.112349e-005, -1.057501e-005, 
    -2.570843e-006, -6.001683e-007, 5.57661e-006, 7.672956e-006, 
    6.801984e-006, 1.025508e-005, 8.501338e-006, 1.6206e-006, 1.101667e-006, 
    -4.634785e-008, 2.899986e-006, 9.428808e-006, 9.422598e-006, 
    3.466233e-006, -3.67465e-006, -1.080908e-005, -1.412421e-005, 
    -1.416818e-005, -1.353277e-005, -7.988418e-006, -4.820677e-006, 
    -3.53297e-006, -2.145671e-006, -4.217057e-006, -7.873059e-007, 
    -4.93008e-007, -9.558125e-007, 7.512399e-007, 2.98095e-006, 
    -3.261766e-006, -5.570819e-007, -1.832872e-006, -3.450641e-006, 
    -3.769277e-006, -3.015901e-006, -4.809752e-006, -6.735727e-006, 
    -1.111284e-006, -6.170594e-007, -2.911216e-006, -1.304625e-006, 
    -2.909728e-006, -3.546005e-006, -5.818312e-006, -6.675004e-006, 
    -5.702828e-006,
  -2.199316e-006, -1.544533e-006, -4.322851e-007, -8.127612e-007, 
    -3.082289e-008, -5.852703e-007, -9.036589e-007, -1.039259e-006, 
    8.665211e-009, 2.818529e-007, -3.845646e-006, -3.739724e-006, 
    -9.645055e-007, -1.681379e-006, -2.793251e-006, -5.074991e-006, 
    -2.106184e-006, -2.192983e-006, -4.85059e-007, 1.877641e-006, 
    4.522723e-006, 1.49816e-006, 1.426011e-006, -1.234837e-006, 
    1.099925e-007, 2.724155e-007, -9.181895e-007, -3.022355e-006, 
    -4.668687e-006, -2.097864e-006, 3.686509e-007, 3.118535e-006, 
    5.016464e-007, 1.0849e-006, 2.426998e-006, 4.540355e-006, 6.933356e-006, 
    6.326135e-006, 3.697944e-006, 1.793698e-006, 4.278845e-007, 
    -3.378866e-006, -2.98026e-006, -3.651805e-006, -4.174342e-006, 
    -4.573569e-006, -4.939142e-006, -9.23167e-006, -1.219898e-005, 
    -2.797842e-006, 1.234042e-006, 3.394744e-007, 4.66255e-006, 
    1.116479e-005, 1.046754e-005, 8.898573e-006, 3.766367e-006, 
    3.963432e-006, 8.470663e-006, 1.050343e-005, 1.39831e-005, 1.071888e-005, 
    1.676974e-006, -4.199177e-006, -9.302199e-006, -1.025675e-005, 
    -8.207217e-006, -6.527109e-006, -2.900289e-006, -1.453761e-006, 
    1.165718e-007, -7.46586e-008, -7.786148e-007, -6.931814e-007, 
    -4.432127e-007, 2.580236e-009, 2.629804e-008, 3.49206e-006, 
    9.357655e-007, -4.037372e-006, -5.564247e-006, -1.047616e-005, 
    -7.747887e-006, -6.04779e-006, -2.229615e-006, -1.006974e-006, 
    -3.742578e-006, 5.010224e-007, 2.105879e-006, 1.672503e-006, 
    9.563792e-007, -2.118741e-007, -1.312945e-006, -2.074767e-006, 
    -2.558558e-006, -1.601283e-006,
  1.574263e-007, -4.553831e-007, -2.074016e-007, -2.903516e-007, 
    5.076078e-008, -3.303364e-007, -1.738744e-006, -1.357026e-006, 
    -1.037894e-006, -2.19733e-006, -4.112127e-006, -3.868743e-006, 
    -1.960773e-006, -3.07861e-006, -6.349415e-006, -3.802308e-006, 
    -2.178578e-006, -3.095247e-006, 8.46856e-007, 3.17752e-006, 
    1.567325e-006, 1.883353e-006, 2.513798e-006, 1.756944e-006, 6.23772e-006, 
    -4.121684e-007, -1.43625e-006, -1.398748e-006, -4.052028e-006, 
    2.222603e-006, 5.988253e-006, -7.325452e-007, 2.405027e-007, 
    2.762772e-006, 2.92147e-006, 9.920172e-007, 2.244211e-006, 2.547451e-006, 
    1.611781e-006, -1.19535e-006, -2.536827e-006, -1.24713e-006, 
    1.175425e-006, 1.734219e-006, 3.396075e-006, 1.772591e-006, 
    -6.201626e-007, -1.195596e-006, -9.398187e-006, -1.225673e-005, 
    -1.185725e-005, -2.082335e-006, 9.098123e-006, 1.211685e-005, 
    8.87796e-006, 7.794395e-006, 1.386997e-005, 1.39749e-005, 1.003181e-005, 
    1.223023e-005, 6.43119e-006, -1.304501e-006, -5.725304e-006, 
    -6.360217e-006, -2.268107e-006, 4.56319e-007, -9.400428e-007, 
    -1.522685e-007, -1.277555e-006, -2.231104e-006, -1.536463e-006, 
    -9.488613e-007, -1.212611e-006, -9.85739e-007, 7.460289e-008, 
    1.188216e-006, 2.67349e-006, 1.807111e-006, -3.318765e-006, 
    -1.140029e-005, -8.173565e-006, -6.834694e-006, -3.37986e-006, 
    -2.912708e-006, -2.183048e-006, -2.250476e-006, -2.349074e-006, 
    1.363427e-006, 2.788101e-006, 4.059546e-006, 1.974498e-006, 
    2.954746e-006, 1.476552e-006, -1.485054e-006, -2.794259e-007, 
    -1.078997e-006,
  -1.577317e-006, -7.218655e-007, -3.227617e-007, 1.43893e-007, 
    2.965058e-007, -7.6396e-007, -1.02858e-006, -5.58324e-007, 
    -1.464811e-006, -1.881052e-006, -3.076994e-006, -5.613065e-007, 
    -4.031035e-007, 3.697696e-007, -5.7787e-006, -3.978514e-006, 
    -3.604371e-006, -1.833738e-006, -2.213719e-006, 2.250543e-006, 
    1.479408e-006, 3.071722e-006, 6.629747e-006, 4.466718e-006, 
    8.018287e-006, -1.885521e-006, 2.995728e-006, 6.141732e-006, 
    7.105094e-006, 7.885543e-006, 7.174507e-006, 3.773443e-006, 
    1.251426e-007, 2.886827e-007, 4.76065e-007, 3.038322e-007, 1.21392e-006, 
    1.87665e-006, -1.00114e-007, -2.341994e-006, -2.072904e-006, 
    4.131194e-006, 3.617104e-006, 2.475304e-006, 2.069373e-006, 
    6.090559e-007, 3.588793e-006, -1.734774e-006, -6.588321e-006, 
    7.289251e-006, 6.485334e-006, 1.4262e-005, 1.480887e-005, 1.476553e-005, 
    1.260027e-005, 1.487816e-005, 1.61732e-005, 1.102149e-005, 9.435142e-006, 
    3.619962e-006, -1.085949e-006, -2.413768e-006, -1.850754e-006, 
    4.815265e-007, 8.533116e-007, 4.439016e-007, -1.267373e-006, 
    -1.747067e-006, -2.155855e-006, -2.911965e-006, -1.734772e-006, 
    -2.20627e-006, -1.35802e-006, -5.107645e-007, -2.244142e-007, 
    2.157911e-007, 4.761891e-007, -1.519698e-006, -1.271059e-005, 
    -9.967787e-006, -5.128387e-006, -1.940159e-006, -1.228752e-006, 
    -1.344112e-006, -5.884248e-006, -7.321589e-006, -3.261517e-006, 
    1.246826e-006, 2.162749e-006, -3.690802e-007, 7.483459e-006, 
    6.759137e-006, 1.370008e-006, -8.819297e-007, -1.107559e-006, 
    -6.062583e-007,
  -1.764573e-006, -9.729497e-007, 3.686523e-007, 1.581979e-006, 
    4.147217e-007, -5.360964e-007, -1.535092e-007, -4.496698e-007, 
    -1.222543e-006, -1.635431e-006, -2.86577e-006, -1.05292e-006, 
    -3.752884e-007, -2.036272e-006, -6.50215e-006, -9.095202e-006, 
    -5.977878e-006, -3.798583e-006, 6.152641e-007, 4.351483e-006, 
    2.396826e-006, 4.70936e-006, 7.132539e-006, -2.147281e-007, 
    5.596477e-006, 2.842367e-006, 1.1981e-005, 1.450526e-005, 1.371239e-005, 
    1.741123e-005, 1.200956e-005, 9.49288e-006, 5.537614e-006, 2.377081e-006, 
    7.307508e-007, 9.566272e-007, 1.569189e-006, 2.415202e-006, 
    -1.126679e-006, -9.383057e-007, 4.00056e-006, 4.843843e-006, 
    5.538361e-006, 3.508572e-006, 1.488475e-006, 7.692695e-006, 
    3.112949e-006, 2.144756e-006, 6.264789e-006, 1.083647e-005, 
    1.532086e-005, 1.403066e-005, 1.677173e-005, 1.949516e-005, 
    1.675596e-005, 9.709693e-006, 6.234121e-006, 4.71768e-006, 3.162122e-006, 
    4.308622e-007, 1.576755e-007, -7.690542e-007, -1.593957e-006, 
    -1.334304e-006, -1.930599e-006, -1.140465e-006, -3.132997e-006, 
    -3.638394e-006, -3.27282e-006, -3.443438e-006, -2.395762e-006, 
    -2.098359e-006, -1.968347e-006, -1.236823e-006, -4.305466e-007, 
    1.810247e-008, -3.479947e-006, -7.112974e-006, -4.66074e-006, 
    -3.646715e-006, -3.027447e-006, -6.120922e-007, 4.422886e-007, 
    1.428497e-006, -3.118593e-006, -3.097357e-006, 1.920707e-007, 
    8.179592e-006, 2.237752e-006, 3.579851e-006, 4.231777e-006, 
    -4.423437e-007, 6.409682e-007, -1.219689e-006, 8.206525e-007, 
    -7.255921e-007,
  -6.613909e-007, 1.779176e-007, 3.472689e-006, 4.193034e-006, 3.028387e-007, 
    -2.262539e-009, 1.171952e-007, 1.036599e-007, -3.607595e-007, 
    5.850916e-007, -2.022985e-006, -2.395389e-006, -2.049684e-006, 
    -3.816217e-006, -5.627453e-006, -8.163257e-006, -5.693517e-006, 
    9.285577e-008, -3.389068e-007, -3.807028e-006, -8.3792e-006, 
    3.077061e-006, 1.390363e-005, 6.531282e-006, -3.761823e-006, 
    -3.390531e-006, 1.141054e-005, 1.449347e-005, 1.524312e-005, 
    1.708279e-005, 2.354294e-005, 1.940774e-005, 1.723925e-005, 
    1.402606e-005, 1.231727e-005, 5.451064e-006, 5.417537e-006, 
    4.548428e-006, 2.739674e-006, 1.936453e-005, 2.335754e-005, 1.02829e-005, 
    4.95337e-006, -3.514957e-006, -5.096845e-006, 9.329095e-006, 
    1.82003e-006, 5.51527e-006, 1.569326e-005, 7.202325e-006, -1.439403e-007, 
    7.248389e-006, 4.715577e-006, 8.268013e-006, 1.176767e-005, 
    1.157867e-005, 1.082976e-005, 6.270755e-006, 1.649531e-006, 
    1.308916e-006, -2.788056e-007, -1.82567e-006, -9.938121e-007, 
    -2.225518e-006, -1.955806e-006, -2.253953e-006, -2.346464e-006, 
    -2.556819e-006, -2.43674e-006, -1.850256e-006, -2.155977e-006, 
    -1.944256e-006, -1.99281e-006, -1.93308e-006, -1.281728e-008, 
    1.05547e-006, -2.777606e-006, -3.807151e-006, -1.709438e-006, 
    -3.617905e-006, -1.615562e-006, -5.883749e-007, -4.070789e-007, 
    2.252035e-006, 2.149836e-006, 6.590981e-007, 2.059811e-006, 
    1.304197e-005, 8.973577e-006, 9.88441e-006, 1.105974e-005, 7.598695e-006, 
    3.680061e-006, 2.628522e-007, 1.716213e-006, 2.968764e-007,
  4.226189e-006, 4.902206e-006, 3.814916e-006, 3.260968e-006, 1.445758e-006, 
    1.029271e-006, 1.276009e-006, 1.114952e-006, 3.266806e-007, 
    -6.86598e-007, -2.882285e-006, -5.39487e-006, -3.859804e-006, 
    -5.199541e-006, -6.767264e-006, -7.166122e-006, -5.79633e-006, 
    -2.679506e-006, -3.417361e-006, -9.933392e-006, -1.550245e-006, 
    5.124111e-006, 4.3043e-006, -5.972783e-006, -2.10776e-005, 
    -1.497482e-005, -1.389308e-006, 1.224478e-006, -1.798348e-006, 
    3.058944e-006, 1.024229e-005, 6.553128e-006, 4.073947e-006, 
    6.016067e-006, 9.341387e-006, 1.441238e-005, 1.343908e-005, 
    3.218324e-005, 1.974078e-005, 1.084082e-005, 2.631617e-005, 
    1.045525e-005, 1.076332e-007, -9.792071e-006, -1.714454e-005, 
    -4.999238e-006, -7.319089e-006, -4.981222e-006, 2.242487e-005, 
    3.228297e-005, 3.3542e-005, 2.511763e-005, 2.162217e-005, 2.778779e-005, 
    2.979062e-005, 2.825406e-005, 1.68594e-005, 1.094276e-005, 6.183083e-006, 
    3.185094e-006, 2.714343e-006, -1.018896e-006, -1.691185e-006, 
    -1.668091e-006, -1.338401e-006, -1.365223e-006, -1.43054e-006, 
    -1.60004e-006, -1.92948e-006, -1.663991e-006, -3.551722e-007, 
    -8.343686e-007, 2.811075e-007, -5.517441e-007, 1.198273e-006, 
    -1.735393e-006, -3.546753e-006, -5.582024e-007, -3.641997e-006, 
    -5.747283e-006, -2.861921e-006, -1.210625e-006, 3.220848e-007, 
    2.073965e-006, 5.455287e-006, -1.161823e-006, -3.689682e-006, 
    4.267051e-006, 1.366608e-005, 1.534184e-005, 1.929375e-005, 
    1.814834e-005, 1.255842e-005, 1.932902e-006, 9.169778e-006, 7.097022e-006,
  5.529051e-006, 4.772692e-006, 4.654472e-006, 8.841062e-007, 6.248276e-006, 
    8.944393e-006, 8.098878e-006, 7.279315e-006, 4.241462e-006, 
    3.140267e-006, 4.70227e-007, -3.407675e-006, -7.6781e-006, 
    -6.208349e-006, -7.192073e-006, -8.008412e-006, -3.47125e-006, 
    7.105082e-007, 2.457797e-006, 3.896006e-006, 5.854639e-006, 
    1.172346e-005, 1.231094e-005, 6.568909e-006, -3.679597e-007, 
    -8.504248e-006, -1.482903e-005, -9.502128e-006, -5.713628e-007, 
    1.057285e-005, -4.73239e-006, -4.776224e-006, -3.118341e-006, 
    1.996734e-006, 5.529051e-006, -1.448414e-006, -8.405696e-007, 
    8.363626e-006, 1.418812e-006, 5.478141e-006, 1.781556e-005, 7.43242e-006, 
    1.230201e-005, 2.49783e-005, 2.406685e-005, 1.165034e-005, 2.658606e-006, 
    1.478565e-005, 2.635394e-005, 4.765191e-005, 5.190258e-005, 
    4.813781e-005, 3.043348e-005, 2.797156e-005, 2.396266e-005, 
    2.070116e-005, 1.381769e-005, 8.686106e-006, 6.57486e-006, 3.525958e-006, 
    2.104141e-006, 5.257352e-007, -2.401844e-007, -7.824624e-007, 
    -5.482661e-007, -1.000765e-006, -1.880058e-006, -3.505775e-007, 
    -1.229628e-007, -9.943078e-007, -4.643243e-007, 1.184986e-006, 
    8.110901e-007, -1.964763e-007, 4.318572e-007, -3.981386e-007, 
    -4.180922e-006, -1.77227e-006, -3.401212e-006, -4.060346e-006, 
    -5.209473e-006, -3.332421e-006, -3.93232e-006, -5.146263e-006, 
    -6.883125e-006, -2.526469e-005, -2.305237e-005, 6.323287e-006, 
    3.598368e-005, 2.30789e-005, 6.987015e-006, 7.017799e-006, 1.537015e-005, 
    3.28332e-006, 3.007404e-006, 6.189919e-006,
  5.245187e-006, 7.454899e-006, 1.578999e-006, 4.78499e-006, 8.437633e-006, 
    1.097182e-005, 3.356708e-006, 8.042625e-006, 1.241587e-005, 
    4.697071e-006, 8.689085e-006, 3.001191e-006, -3.352292e-006, 
    -8.794196e-006, -8.784262e-006, -9.198517e-006, -3.229852e-006, 
    -1.244149e-006, 4.376925e-007, 2.320594e-007, 7.387102e-006, 
    1.151919e-005, 1.475051e-005, 8.611598e-006, 1.210257e-005, 
    1.672386e-006, -9.378018e-007, 4.615358e-007, -4.368776e-007, 
    1.063891e-005, -4.952801e-006, 1.016505e-005, 7.241317e-006, 
    6.645641e-006, 4.73953e-006, -1.045708e-006, -2.299392e-006, 
    9.360156e-007, 2.604203e-006, 3.486639e-007, -1.14913e-005, 
    -1.456951e-005, -1.772758e-006, 1.432882e-005, 1.688374e-005, 
    9.143827e-006, 2.835179e-006, -9.534037e-006, -1.032095e-005, 
    1.492946e-006, 1.078581e-005, 1.114716e-005, 1.277573e-005, 
    1.463602e-005, 1.240606e-005, 7.279312e-006, 7.304768e-006, 
    4.597849e-006, 3.719303e-006, 2.29798e-006, 2.105755e-006, 1.847096e-006, 
    9.653195e-007, -2.268976e-007, 4.969261e-007, 1.37982e-006, 
    2.857023e-007, -9.86247e-008, -1.079379e-007, -2.431401e-006, 
    6.37865e-007, -1.488652e-006, -2.719717e-007, -1.318404e-008, 
    -3.427165e-006, 9.133895e-006, 6.147711e-007, 1.049048e-007, 
    3.356254e-007, -2.848261e-006, -4.064568e-007, -7.874045e-006, 
    -2.350673e-005, -3.139988e-005, -3.862508e-005, -4.372238e-005, 
    -3.479796e-005, 9.326614e-006, 1.545087e-005, 1.737609e-005, 
    2.779168e-006, -1.225598e-005, -9.421281e-006, 1.391621e-006, 
    -3.324349e-006, 4.45878e-006,
  -2.505658e-006, -6.477203e-007, -1.150896e-006, -1.083056e-005, 
    1.373613e-006, 5.441252e-006, -6.124148e-006, -8.07162e-006, 
    -1.204164e-006, -5.614413e-006, 2.200378e-005, 8.375167e-006, 
    -5.415602e-007, -5.715618e-006, -7.10689e-006, -1.068254e-005, 
    -4.228234e-006, 1.142151e-006, 3.1569e-006, -3.89562e-007, 7.794653e-006, 
    5.14782e-006, 3.216635e-006, 5.825823e-006, 1.801636e-005, 5.443864e-006, 
    -3.765801e-006, 3.636727e-006, 4.255373e-006, 2.700312e-006, 
    -8.03826e-007, -3.105299e-006, 3.308029e-006, 7.241448e-006, 
    -1.002001e-006, -2.076005e-006, 1.479166e-006, 3.395828e-006, 
    4.467103e-006, -9.037758e-007, -1.992076e-005, -2.065973e-005, 
    -8.753705e-006, 7.034541e-007, 3.523615e-006, -2.441695e-006, 
    -1.523411e-006, -8.871546e-006, -1.045827e-005, -1.179839e-005, 
    -4.372276e-006, -3.713511e-006, -2.398883e-008, 2.563473e-006, 
    3.047266e-006, 4.643669e-006, 3.466361e-006, 2.355373e-007, 
    -3.710666e-007, 1.647666e-006, 3.623314e-006, 5.624539e-006, 
    6.979802e-006, 2.50113e-006, 9.996169e-006, 7.865427e-006, 1.23431e-005, 
    1.577795e-005, 1.449521e-005, 1.359505e-005, 1.284199e-006, 
    1.173303e-005, 2.825928e-005, 2.580792e-005, 5.018301e-006, 
    9.442971e-006, 2.59489e-006, -9.274954e-007, -1.310436e-005, 
    -6.84413e-006, -4.48888e-006, -9.314372e-006, -1.167322e-005, 
    -1.479924e-005, -1.550928e-005, -6.869217e-006, -1.992066e-006, 
    -2.42173e-007, -2.951929e-007, 2.901479e-006, 7.593728e-006, 
    -2.952809e-006, 1.730994e-006, 4.737922e-006, -1.237437e-006, 
    -2.622619e-008,
  -1.652169e-005, -1.903229e-005, -8.820269e-006, -3.847752e-006, 
    -3.952737e-007, 3.786852e-006, 3.114568e-006, -4.990543e-006, 
    -1.258095e-005, -1.323598e-005, -3.032779e-006, 1.798541e-006, 
    -5.352272e-007, -3.168636e-006, -6.53369e-006, -4.331425e-006, 
    6.239643e-007, 4.416928e-006, 1.342604e-005, 9.256204e-006, 
    1.251359e-005, 1.001045e-005, 2.480407e-005, 2.912541e-005, 
    1.525119e-005, 1.452612e-005, 1.142766e-006, 2.087625e-006, 7.75118e-006, 
    2.550158e-005, 2.012051e-005, 3.661567e-006, 6.170179e-006, 
    1.783519e-006, -4.433314e-007, -2.16566e-006, 8.801719e-006, 
    5.589274e-006, 1.137987e-005, 1.871199e-005, 7.954965e-006, 
    6.784612e-006, 2.151457e-006, 1.459989e-005, 1.370395e-005, 
    3.990506e-006, 4.253961e-007, 8.285933e-007, 3.855654e-006, 
    3.323432e-006, -2.39948e-006, -5.426773e-006, -2.943256e-006, 
    -2.687448e-006, 1.046159e-006, -3.75534e-007, 1.359087e-006, 
    1.077704e-006, 2.615128e-006, 5.119517e-006, -2.121451e-006, 
    -4.882884e-006, -2.450895e-006, 2.802262e-006, 9.2911e-006, 
    7.898205e-006, 9.56242e-006, 1.33539e-005, 2.238761e-005, 8.411444e-007, 
    1.420613e-005, 3.016005e-005, 5.320428e-006, -8.710354e-006, 
    -7.230046e-006, 5.544935e-006, -3.326211e-006, -1.179578e-005, 
    -6.160913e-006, -4.381715e-006, -8.470595e-006, -6.028543e-006, 
    -6.117079e-006, -6.353263e-006, -5.402692e-006, -2.731785e-006, 
    -2.628221e-006, -2.271958e-006, -1.361994e-006, -3.35056e-007, 
    3.66912e-007, -1.584023e-006, -3.482048e-006, -4.189111e-006, 
    -9.690866e-006, -8.273895e-006,
  -1.834858e-006, -1.40235e-006, -8.209536e-007, -2.836459e-007, 
    -5.88152e-006, -6.152843e-006, -3.940888e-006, -1.833243e-006, 
    4.016088e-006, -2.421093e-006, -2.458969e-006, -5.677616e-007, 
    -1.015045e-006, -5.388283e-007, -3.347079e-006, 2.278983e-006, 
    3.390112e-006, 7.474773e-006, 1.208444e-005, 1.333464e-005, 4.23898e-006, 
    1.498148e-005, 3.989808e-005, 3.76274e-005, 3.657327e-005, 2.341058e-005, 
    5.463735e-006, -3.368041e-008, 9.13538e-006, 1.490536e-005, 
    2.096988e-005, 2.375353e-006, 2.225213e-006, -3.379606e-006, 
    -4.632551e-006, -2.96846e-006, 6.028611e-006, 2.153054e-005, 
    2.293845e-005, 1.495851e-005, 9.593219e-006, 1.094115e-005, 
    1.974886e-005, 1.210927e-005, 3.531426e-006, 5.222584e-006, 
    1.104272e-006, 2.141889e-006, 2.493929e-006, 2.447738e-006, 
    -1.326105e-006, -3.361729e-006, 1.123521e-006, -1.635681e-006, 
    -1.525186e-007, 8.462321e-007, 6.51773e-007, -1.515105e-006, 
    -2.455119e-006, -3.278036e-006, -2.266619e-006, 6.625751e-007, 
    1.966552e-006, 3.468713e-006, 8.745095e-006, 5.789694e-006, 
    1.111184e-007, 1.073987e-005, 5.002541e-006, -6.484624e-006, 
    1.659665e-005, -7.497911e-006, -2.440105e-005, -8.281222e-006, 
    -8.706265e-007, -3.920028e-006, 1.617491e-006, 8.847273e-007, 
    -1.223787e-006, -1.781463e-006, -4.435485e-006, -1.473878e-006, 
    -1.034169e-006, -4.371295e-007, -3.894465e-007, -1.689198e-006, 
    -1.564154e-006, -1.583773e-006, -8.826728e-007, -3.302121e-007, 
    -1.649332e-007, -4.433368e-007, -5.969806e-006, -8.889936e-006, 
    -6.967563e-006, -1.645363e-006,
  -4.874077e-006, -3.705572e-006, -3.594934e-006, -3.555941e-006, 
    -2.962254e-006, -1.162566e-006, -1.129163e-006, -1.00747e-006, 
    -2.624117e-007, 6.782238e-007, -1.103334e-006, -5.877539e-007, 
    -7.099434e-007, 5.009002e-007, 2.961701e-006, 5.464975e-006, 
    -1.589982e-006, 7.492028e-006, 1.044122e-005, 2.029859e-005, 
    1.207078e-005, 2.098987e-005, 3.075821e-005, -2.290658e-005, 
    3.913898e-006, 2.351413e-005, 9.891592e-007, 4.118156e-006, 
    6.257465e-006, -3.074747e-006, -2.06046e-005, -2.423576e-005, 
    -2.261439e-005, -1.34934e-005, -1.083366e-005, 3.235393e-006, 
    1.402893e-005, 2.185215e-005, 1.909916e-005, 1.66288e-005, 
    -4.379603e-006, -5.777078e-006, 6.544069e-006, -2.406814e-007, 
    5.735419e-007, 1.793454e-006, 1.347285e-006, 6.479258e-007, 
    -1.715276e-006, -4.203521e-006, 1.530825e-007, -1.576076e-006, 
    -8.385923e-007, -2.011935e-006, -3.675401e-006, -1.442835e-006, 
    -8.542384e-007, -2.946734e-006, -4.30336e-006, -7.378213e-006, 
    -4.299013e-006, -2.781703e-006, -2.385952e-006, -9.3669e-007, 
    -2.359751e-006, -8.027037e-007, -2.90079e-006, 7.115526e-006, 
    8.51338e-006, -8.060524e-007, -6.409013e-006, -2.424124e-005, 
    -1.788539e-005, -1.396726e-005, -1.02529e-005, -2.58687e-006, 
    2.761777e-006, -4.82205e-007, -2.72272e-006, -2.383841e-006, 
    -1.362243e-006, 6.250748e-007, 1.971512e-008, -1.021379e-006, 
    -1.413777e-006, -1.259301e-006, -1.24291e-006, -2.105686e-006, 
    -1.307356e-006, -2.072775e-007, -2.087677e-007, -6.757909e-008, 
    -3.72954e-006, -1.329944e-005, -1.159909e-005, -5.598891e-006,
  -3.818824e-006, -1.613202e-006, -1.341753e-006, -1.33008e-006, 
    -6.692136e-007, -3.1171e-007, -3.129517e-007, -1.594698e-007, 
    -4.423412e-008, -2.256558e-007, -3.064202e-006, -6.862259e-007, 
    -2.684945e-008, 9.995922e-007, 3.076814e-006, 8.958676e-006, 
    6.506314e-006, 4.139016e-006, 1.039229e-005, 1.351594e-005, 
    9.090549e-006, 9.379137e-006, 1.722695e-005, 1.400619e-005, 
    1.395516e-005, 6.790317e-006, 5.919705e-006, 1.543223e-005, 
    9.209514e-006, -1.898185e-006, -8.755946e-006, -6.402683e-006, 
    -2.190597e-005, -2.838326e-005, -7.508723e-006, 6.88916e-006, 
    1.783704e-005, 5.024027e-006, 3.391608e-006, 5.831302e-006, 
    -6.838789e-006, -1.544433e-005, -8.496918e-006, -2.487777e-006, 
    1.417196e-006, 1.73568e-008, 7.973067e-007, 2.552788e-006, 2.292638e-006, 
    -6.666087e-007, -1.688828e-006, -3.495345e-006, -3.810381e-006, 
    -2.428297e-006, -1.419738e-006, -1.468197e-008, -1.776993e-006, 
    -1.945127e-006, -1.553102e-006, -3.914316e-006, -3.006586e-006, 
    -2.749913e-006, -1.830387e-006, -1.884652e-006, -2.089294e-006, 
    -1.622016e-007, -1.000765e-006, -3.661007e-007, -5.91181e-006, 
    -2.43027e-005, -7.438437e-006, -9.091478e-006, -9.216397e-006, 
    -1.663196e-005, -1.539901e-005, -2.82417e-006, -6.608752e-008, 
    -2.746065e-006, -1.771403e-006, 7.298695e-008, -1.340512e-006, 
    -6.195442e-007, -1.136118e-006, -3.420109e-007, -1.524418e-006, 
    -1.508647e-006, -1.841812e-006, -1.602772e-006, -2.186401e-006, 
    -1.050062e-006, -6.569203e-007, -2.831494e-007, -1.510136e-006, 
    -7.80389e-006, -1.001982e-005, -6.824885e-006,
  -3.460077e-006, -2.057629e-006, -3.192849e-006, -2.991684e-006, 
    -2.117855e-006, -1.457858e-006, -8.168594e-007, -5.164768e-007, 
    -2.455239e-007, -1.764819e-007, -1.640643e-007, -2.016897e-007, 
    -4.766162e-007, 3.202235e-007, 6.872887e-007, 4.701662e-006, 
    1.029258e-005, 6.417901e-006, 3.343297e-006, 2.6756e-006, 3.305297e-006, 
    1.099889e-005, 1.386128e-005, 1.688758e-005, 1.889776e-005, 
    1.532656e-005, 1.287855e-005, 5.255235e-006, -1.751163e-006, 
    1.159166e-006, -2.939032e-006, -5.659862e-006, -2.127785e-006, 
    -1.839017e-005, -9.157906e-006, 3.84323e-006, 4.761139e-006, 
    -5.373135e-006, -7.807612e-006, -4.410893e-006, -7.223112e-006, 
    -6.754475e-006, -5.359725e-007, 1.430235e-007, 3.122732e-007, 
    3.280456e-007, 3.216015e-006, 1.163382e-006, 2.911675e-007, 
    -2.214338e-007, -2.03528e-006, -3.107914e-006, -2.628221e-006, 
    -3.178322e-006, -1.461088e-006, 1.057581e-006, 9.397263e-008, 
    -2.75204e-007, 8.205188e-008, -1.070802e-006, -5.774482e-007, 
    3.81192e-007, -3.148148e-007, -6.113473e-007, 1.88224e-007, 
    7.668859e-007, 1.162018e-007, -1.441591e-006, 5.392703e-007, 
    2.910419e-006, 6.999551e-006, 1.986518e-007, -6.965816e-006, 
    -8.787487e-006, -5.7176e-006, -8.19876e-006, -4.13572e-006, 
    1.401426e-006, -7.440922e-007, -2.132011e-006, -1.621276e-006, 
    -1.003374e-006, -7.394992e-007, 4.982903e-007, -9.277501e-007, 
    -2.040506e-007, -3.462328e-007, -7.049775e-007, -8.469115e-007, 
    -1.554715e-006, -4.987191e-007, -4.429644e-007, -8.774572e-007, 
    -2.544028e-006, -3.862408e-006, -4.949448e-006,
  -2.588856e-006, -2.282389e-006, -3.753009e-006, -3.271205e-006, 
    -3.289583e-006, -2.782695e-006, -1.615437e-006, -1.063225e-006, 
    -7.206227e-007, -4.524018e-007, -3.303364e-007, -4.475588e-007, 
    -2.790516e-007, -3.492112e-007, 3.573788e-009, 6.36004e-007, 
    1.275388e-006, 1.178282e-006, 2.946553e-006, 3.156162e-006, 
    7.065481e-006, 1.313472e-005, 1.449222e-005, 1.789118e-005, 
    3.337696e-005, 4.388687e-005, 3.197749e-005, 1.287408e-007, 
    -6.330534e-006, 1.176295e-005, 6.139504e-006, 6.163715e-006, 
    4.683163e-006, -4.033398e-006, -9.473184e-006, 2.881898e-007, 
    5.476522e-006, 9.135132e-006, -7.072122e-007, -1.900171e-006, 
    -3.773501e-006, -2.543655e-006, -2.187007e-007, 2.014112e-006, 
    3.970854e-008, -1.536463e-006, 2.306751e-008, 7.672588e-007, 
    1.54398e-006, 2.856524e-006, 2.639712e-006, -1.261785e-006, 
    -6.014152e-007, -8.258021e-007, -2.0133e-006, -1.610844e-006, 
    2.407487e-007, -6.079972e-007, 1.066398e-006, 2.151683e-007, 
    -6.797691e-007, -7.438443e-007, -5.103921e-007, -1.537574e-007, 
    1.340704e-006, 1.935758e-006, 9.085711e-007, -1.626981e-007, 
    6.524071e-006, 9.653319e-006, 8.551007e-006, 1.162164e-005, 
    1.572917e-006, 7.101371e-007, -2.301014e-006, -7.320345e-006, 
    -1.13084e-005, -5.174083e-006, -1.918801e-006, -2.274443e-006, 
    -1.514235e-006, -2.534734e-007, -4.099338e-007, 2.413708e-007, 
    -5.491529e-009, -5.106413e-007, -4.548856e-007, -2.836478e-007, 
    2.989891e-007, -1.077506e-006, -1.316421e-006, -2.374527e-007, 
    -9.827588e-007, -9.579236e-007, -2.376638e-006, -3.110023e-006,
  -2.951451e-006, -4.045196e-006, -4.641739e-006, -3.112507e-006, 
    -2.849999e-006, -2.894826e-006, -2.738736e-006, -2.536081e-006, 
    -7.999713e-007, -4.265729e-007, -1.509391e-006, -9.686028e-007, 
    -5.170976e-007, -5.019481e-007, -5.904857e-007, -7.776157e-008, 
    4.25401e-007, 1.637612e-007, 1.341326e-006, 2.510446e-006, 2.829083e-006, 
    5.309752e-006, 5.154407e-006, 3.160509e-006, 5.208797e-006, 
    1.452625e-005, 2.409094e-005, 1.146892e-005, -1.275694e-006, 
    7.840223e-006, 7.688854e-006, 1.528112e-005, 1.536369e-005, 1.63314e-006, 
    -5.639489e-006, -6.77037e-006, -2.656649e-006, 7.685623e-006, 
    3.259975e-006, -3.72035e-006, 1.885201e-008, 1.44315e-006, 4.283311e-006, 
    5.643909e-006, 6.357302e-006, 2.602583e-006, -1.127425e-006, 
    -1.762338e-006, 2.042797e-006, 2.73421e-006, 4.269402e-006, 
    2.432461e-006, 1.337598e-006, -1.26689e-007, -2.0775e-006, 
    -2.297292e-006, -9.751866e-007, -8.284087e-007, 7.711069e-007, 
    2.335473e-007, -7.99972e-007, -4.854323e-007, -4.422195e-007, 
    3.803248e-007, 3.06444e-008, 8.523191e-007, 1.635003e-006, 1.526968e-006, 
    6.651973e-006, 1.176233e-005, 6.826567e-006, 8.502066e-007, 
    -1.552729e-006, 6.825685e-007, 2.316112e-006, -3.451059e-007, 
    -7.376475e-006, -7.670527e-006, -5.149743e-006, -2.835968e-006, 
    -3.692909e-006, -2.727935e-006, -1.548383e-006, 1.155804e-007, 
    -2.062848e-007, -5.290185e-007, -8.665311e-007, -1.826911e-007, 
    -4.535195e-008, -4.427166e-007, -1.569861e-007, -3.403945e-007, 
    1.005556e-007, -2.937041e-007, -1.243405e-006, -4.367806e-006,
  -4.918156e-006, -5.729275e-006, -6.361582e-006, -3.287969e-006, 
    -3.101705e-006, -3.4869e-006, -3.370174e-006, -2.624867e-006, 
    -3.328326e-006, -1.700622e-006, -4.126653e-007, -6.657366e-007, 
    -8.47779e-007, -2.695524e-006, -2.299897e-006, -1.26824e-006, 
    -3.001616e-007, 3.528819e-007, 1.131095e-006, 1.865722e-006, 
    1.989033e-007, 1.85206e-006, 3.238238e-007, -6.712016e-007, 
    -5.994261e-007, 5.67632e-006, 1.416973e-005, 1.952707e-005, 
    1.565066e-005, 1.081127e-005, 1.737958e-005, 2.103383e-005, 
    1.811147e-005, 9.577449e-006, 9.241798e-006, 1.375785e-005, 
    9.057636e-006, 6.465962e-006, 6.881957e-006, 8.486932e-006, 
    -9.637588e-007, -8.183739e-006, -6.461043e-006, 3.611422e-008, 
    4.91699e-006, 5.320806e-006, 2.769475e-006, 2.969649e-006, 2.030378e-006, 
    -9.006781e-007, -2.486412e-006, -7.729022e-007, 1.109838e-007, 
    2.269653e-007, 1.990256e-007, -1.902038e-006, -2.334668e-006, 
    -2.076008e-006, -1.184422e-006, -4.172607e-007, -5.27777e-007, 
    -8.060556e-007, -2.241654e-007, -2.566997e-007, -2.200647e-008, 
    -3.389046e-007, 1.593528e-006, 2.540497e-006, 1.229193e-006, 
    3.46325e-006, 6.864073e-006, 1.417695e-006, -3.7396e-006, 1.200136e-006, 
    3.988145e-006, 3.38117e-006, -2.23222e-006, -6.88573e-006, 
    -7.032628e-006, -9.030877e-006, -7.802648e-006, -3.699988e-006, 
    -1.677527e-006, 9.024734e-008, -1.127675e-006, -1.234962e-006, 
    3.39347e-007, 2.316856e-007, -4.117965e-007, 1.82139e-007, 
    -6.746777e-007, -1.249117e-006, -7.407389e-007, -6.688406e-007, 
    -2.175472e-006, -2.983985e-006,
  -4.3236e-006, -1.733654e-006, -2.661872e-006, -4.404936e-006, 
    -3.893205e-006, -4.625721e-006, -5.813965e-006, -3.846391e-006, 
    -6.864495e-006, -7.998598e-006, -3.793863e-006, -5.907717e-006, 
    -7.931544e-006, -4.6328e-006, -2.324857e-006, -2.041486e-006, 
    -1.977784e-006, 4.525957e-007, 1.40093e-006, -5.03187e-008, 
    -2.307348e-006, 1.020578e-006, 1.29389e-006, 1.496295e-006, 
    2.681561e-006, 2.813311e-006, 5.535134e-006, 6.847429e-006, 
    1.111959e-005, 1.509871e-005, 2.134241e-005, 1.956893e-005, 1.59616e-005, 
    1.299714e-005, 1.460286e-005, 8.320909e-006, 1.090253e-005, 
    1.476902e-005, 8.833882e-006, 4.670375e-006, 7.905161e-006, 
    6.951741e-006, 3.150577e-006, -4.369213e-009, -6.8386e-007, 
    -1.068147e-007, -1.39192e-006, -1.248991e-006, -4.239664e-007, 
    -2.396882e-007, 1.724531e-006, -8.911193e-007, -3.738482e-006, 
    -4.312174e-006, -2.283134e-006, -2.691551e-006, -1.073657e-006, 
    -2.492745e-006, -2.282018e-006, -6.304717e-007, -1.643378e-006, 
    -9.602836e-007, -1.038762e-006, -3.900652e-007, -6.782793e-007, 
    -2.606242e-006, 1.106137e-007, 1.797425e-006, -1.207023e-006, 
    1.644818e-006, 8.400129e-006, 4.179252e-006, 3.55496e-007, 
    -2.397373e-006, -4.076115e-006, -1.758737e-006, 1.419805e-006, 
    -4.056992e-006, -9.540494e-006, -1.273133e-005, -1.076003e-005, 
    -7.143022e-006, -7.165003e-006, -2.595685e-006, -1.347466e-006, 
    -1.911352e-006, -1.124446e-006, -5.207003e-007, -1.064966e-006, 
    -2.144305e-006, -2.585007e-006, -1.709316e-006, -1.612084e-006, 
    -1.96015e-006, -1.337904e-006, -2.663983e-006,
  -7.204613e-006, -7.082053e-007, -3.551968e-006, -4.996885e-006, 
    -2.698257e-006, -3.931696e-006, -3.77648e-006, 1.196784e-006, 
    3.44191e-007, -1.338647e-006, -3.689547e-007, -2.976289e-006, 
    -5.381335e-006, -5.10021e-007, -1.000765e-006, -1.49685e-006, 
    -1.238935e-006, 4.332242e-007, 8.610116e-007, 8.287257e-007, 
    1.78811e-006, 8.053785e-007, 4.164576e-007, 2.704407e-006, 1.659465e-006, 
    9.92266e-007, 2.457297e-006, 3.197389e-006, 3.786232e-006, 5.519485e-006, 
    6.748709e-006, 6.154156e-006, 5.625534e-006, 3.412337e-006, 
    3.440531e-006, 1.295626e-006, 4.443253e-006, 2.418063e-006, 
    5.061898e-006, 6.714065e-006, 9.160587e-006, 9.422602e-006, 
    6.169306e-006, 3.646168e-006, 3.809833e-006, 2.157783e-006, 
    -2.589331e-007, 6.204828e-007, 9.686737e-007, 2.53168e-006, 
    4.998939e-006, 4.486959e-006, 7.455274e-007, 1.18362e-006, 
    -3.081095e-007, -1.587498e-006, -3.691914e-006, -3.891342e-006, 
    -3.761828e-006, -1.276809e-006, -6.433866e-007, -3.294681e-007, 
    -3.643613e-007, -1.256568e-006, -1.613453e-006, -2.144679e-006, 
    -7.103172e-007, 7.871258e-007, 5.994087e-006, 6.471306e-006, 
    3.269288e-006, 8.166826e-007, 1.340337e-006, -2.515593e-006, 
    -4.615042e-006, -9.073847e-007, -1.430664e-006, -3.559544e-006, 
    -5.494705e-006, -5.308693e-006, -8.048395e-006, -7.297251e-006, 
    -6.368165e-006, -8.350515e-006, -4.369298e-006, -3.542407e-006, 
    -4.305346e-006, -5.824766e-006, -3.648205e-006, -4.097227e-006, 
    -6.43075e-006, -5.174458e-006, -3.522414e-006, -5.670168e-006, 
    -5.512466e-006, -1.060879e-005,
  -3.710542e-006, -3.710169e-006, -1.459621e-005, -6.806375e-006, 
    3.089106e-006, 2.764635e-006, 3.341338e-007, 1.25614e-006, 3.047007e-007, 
    -6.86352e-007, 2.664052e-006, 5.963042e-006, 2.641204e-006, 
    1.569684e-006, 1.250178e-006, 2.228191e-006, 2.73508e-006, 3.615863e-006, 
    2.966668e-006, 1.993872e-006, 2.440783e-006, 3.032357e-006, 
    3.180872e-006, 3.956353e-006, 2.40328e-006, 3.097054e-006, 4.931262e-006, 
    2.241477e-006, 2.93152e-007, 5.937836e-007, 3.011122e-006, 2.61401e-006, 
    6.592236e-007, 2.445751e-006, 2.40589e-006, 5.621434e-006, 5.075184e-006, 
    3.746136e-007, -1.924516e-006, -4.727663e-007, 4.347261e-006, 
    8.645631e-006, 7.751685e-006, 6.348739e-006, 5.143735e-006, 
    4.412454e-006, 9.18506e-007, 2.390367e-006, 4.817775e-007, 1.3073e-006, 
    2.690627e-006, 4.644664e-006, 9.442094e-006, 8.940669e-006, 
    6.354823e-006, 2.070612e-006, -1.326231e-006, -4.591944e-006, 
    -1.293696e-006, -5.120073e-007, -7.26337e-007, 1.015609e-006, 
    1.123146e-006, -1.408933e-006, -1.216213e-006, -1.159959e-006, 
    -2.284001e-006, -5.178677e-006, -9.596624e-007, 2.51181e-006, 
    4.652738e-006, 4.592137e-006, 2.959594e-006, -2.700865e-006, 
    -4.126783e-006, -2.651192e-006, -1.297791e-006, -4.211091e-006, 
    -3.142057e-006, -2.139339e-006, -1.20702e-006, 1.151089e-006, 
    -3.391542e-007, -4.976271e-006, -7.114835e-006, -2.120836e-006, 
    -1.486915e-006, -4.957292e-008, -1.887631e-006, -4.603617e-006, 
    -3.973917e-006, -3.590216e-006, -5.448763e-006, -3.336771e-006, 
    -3.886749e-006, -5.284724e-006,
  -2.571969e-006, -2.419854e-006, -1.541175e-006, 3.842735e-006, 
    4.408977e-006, 2.620094e-006, 2.521372e-006, 1.906823e-006, 
    1.650023e-007, -6.89206e-007, -1.174983e-006, 1.709135e-006, 
    1.853055e-006, 5.931615e-007, 1.30109e-006, 3.345408e-006, 1.36827e-006, 
    3.078048e-007, 2.558982e-007, 1.098188e-006, 1.585579e-006, 
    1.269551e-006, 1.214291e-006, 2.530933e-006, 4.447842e-006, 
    4.355084e-006, 3.45915e-006, 3.166469e-006, 1.056465e-006, -9.45256e-008, 
    2.268922e-006, 4.467962e-006, 5.442624e-006, 6.788199e-006, 5.72028e-006, 
    6.481481e-006, 7.275961e-006, 5.522345e-006, -9.152063e-007, 
    -1.5608e-006, 3.481133e-006, 8.39864e-006, 6.820856e-006, 3.49057e-006, 
    3.763385e-006, 4.761268e-006, 2.239742e-006, -4.402318e-007, 
    7.671224e-008, 3.335099e-007, 4.068983e-006, 3.36304e-006, 4.179748e-006, 
    7.742867e-006, 7.347488e-006, 2.701303e-006, 2.784254e-006, 
    -3.890709e-007, 1.348153e-006, 1.451594e-006, 1.307671e-006, 
    6.995797e-007, 1.799035e-007, 5.659695e-007, -1.707576e-006, 
    -4.163787e-006, 1.281473e-006, -1.610844e-006, -4.323723e-006, 
    1.079685e-006, 4.44561e-006, 3.545952e-006, 3.267058e-006, 3.675723e-006, 
    5.540474e-006, 3.43407e-006, 2.616616e-006, 1.762659e-006, 
    -1.657405e-006, -8.425763e-006, -3.775236e-006, -1.416633e-006, 
    2.731853e-006, 5.095673e-006, 3.036454e-006, 1.662072e-006, 
    1.300843e-006, 2.921097e-006, 3.32355e-006, 2.376459e-006, 
    -1.754017e-006, -4.054758e-006, -3.040235e-006, -1.719251e-006, 
    -2.068185e-006, -1.379381e-006,
  -2.11537e-006, 1.349891e-006, 9.755004e-007, 1.655242e-006, 1.463764e-006, 
    9.022388e-007, 1.021572e-006, 1.797671e-006, 8.616298e-007, 
    2.171069e-006, 4.725862e-007, -8.343686e-007, 8.882071e-007, 
    8.683364e-007, 1.844983e-006, 3.07048e-006, 1.362432e-006, 
    -1.424578e-007, -5.149868e-007, 2.342682e-006, 2.882478e-006, 
    2.049253e-006, 3.837269e-006, 5.093811e-006, 5.794534e-006, 
    5.448457e-006, 6.45056e-006, 7.38213e-006, 6.001292e-006, 6.7152e-007, 
    -1.634808e-006, -1.795121e-006, 3.26519e-006, 1.017833e-005, 
    7.966137e-006, 6.876238e-006, 6.656319e-006, 4.104619e-006, 
    3.951014e-006, 4.513657e-006, 6.780743e-006, 8.542309e-006, 
    3.253142e-006, 2.285562e-006, 4.55774e-006, 8.452778e-006, 7.987364e-006, 
    6.522954e-006, 4.463862e-006, 2.885829e-006, 1.82375e-006, 2.79965e-006, 
    4.313733e-006, 5.677935e-006, 4.723517e-006, 3.5462e-006, 2.201867e-006, 
    1.053235e-006, 2.225212e-006, 2.952884e-006, 2.216644e-006, 
    1.214416e-006, 3.095447e-007, 4.299083e-006, 3.940582e-006, 
    1.673001e-006, 9.44332e-007, 1.871307e-006, 6.83675e-006, 7.381635e-006, 
    8.394292e-006, 7.370711e-006, 7.560328e-006, 4.325653e-006, 
    1.667659e-006, 3.597113e-006, 6.505819e-006, 6.078033e-006, 6.15192e-006, 
    1.49816e-006, 2.468227e-006, 1.497168e-006, 5.083009e-006, 7.542816e-006, 
    6.710712e-006, 5.933864e-006, 3.166966e-006, 2.062663e-006, 
    4.559977e-006, 3.952506e-006, 2.483375e-006, 2.106497e-006, 
    1.475311e-006, 1.609047e-006, -2.177076e-007, -9.135929e-007,
  -2.333563e-007, 1.474192e-006, 4.284428e-006, 4.509062e-006, -6.02533e-007, 
    -9.587948e-007, -6.509608e-007, 3.220732e-006, 3.740164e-006, 
    3.169076e-006, 1.47233e-006, 2.200499e-006, 4.393205e-006, 3.564081e-006, 
    3.050485e-006, 1.808727e-006, 2.531056e-006, 3.145233e-006, 
    7.951976e-007, 5.746606e-007, 1.248067e-006, 1.844364e-006, 
    2.788973e-006, 4.614861e-006, 4.74388e-006, 4.236246e-006, 6.878099e-006, 
    6.33433e-006, 5.723632e-006, 4.894257e-006, 1.286066e-006, 3.895129e-007, 
    4.192289e-006, 7.556349e-006, 8.336798e-006, 9.253346e-006, 
    4.071093e-006, 4.793179e-006, 4.857129e-006, 5.96565e-006, 9.010206e-006, 
    8.161584e-006, 6.085108e-006, 6.804587e-006, 6.732067e-006, 5.97695e-006, 
    6.665509e-006, 6.456147e-006, 4.172295e-006, 1.964816e-006, 
    1.160895e-006, 1.179769e-006, 2.255882e-006, 2.873785e-006, 3.3577e-006, 
    2.261595e-006, 2.422403e-007, 1.310529e-006, 2.176408e-006, 
    5.227052e-006, 7.771923e-006, 8.13017e-006, 7.694805e-006, 6.070335e-006, 
    5.779013e-006, 3.471197e-006, 4.279213e-006, 7.779743e-006, 
    1.066436e-005, 1.081511e-005, 6.691338e-006, 6.998052e-006, 
    9.592595e-006, 6.669234e-006, 4.695452e-006, 3.168703e-006, 
    2.717941e-006, 2.611152e-006, 5.728351e-006, 7.750934e-006, 
    4.691105e-006, 4.2057e-006, 5.571763e-006, 7.505934e-006, 4.380043e-006, 
    4.085372e-006, 4.249658e-006, 5.346135e-006, 3.365647e-006, 
    3.074329e-006, 2.747993e-006, 2.034973e-006, 8.165553e-007, 
    2.209812e-006, 3.312498e-006, 6.238333e-007,
  1.915267e-006, 3.359562e-006, 3.869305e-006, 8.990213e-006, 9.189516e-006, 
    3.77518e-006, 1.388636e-006, 8.22889e-007, 2.180135e-006, 3.24234e-006, 
    4.222091e-006, 5.994709e-006, 5.775537e-006, 4.479507e-006, 
    2.926063e-006, 1.028402e-006, 7.557082e-007, 1.344182e-006, 
    1.712735e-006, 2.554529e-006, 1.931287e-006, 2.084147e-006, 
    1.956865e-006, 5.50197e-007, 6.898954e-007, 1.509832e-006, 1.616747e-006, 
    1.811582e-006, 2.048884e-006, 3.97262e-006, 4.939207e-006, 1.175673e-006, 
    8.329453e-007, 2.865961e-006, 3.76835e-006, 4.131318e-006, 3.716197e-006, 
    3.428231e-006, 4.914746e-006, 7.124838e-006, 8.250123e-006, 
    5.168315e-006, 3.575628e-006, 2.311389e-006, 2.996101e-006, 
    2.521497e-006, 4.13852e-006, 3.766115e-006, 5.266029e-007, -1.75366e-007, 
    3.033338e-007, 2.145862e-006, 2.673365e-006, 3.544708e-006, 
    4.508938e-006, 6.108083e-006, 7.529283e-006, 7.067221e-006, 
    3.880112e-006, 4.257607e-006, 6.148563e-006, 5.742382e-006, 
    3.602701e-006, 2.115812e-006, 4.471933e-006, 2.293384e-006, 
    1.629537e-006, 4.561093e-006, 7.425468e-006, 9.560556e-006, 
    4.805967e-006, 2.841499e-006, 3.193414e-006, 4.34341e-006, 3.040304e-006, 
    2.507712e-006, 4.260463e-006, 5.850542e-006, 6.859597e-006, 
    7.977929e-006, 8.062369e-006, 7.172148e-006, 6.184821e-006, 6.24691e-006, 
    7.3265e-006, 5.614607e-006, 2.950774e-006, 3.950516e-006, 1.682312e-006, 
    4.383128e-007, 1.137178e-006, 1.696841e-006, 1.616996e-006, 
    1.075214e-006, 1.399314e-006, 5.424972e-007,
  2.729863e-006, 1.754831e-006, 5.521824e-007, 1.949911e-006, 5.518741e-006, 
    6.38251e-006, 6.395674e-006, 4.530173e-006, 1.230683e-006, 2.528946e-006, 
    9.75253e-007, 3.841742e-006, 6.866426e-006, 3.436055e-006, 1.22112e-006, 
    -5.998008e-007, -1.459357e-007, -9.216819e-008, 1.393355e-006, 
    1.626184e-006, 4.486201e-007, -4.701615e-007, -5.508755e-007, 
    4.533395e-007, 8.051302e-007, 1.270916e-006, -7.365197e-007, 
    -2.414017e-006, 3.262903e-008, 8.61507e-007, 2.44016e-006, 2.356092e-006, 
    2.421038e-006, 2.591409e-006, 3.836027e-006, 5.247538e-006, 
    4.690608e-006, 4.376443e-006, 3.439531e-006, 2.54211e-006, 2.847086e-006, 
    1.894902e-006, 1.002199e-006, 1.926691e-006, 3.229053e-006, 
    3.664788e-006, 3.541977e-006, 2.212918e-006, 1.222735e-006, 6.39976e-007, 
    1.579228e-007, 6.607133e-007, 2.562711e-007, 3.485338e-007, 
    1.496048e-006, 3.515526e-006, 4.056688e-006, 2.756189e-006, 
    1.350763e-006, 4.590771e-006, 7.908266e-006, 8.591112e-006, 
    7.670592e-006, 4.480874e-006, 2.513672e-006, 2.401914e-006, 
    3.220734e-006, 5.131186e-006, 6.1806e-006, 5.448207e-006, 4.721031e-006, 
    4.512292e-006, 4.066125e-006, 4.052714e-006, 3.12996e-006, 3.344909e-006, 
    3.827955e-006, 3.133188e-006, 6.484211e-006, 1.05485e-005, 7.925153e-006, 
    4.496894e-006, 2.816167e-006, 1.921104e-006, 3.346398e-006, 
    5.140622e-006, 3.90718e-006, 2.043294e-006, 7.228045e-007, 3.546193e-007, 
    9.586129e-007, 2.094826e-006, 7.548388e-007, -2.740853e-007, 
    4.278827e-007, 9.684227e-007,
  1.076209e-006, 8.818706e-007, 9.100595e-007, -1.196104e-007, 
    -8.782026e-007, -7.974995e-008, 1.627922e-006, 1.554286e-006, 
    2.352121e-006, 2.866085e-006, 3.451949e-006, 2.609288e-006, 
    1.483878e-006, 1.551679e-006, 2.70478e-006, 2.274261e-006, 8.463567e-007, 
    1.545718e-006, 9.937539e-007, -6.587852e-007, -1.090298e-006, 
    -1.033177e-006, -4.299272e-007, -2.872493e-007, 3.942305e-007, 
    1.954231e-007, -1.240673e-006, 4.277572e-007, 1.561364e-006, 
    7.283898e-007, 8.785191e-007, 1.209572e-006, 1.469723e-006, 1.75036e-006, 
    2.261223e-006, 1.589056e-006, 1.83269e-006, 1.137427e-006, 2.017339e-006, 
    3.571407e-006, 2.860746e-006, 1.857527e-006, 1.853801e-006, 
    2.457795e-006, 2.21056e-006, 1.8389e-006, 2.386021e-006, 1.392362e-006, 
    1.368767e-006, 2.231047e-006, 1.828469e-006, 1.044419e-006, 
    9.959904e-007, 1.293019e-006, 1.702429e-006, 1.656111e-006, 
    7.965618e-007, 1.033864e-006, 9.932573e-007, 1.579618e-006, 
    2.632137e-006, 3.390109e-006, 3.238241e-006, 3.349752e-006, 
    4.300942e-006, 4.692472e-006, 3.883462e-006, 2.594884e-006, 
    2.479774e-006, 3.118538e-006, 3.713466e-006, 4.086118e-006, 
    3.594007e-006, 3.744509e-006, 2.969526e-006, 2.775811e-006, 
    2.259238e-006, 3.287788e-006, 5.969376e-006, 7.659913e-006, 5.54457e-006, 
    3.894888e-006, 3.751091e-006, 2.789717e-006, 1.355852e-006, 
    7.856379e-007, 1.112718e-006, -1.146301e-006, -1.277183e-006, 
    9.673049e-007, 2.778665e-006, 2.622329e-006, 3.218249e-006, 
    1.906823e-006, 8.940415e-007, 6.150167e-007,
  -4.310436e-007, -5.195811e-007, -2.179577e-007, -1.310345e-007, 
    -9.241558e-008, 8.105944e-007, 1.558135e-006, 1.816795e-006, 
    9.969835e-007, 5.437396e-007, 8.319539e-007, 4.407984e-007, 
    6.261935e-007, 1.853924e-006, 1.887203e-006, 1.713232e-006, 
    1.614388e-006, 7.225544e-007, -6.596565e-008, 3.620698e-007, 
    9.538944e-007, 1.234534e-006, 1.244965e-006, 7.143581e-007, 
    6.251994e-007, 1.291281e-006, 1.702429e-006, 1.020452e-006, 
    -2.821707e-008, 3.852892e-007, 1.01176e-006, 7.662643e-007, 
    1.054602e-006, 1.390995e-006, 9.250866e-007, 1.307425e-006, 
    1.080183e-006, 9.928867e-007, 1.301092e-006, 8.603906e-007, 
    5.966403e-007, 8.458624e-007, 1.194797e-006, 1.675111e-006, 
    1.783145e-006, 2.161138e-006, 2.670385e-006, 2.482009e-006, 
    1.743284e-006, 6.417158e-007, 2.289535e-007, -2.108786e-007, 
    -1.239555e-007, 9.347741e-008, 3.761029e-007, 7.349727e-007, 
    5.509432e-007, -1.459343e-007, -3.513219e-007, 6.951177e-008, 
    8.255029e-008, 5.013999e-008, 3.051982e-007, 1.974131e-007, 
    3.911282e-007, 1.604455e-006, 1.694732e-006, 8.731809e-007, 
    3.120281e-007, 3.096688e-007, 1.694732e-006, 2.818031e-006, 
    3.448101e-006, 3.034098e-006, 2.575141e-006, 2.372983e-006, 
    2.171442e-006, 3.466602e-006, 4.085125e-006, 3.308155e-006, 
    2.466984e-006, 2.007904e-006, 1.658969e-006, 1.565961e-006, 
    1.848586e-006, 1.141029e-006, 1.321954e-006, 1.625689e-006, 
    1.033243e-006, 1.374604e-006, 2.043542e-006, 2.766994e-006, 
    2.824736e-006, 2.093459e-006, 5.991214e-007, -3.628793e-008,
  5.46097e-008, -2.394399e-007, -2.586871e-007, -1.081844e-007, 
    3.547448e-007, 1.397205e-006, 1.917131e-006, 1.757813e-006, 
    1.501513e-006, 8.031448e-007, 3.076811e-007, 1.632643e-007, 
    -1.341377e-007, -4.124172e-007, -5.010788e-007, -5.265356e-007, 
    -1.290468e-007, 5.134416e-007, 1.314379e-006, 1.7937e-006, 1.889067e-006, 
    1.328411e-006, 8.359279e-007, 1.021695e-006, 1.387767e-006, 
    1.239128e-006, 1.061928e-006, 1.141277e-006, 5.565307e-007, 
    -1.959779e-007, -8.780785e-007, -5.58573e-007, 3.881478e-007, 
    4.594244e-007, -6.758e-008, -3.559171e-007, -1.959779e-007, 
    1.767999e-007, 4.856265e-007, 8.235102e-007, 8.05132e-007, 5.469697e-007, 
    2.989896e-007, 3.076821e-008, 3.259356e-007, 7.076537e-007, 
    8.302159e-007, 8.432544e-007, 7.230515e-007, 8.949119e-007, 1.10328e-006, 
    1.087261e-006, 1.085647e-006, 1.061556e-006, 9.480591e-007, 
    1.013997e-006, 1.243971e-006, 1.377213e-006, 1.37237e-006, 9.080741e-007, 
    4.826466e-007, -2.31616e-007, -7.782405e-007, -9.251407e-007, 
    -1.005607e-006, -9.140895e-007, -5.396973e-007, 1.314756e-007, 
    3.444384e-007, 5.585207e-008, 3.672862e-007, 1.878516e-007, 
    -1.173739e-007, 2.551551e-007, 4.511053e-007, 5.725501e-007, 
    8.448687e-007, 1.423779e-006, 1.969161e-006, 2.417438e-006, 2.28966e-006, 
    1.82698e-006, 1.315125e-006, 7.629121e-007, 6.268153e-007, 1.11458e-006, 
    1.466495e-006, 1.67002e-006, 1.38665e-006, 1.11371e-006, 1.032375e-006, 
    1.02331e-006, 5.719294e-007, -7.490598e-008, 1.975359e-007, 2.403776e-007,
  5.011484e-007, 9.222304e-007, 1.326548e-006, 1.484501e-006, 1.405152e-006, 
    1.343809e-006, 1.160152e-006, 1.027656e-006, 1.16723e-006, 1.17704e-006, 
    1.046904e-006, 7.897343e-007, 3.48411e-007, 2.654615e-007, 6.135278e-007, 
    9.009959e-007, 8.226407e-007, 8.317056e-007, 1.106136e-006, 
    1.471587e-006, 1.566953e-006, 1.549693e-006, 1.517035e-006, 
    1.314751e-006, 1.026787e-006, 7.1349e-007, 3.356217e-007, -4.833146e-008, 
    -2.865022e-007, -9.005498e-008, 2.326797e-007, 2.729125e-007, 
    1.596632e-007, 2.479524e-007, 4.553272e-007, 5.256115e-007, 
    4.970507e-007, 4.650133e-007, 2.673246e-007, -6.037681e-008, 
    5.771426e-008, 8.967741e-007, 1.468606e-006, 1.325679e-006, 
    1.077824e-006, 9.810901e-007, 8.791412e-007, 8.29843e-007, 9.414775e-007, 
    1.104894e-006, 1.193183e-006, 1.26682e-006, 1.070497e-006, 7.211893e-007, 
    4.602944e-007, 3.890173e-007, 3.299097e-007, 3.525097e-007, 
    5.901829e-007, 8.574102e-007, 9.80966e-007, 7.744607e-007, 3.3885e-007, 
    3.710147e-008, 4.716003e-008, 2.083407e-007, 4.593012e-007, 
    7.565791e-007, 8.097268e-007, 5.737916e-007, 3.073092e-007, 
    1.990275e-007, 2.254774e-007, 5.937841e-007, 1.088254e-006, 
    1.302334e-006, 1.215535e-006, 1.03908e-006, 1.232671e-006, 1.857154e-006, 
    2.663679e-006, 3.04875e-006, 2.636485e-006, 1.731736e-006, 8.18171e-007, 
    3.513917e-007, 3.869063e-007, 5.85216e-007, 7.334825e-007, 7.542199e-007, 
    6.343896e-007, 4.21303e-007, 9.72027e-008, -3.511977e-007, 
    -5.334891e-007, -1.294193e-007,
  7.807921e-008, 1.442659e-007, 2.970028e-007, 4.816525e-007, 6.470555e-007, 
    7.829049e-007, 9.430923e-007, 1.184243e-006, 1.471214e-006, 
    1.746141e-006, 1.921229e-006, 1.948548e-006, 1.893662e-006, 
    1.830705e-006, 1.793328e-006, 1.822757e-006, 1.871932e-006, 
    1.791341e-006, 1.473697e-006, 9.864298e-007, 5.949018e-007, 4.76934e-007, 
    5.988754e-007, 8.490906e-007, 1.034734e-006, 1.059197e-006, 
    9.091918e-007, 6.213513e-007, 3.038322e-007, 9.260839e-008, 
    3.300374e-008, 1.333378e-007, 3.192299e-007, 5.530542e-007, 
    6.843088e-007, 5.554134e-007, 1.991516e-007, -2.139836e-007, 
    -4.884132e-007, -5.475208e-007, -4.419717e-007, -2.285119e-007, 
    3.747436e-008, 1.894659e-007, 2.782517e-007, 3.741161e-007, 4.04043e-007, 
    4.514777e-007, 5.582697e-007, 6.564933e-007, 6.812043e-007, 
    6.603423e-007, 6.17129e-007, 5.797524e-007, 6.408468e-007, 7.759509e-007, 
    9.124205e-007, 1.031009e-006, 1.082046e-006, 1.015984e-006, 
    8.787688e-007, 7.159738e-007, 5.616225e-007, 4.734575e-007, 
    4.857507e-007, 4.961817e-007, 4.504845e-007, 3.356213e-007, 
    2.395091e-007, 1.748131e-007, 1.112348e-007, -1.703938e-008, 
    -1.667963e-007, -1.797102e-007, 1.810258e-008, 3.114073e-007, 
    5.243696e-007, 6.68414e-007, 7.925905e-007, 9.366347e-007, 1.071863e-006, 
    1.157172e-006, 1.197405e-006, 1.166113e-006, 1.002573e-006, 
    7.836495e-007, 5.647269e-007, 3.36739e-007, 1.643823e-007, 6.702817e-008, 
    8.677216e-008, 1.724538e-007, 2.429861e-007, 2.573906e-007, 
    2.170332e-007, 1.315993e-007,
  9.243413e-007, 1.026291e-006, 1.134076e-006, 1.241488e-006, 1.333254e-006, 
    1.40242e-006, 1.440543e-006, 1.447869e-006, 1.436445e-006, 1.414962e-006, 
    1.381807e-006, 1.33015e-006, 1.264585e-006, 1.195294e-006, 1.123148e-006, 
    1.056093e-006, 1.000834e-006, 9.555097e-007, 9.176356e-007, 
    8.813768e-007, 8.493389e-007, 8.170532e-007, 7.850158e-007, 
    7.585659e-007, 7.344756e-007, 7.116273e-007, 6.769824e-007, 
    6.342657e-007, 5.797519e-007, 5.186571e-007, 4.540857e-007, 
    3.859132e-007, 3.146356e-007, 2.412476e-007, 1.759308e-007, 
    1.221624e-007, 8.292272e-008, 5.063703e-008, 1.785429e-008, 
    -1.592161e-008, -5.143602e-008, -8.322513e-008, -1.039625e-007, 
    -1.155108e-007, -1.136486e-007, -9.713267e-008, -6.074924e-008, 
    -1.008539e-008, 5.932907e-008, 1.484877e-007, 2.509332e-007, 
    3.621949e-007, 4.69111e-007, 5.731708e-007, 6.704008e-007, 7.545923e-007, 
    8.223924e-007, 8.740499e-007, 9.07205e-007, 9.09813e-007, 8.752918e-007, 
    8.083607e-007, 7.231761e-007, 6.321548e-007, 5.463489e-007, 
    4.739541e-007, 4.334725e-007, 4.218e-007, 4.232902e-007, 4.334725e-007, 
    4.563212e-007, 4.893518e-007, 5.328134e-007, 5.718048e-007, 
    5.983788e-007, 6.115415e-007, 6.09803e-007, 5.978818e-007, 5.778893e-007, 
    5.603811e-007, 5.494535e-007, 5.401398e-007, 5.310749e-007, 
    5.225065e-007, 5.126972e-007, 5.000306e-007, 4.923322e-007, 
    4.883586e-007, 4.903454e-007, 5.05991e-007, 5.456036e-007, 6.116657e-007, 
    6.812043e-007, 7.403119e-007, 7.898584e-007, 8.479728e-007,
  -3.141645e-008, -3.141668e-008, -3.091986e-008, -3.166497e-008, 
    -3.30308e-008, -3.576281e-008, -3.390016e-008, -2.967806e-008, 
    -2.073739e-008, -5.712081e-009, 1.452861e-008, 3.663195e-008, 
    5.997708e-008, 8.481254e-008, 1.082818e-007, 1.277774e-007, 
    1.395742e-007, 1.4926e-007, 1.492599e-007, 1.470247e-007, 1.403193e-007, 
    1.301369e-007, 1.189609e-007, 1.030663e-007, 8.828931e-008, 7.50025e-008, 
    6.780022e-008, 6.668267e-008, 7.47541e-008, 9.189046e-008, 1.233071e-007, 
    1.646579e-007, 2.150733e-007, 2.678483e-007, 3.204991e-007, 3.65451e-007, 
    4.044424e-007, 4.364798e-007, 4.631778e-007, 4.840393e-007, 
    5.008033e-007, 5.127241e-007, 5.201747e-007, 5.296121e-007, 
    5.424023e-007, 5.627672e-007, 5.898376e-007, 6.183983e-007, 
    6.475797e-007, 6.840874e-007, 7.268042e-007, 7.737428e-007, 
    8.250274e-007, 8.698553e-007, 9.104608e-007, 9.401392e-007, 
    9.510666e-007, 9.385249e-007, 9.05618e-007, 8.537124e-007, 7.891408e-007, 
    7.087988e-007, 6.179014e-007, 5.180636e-007, 4.123895e-007, 
    3.046046e-007, 1.978128e-007, 1.040596e-007, 2.595289e-008, 
    -3.948799e-008, -9.449832e-008, -1.333653e-007, -1.631679e-007, 
    -1.821668e-007, -1.9148e-007, -1.934668e-007, -1.924734e-007, 
    -1.84526e-007, -1.739711e-007, -1.616777e-007, -1.513711e-007, 
    -1.425544e-007, -1.312544e-007, -1.123797e-007, -9.15179e-008, 
    -6.904202e-008, -4.457911e-008, -2.582874e-008, -1.365947e-008, 
    -6.581558e-009, -3.849664e-009, -4.842832e-009, -1.055491e-008, 
    -1.589456e-008, -2.371758e-008, -2.992647e-008,
  4.965812e-007, 4.839152e-007, 4.670271e-007, 4.526228e-007, 4.34493e-007, 
    4.152457e-007, 4.102786e-007, 3.968676e-007, 3.742675e-007, 
    3.424783e-007, 3.082056e-007, 2.826253e-007, 2.623846e-007, 
    2.401571e-007, 2.22524e-007, 2.053877e-007, 1.907349e-007, 1.789381e-007, 
    1.733501e-007, 1.666447e-007, 1.557171e-007, 1.454105e-007, 
    1.358489e-007, 1.254181e-007, 1.257906e-007, 1.262873e-007, 1.35228e-007, 
    1.524885e-007, 1.829118e-007, 2.12714e-007, 2.397846e-007, 2.523263e-007, 
    2.59156e-007, 2.704561e-007, 2.941738e-007, 3.319234e-007, 3.740191e-007, 
    4.123896e-007, 4.291534e-007, 4.281601e-007, 4.378458e-007, 
    4.444272e-007, 4.736086e-007, 5.381802e-007, 6.73905e-007, 8.56941e-007, 
    1.036748e-006, 1.212209e-006, 1.390775e-006, 1.590451e-006, 1.78131e-006, 
    1.961614e-006, 2.16191e-006, 2.3745e-006, 2.589077e-006, 2.783413e-006, 
    2.859657e-006, 2.803902e-006, 2.643342e-006, 2.444039e-006, 
    2.222508e-006, 1.99539e-006, 1.817693e-006, 1.636893e-006, 1.459196e-006, 
    1.287584e-006, 1.119822e-006, 9.934106e-007, 9.092191e-007, 
    8.283803e-007, 7.439405e-007, 6.290775e-007, 4.112719e-007, 1.56338e-007, 
    -2.545607e-008, -1.203268e-007, -1.531096e-007, -1.738467e-007, 
    -1.698736e-007, -1.428025e-007, -1.013277e-007, -4.557296e-008, 
    6.581331e-008, 1.899898e-007, 2.904485e-007, 3.298123e-007, 
    3.228583e-007, 2.832462e-007, 2.558031e-007, 2.919387e-007, 
    3.886721e-007, 4.978231e-007, 5.621462e-007, 5.553165e-007, 
    5.184361e-007, 4.981955e-007,
  2.659857e-007, 3.499289e-007, 3.935148e-007, 3.845742e-007, 3.213685e-007, 
    2.181779e-007, 1.918525e-007, 2.052635e-007, 2.096097e-007, 
    1.976887e-007, 1.917282e-007, 1.873821e-007, 1.844019e-007, 
    2.086163e-007, 2.571692e-007, 3.007551e-007, 3.272046e-007, 
    3.212442e-007, 2.764165e-007, 2.30223e-007, 2.084921e-007, 1.947084e-007, 
    1.702457e-007, 1.642853e-007, 1.606842e-007, 1.835326e-007, 2.43634e-007, 
    3.085782e-007, 3.50674e-007, 3.618499e-007, 3.173948e-007, 2.867232e-007, 
    2.966572e-007, 3.439684e-007, 3.658235e-007, 3.231068e-007, 
    2.777825e-007, 2.975265e-007, 3.736466e-007, 5.06267e-007, 6.843358e-007, 
    8.81652e-007, 1.099706e-006, 1.340856e-006, 1.703327e-006, 2.247716e-006, 
    2.66557e-006, 2.879029e-006, 2.897034e-006, 2.957259e-006, 3.017486e-006, 
    3.01823e-006, 2.922491e-006, 2.895668e-006, 3.113101e-006, 3.308679e-006, 
    3.472095e-006, 3.691018e-006, 3.814946e-006, 3.57243e-006, 2.95577e-006, 
    2.298131e-006, 1.89431e-006, 1.718601e-006, 1.486887e-006, 1.114483e-006, 
    6.837149e-007, 2.620122e-007, 1.477702e-008, -1.87506e-008, 
    -2.409024e-008, -6.022583e-008, -1.192093e-007, -1.610565e-007, 
    -1.821668e-007, -2.33576e-007, -2.024076e-007, -1.493841e-007, 
    -2.165634e-007, -3.543992e-007, -4.212061e-007, -4.420676e-007, 
    -2.546853e-007, 8.30737e-008, 3.679347e-007, 5.291154e-007, 
    6.288287e-007, 6.477039e-007, 6.400051e-007, 5.047768e-007, 
    3.361456e-007, 2.833708e-007, 3.213684e-007, 3.180155e-007, 2.84612e-007, 
    2.529471e-007,
  2.371768e-007, 3.209958e-007, 3.429751e-007, 3.68307e-007, 3.894171e-007, 
    4.178535e-007, 5.03535e-007, 5.969157e-007, 5.638848e-007, 4.786998e-007, 
    4.995615e-007, 5.754332e-007, 5.397947e-007, 3.955016e-007, 
    2.983958e-007, 1.973162e-007, 1.670172e-007, 1.991789e-007, 
    2.189229e-007, 2.517054e-007, 3.160287e-007, 3.187607e-007, 3.30309e-007, 
    3.00631e-007, 2.684693e-007, 2.056361e-007, 1.470248e-007, 2.284845e-007, 
    4.046907e-007, 4.763405e-007, 3.97116e-007, 3.073364e-007, 1.621743e-007, 
    1.465276e-008, 1.175951e-007, 3.491839e-007, 6.51305e-007, 8.856256e-007, 
    9.300808e-007, 8.640189e-007, 8.70352e-007, 1.128639e-006, 1.494338e-006, 
    1.79174e-006, 2.025316e-006, 2.52674e-006, 3.270432e-006, 3.742675e-006, 
    3.715232e-006, 3.229951e-006, 2.81396e-006, 2.779314e-006, 2.92485e-006, 
    3.134708e-006, 3.411124e-006, 3.833075e-006, 4.197657e-006, 
    4.234663e-006, 3.891066e-006, 3.46986e-006, 3.214305e-006, 2.970547e-006, 
    2.70456e-006, 2.193698e-006, 1.696001e-006, 1.515945e-006, 1.139442e-006, 
    9.205196e-007, 1.684451e-006, 2.409269e-006, 2.131114e-006, 
    1.234809e-006, 4.683934e-007, -2.513325e-007, -8.111192e-007, 
    -5.359443e-007, 3.453342e-007, 7.321441e-007, 7.374838e-007, 
    1.062329e-006, 1.339863e-006, 1.332288e-006, 1.156081e-006, 
    1.133854e-006, 9.98999e-007, 3.904106e-007, -7.785911e-008, 4.75593e-008, 
    4.893791e-007, 8.229167e-007, 1.014272e-006, 8.527186e-007, 
    5.453826e-007, 3.142904e-007, 1.600633e-007, 1.34359e-007,
  7.220856e-007, 5.851191e-007, 6.028761e-007, 7.527572e-007, 1.055995e-006, 
    1.09151e-006, 1.051153e-006, 1.045937e-006, 1.082693e-006, 1.278147e-006, 
    1.415858e-006, 1.51073e-006, 1.593928e-006, 1.446406e-006, 1.095732e-006, 
    8.930764e-007, 6.519259e-007, 5.309779e-007, 4.857778e-007, 
    5.491079e-007, 7.774679e-007, 7.941078e-007, 7.516394e-007, 
    7.169942e-007, 5.140901e-007, 3.222376e-007, 3.911555e-008, 
    -1.103926e-007, 8.506095e-008, 3.190091e-007, 2.621362e-007, 
    1.70121e-008, 5.50101e-008, 2.197921e-007, 4.764647e-007, 1.023462e-006, 
    1.963476e-006, 2.489984e-006, 2.508859e-006, 2.300739e-006, 
    2.332777e-006, 2.89008e-006, 3.670528e-006, 4.169593e-006, 4.078572e-006, 
    3.673757e-006, 4.314507e-006, 5.763149e-006, 6.029506e-006, 
    4.836545e-006, 4.004066e-006, 4.493818e-006, 4.918625e-006, 
    3.911679e-006, 2.145272e-006, 4.56721e-007, 3.001351e-007, 1.471117e-006, 
    3.070385e-006, 3.938625e-006, 3.543621e-006, 2.64359e-006, 2.531086e-006, 
    2.362331e-006, 2.235174e-006, 1.703203e-006, 7.54495e-007, 
    -2.135857e-008, 4.325047e-007, 1.732011e-006, 2.049033e-006, 
    1.211962e-006, 2.332035e-007, 3.51667e-007, 7.869048e-007, 1.078844e-006, 
    1.447896e-006, 2.27193e-006, 2.571692e-006, 2.385552e-006, 2.452607e-006, 
    2.224495e-006, 1.966457e-006, 1.687805e-006, 1.569962e-006, 
    1.295283e-006, 5.610282e-007, 2.550587e-007, 4.687663e-007, 
    1.336138e-006, 1.775101e-006, 1.551708e-006, 1.303975e-006, 
    1.220157e-006, 9.207679e-007, 6.804862e-007,
  3.070757e-006, 3.182143e-006, 3.526236e-006, 4.130478e-006, 4.890437e-006, 
    5.049258e-006, 5.034605e-006, 4.612531e-006, 3.682449e-006, 
    3.033629e-006, 3.411e-006, 4.880502e-006, 5.366404e-006, 4.617994e-006, 
    4.048024e-006, 3.686174e-006, 3.047785e-006, 2.215306e-006, 
    1.441811e-006, 1.594424e-006, 2.346312e-006, 2.985944e-006, 
    3.091991e-006, 3.067404e-006, 2.907714e-006, 2.183393e-006, 
    1.561642e-006, 1.647075e-006, 1.97577e-006, 1.630684e-006, 4.054364e-007, 
    -4.034491e-007, -5.014244e-007, -1.459075e-007, -1.134977e-007, 
    8.787956e-007, 2.852456e-006, 5.288794e-006, 6.828704e-006, 
    7.625917e-006, 7.651623e-006, 7.071347e-006, 5.541246e-006, 
    4.795442e-006, 4.512196e-006, 4.000962e-006, 4.457062e-006, 
    4.884849e-006, 5.624692e-006, 5.11743e-006, 3.931298e-006, 3.798306e-006, 
    4.675239e-006, 5.046153e-006, 3.965322e-006, 3.024066e-006, 2.70158e-006, 
    3.453842e-006, 4.161273e-006, 3.532692e-006, 3.250068e-006, 
    2.969678e-006, 2.215555e-006, 1.962607e-006, 2.78751e-006, 3.717344e-006, 
    2.363571e-006, 1.319002e-006, 1.780812e-006, 2.217665e-006, 
    1.681101e-006, 2.18836e-006, 2.096594e-006, 1.21519e-006, 2.150609e-006, 
    3.470728e-006, 4.055228e-006, 3.759315e-006, 3.556907e-006, 
    2.310177e-006, 1.539289e-006, 1.507749e-006, 1.77299e-006, 1.680231e-006, 
    1.862645e-006, 1.173343e-006, 1.635279e-006, 2.46726e-006, 2.559771e-006, 
    2.294655e-006, 2.12056e-006, 1.302611e-006, 9.955211e-007, 1.848986e-006, 
    2.379344e-006, 2.591684e-006,
  2.595782e-006, 3.24063e-006, 4.790723e-006, 5.974745e-006, 6.35162e-006, 
    5.808226e-006, 4.884725e-006, 4.165744e-006, 3.953775e-006, 
    4.026169e-006, 4.472708e-006, 4.606072e-006, 5.27526e-006, 5.988779e-006, 
    6.021932e-006, 7.577861e-006, 8.739531e-006, 7.40476e-006, 4.609054e-006, 
    4.067148e-006, 4.58074e-006, 4.072612e-006, 2.310922e-006, 1.661107e-006, 
    3.241872e-006, 5.225216e-006, 5.053605e-006, 4.177167e-006, 4.98568e-006, 
    4.895527e-006, 4.18797e-006, 2.998859e-006, 1.572322e-006, 1.717979e-006, 
    2.670162e-006, 1.429642e-006, 8.307325e-008, 1.715991e-006, 
    4.442285e-006, 4.198653e-006, 2.23505e-006, 1.880027e-006, 2.39176e-006, 
    3.322835e-006, 4.341206e-006, 5.973629e-006, 6.046395e-006, 
    4.895031e-006, 4.875536e-006, 5.035476e-006, 4.649162e-006, 
    3.845369e-006, 2.078961e-006, 2.521898e-006, 4.037967e-006, 
    4.280233e-006, 4.555781e-006, 4.493197e-006, 4.202377e-006, 3.84425e-006, 
    3.008792e-006, 1.784911e-006, 1.747036e-006, 3.225356e-006, 
    3.645942e-006, 3.787502e-006, 3.985191e-006, 3.280864e-006, 
    2.332778e-006, 2.984951e-006, 3.60695e-006, 4.107629e-006, 2.955025e-006, 
    1.337254e-006, 1.099705e-006, 3.448386e-007, 2.067783e-006, 2.00011e-006, 
    1.861032e-006, 1.798073e-006, 1.781185e-006, 2.286086e-006, 
    2.658491e-006, 2.864624e-006, 2.454345e-006, 2.317876e-006, 3.1434e-006, 
    3.27391e-006, 2.472102e-006, 2.154087e-006, 2.102926e-006, 2.104788e-006, 
    2.289687e-006, 2.204627e-006, 2.589324e-006, 2.673889e-006,
  2.277146e-006, 2.528355e-006, 2.362331e-006, 2.641975e-006, 3.526484e-006, 
    4.575029e-006, 4.901985e-006, 4.626561e-006, 5.326048e-006, 
    6.052604e-006, 4.817546e-006, 4.311776e-006, 3.994381e-006, 
    5.527088e-006, 7.156532e-006, 6.585196e-006, 5.201997e-006, 
    4.589187e-006, 5.382051e-006, 6.294125e-006, 6.351123e-006, 
    5.453701e-006, 4.264837e-006, 4.459545e-006, 4.992882e-006, 4.46501e-006, 
    6.298969e-006, 7.806966e-006, 6.799897e-006, 3.977244e-006, 
    3.304705e-006, 5.169461e-006, 4.803887e-006, 2.391636e-006, 
    1.888598e-006, 3.189343e-006, 4.399693e-006, 6.150207e-006, 
    6.216267e-006, 8.189183e-006, 7.742145e-006, 6.732842e-006, 
    5.028645e-006, 3.602232e-006, 3.529587e-006, 6.005044e-006, 
    5.715588e-006, 4.25602e-006, 4.926946e-006, 5.883972e-006, 6.446366e-006, 
    5.391365e-006, 3.819539e-006, 2.618879e-006, 2.629435e-006, 
    1.904989e-006, 1.443177e-006, 2.607703e-006, 3.867348e-006, 
    4.351015e-006, 3.932913e-006, 3.689651e-006, 3.883739e-006, 
    5.083779e-006, 3.332272e-006, 4.665306e-006, 3.290301e-006, 
    3.358226e-006, 3.385792e-006, 2.981598e-006, 2.848854e-006, 
    2.381206e-006, 3.754969e-006, 5.109485e-006, 5.125006e-006, 
    4.041443e-006, 3.71014e-006, 3.130983e-006, 4.746889e-006, 5.971267e-006, 
    5.387514e-006, 4.337604e-006, 4.477675e-006, 4.880751e-006, 
    4.636745e-006, 4.014497e-006, 4.282096e-006, 4.166241e-006, 
    4.299482e-006, 3.187482e-006, 2.04655e-006, 9.980049e-007, 4.582034e-008, 
    1.488879e-007, 9.98627e-007, 1.804779e-006,
  4.357098e-006, 4.136189e-006, 2.815575e-006, 3.314266e-006, 4.91167e-006, 
    5.358581e-006, 6.135428e-006, 5.541868e-006, 5.672995e-006, 
    5.978471e-006, 6.183363e-006, 6.129841e-006, 5.311147e-006, 
    4.427258e-006, 5.55031e-006, 6.974364e-006, 7.83615e-006, 9.631862e-006, 
    1.027696e-005, 9.219348e-006, 8.691848e-006, 9.687992e-006, 
    1.150059e-005, 1.049824e-005, 8.92207e-006, 9.588026e-006, 1.002389e-005, 
    7.972123e-006, 6.518885e-006, 6.976599e-006, 6.011376e-006, 
    4.782405e-006, 4.030515e-006, 3.324945e-006, 3.248078e-006, 
    4.257388e-006, 5.358208e-006, 5.772585e-006, 5.183618e-006, 
    5.220747e-006, 4.026911e-006, 1.936034e-006, 3.949304e-006, 
    6.359567e-006, 6.414577e-006, 6.612887e-006, 7.332364e-006, 5.39571e-006, 
    6.201368e-006, 5.925447e-006, 4.333506e-006, 3.738453e-006, 
    2.516557e-006, 2.680843e-006, 3.391877e-006, 2.859035e-006, 
    4.502137e-006, 4.0669e-006, 2.14912e-006, 9.218857e-007, 2.043695e-006, 
    2.597024e-006, 3.358473e-006, 2.94745e-006, 4.549325e-006, 5.064656e-006, 
    2.790242e-006, 2.367173e-006, 2.776211e-006, 2.119938e-006, 
    4.489595e-006, 4.881993e-006, 4.029771e-006, 4.50313e-006, 4.038959e-006, 
    4.451596e-006, 3.662706e-006, 2.851211e-006, 2.563993e-006, 
    5.118922e-006, 6.072843e-006, 6.590657e-006, 6.673858e-006, 
    5.606065e-006, 4.935637e-006, 4.540136e-006, 4.708643e-006, 
    4.757196e-006, 4.649162e-006, 2.699968e-006, 1.21817e-006, 1.210843e-006, 
    2.139932e-006, 2.166504e-006, 1.433988e-006, 1.806144e-006,
  4.709511e-006, 5.124883e-006, 6.206581e-006, 6.310642e-006, 7.684281e-006, 
    6.45953e-006, 5.714472e-006, 6.062786e-006, 5.244339e-006, 4.701316e-006, 
    5.264581e-006, 4.586949e-006, 3.14787e-006, 7.674967e-006, 1.089014e-005, 
    1.168822e-005, 1.373837e-005, 1.387199e-005, 1.323794e-005, 
    1.232562e-005, 1.202586e-005, 9.31571e-006, 9.271005e-006, 9.374693e-006, 
    8.32056e-006, 6.396942e-006, 6.127233e-006, 6.048507e-006, 6.757429e-006, 
    5.793696e-006, 4.034118e-006, 1.933797e-006, 2.944842e-006, 4.22063e-006, 
    6.376329e-006, 6.281338e-006, 4.774458e-006, 2.874061e-006, 
    2.211455e-006, 4.861133e-006, 4.610294e-006, 2.589448e-006, 3.91379e-006, 
    7.678074e-006, 8.219355e-006, 6.808588e-006, 5.653128e-006, 
    6.402533e-006, 4.220754e-006, -1.153101e-006, -7.538747e-007, 
    5.82264e-007, 1.163655e-006, 1.371403e-006, 5.101156e-007, 1.989181e-006, 
    2.318497e-006, 9.609994e-007, -9.362884e-008, -1.884129e-006, 
    2.463412e-006, 3.749379e-006, 1.370783e-006, -4.38964e-007, 
    1.703451e-006, 2.814333e-006, 1.42629e-006, 1.130253e-006, 2.317753e-006, 
    4.152083e-006, 3.441921e-006, 3.924344e-006, 5.046279e-006, 
    3.575409e-006, 1.780936e-006, 3.374244e-006, 6.338581e-006, 
    5.040814e-006, 3.457069e-006, 2.138813e-006, 1.203765e-006, 
    3.199777e-006, 3.538033e-006, 3.38306e-006, 2.949437e-006, 3.567462e-006, 
    3.160785e-006, 2.408151e-006, 1.607834e-006, 1.105418e-006, 
    4.147478e-008, 1.562386e-006, 9.570267e-007, 1.676628e-006, 
    3.954025e-006, 4.370138e-006,
  7.043283e-006, 6.791946e-006, 4.888574e-006, 5.510203e-006, 3.72529e-006, 
    3.674751e-006, 3.098572e-006, 4.230191e-006, 5.548696e-006, 
    9.436782e-006, 1.040461e-005, 1.219685e-005, 1.516032e-005, 
    1.525854e-005, 1.495096e-005, 1.542816e-005, 1.266946e-005, 
    9.747841e-006, 9.195879e-006, 8.812425e-006, 7.912269e-006, 
    9.272993e-006, 9.883694e-006, 1.020854e-005, 9.030726e-006, 
    8.198866e-006, 5.68926e-006, 4.569069e-006, 5.481765e-006, 4.6735e-006, 
    4.995614e-006, 2.479428e-006, 8.282586e-007, 3.090718e-007, 
    5.298607e-007, 6.498121e-007, 3.982212e-006, 3.863744e-006, 
    4.128851e-007, 1.63155e-006, 4.979596e-006, 5.246078e-006, 4.494934e-006, 
    5.051368e-006, 4.459172e-006, 4.864609e-006, 3.975008e-006, 
    4.260366e-006, 3.22461e-006, 2.225224e-007, 2.318744e-006, 5.133821e-006, 
    6.222725e-006, 2.089888e-006, 2.507617e-006, 3.80116e-006, 2.143781e-006, 
    2.596535e-007, -1.552826e-006, -2.684941e-006, -1.974331e-008, 
    1.479313e-006, 1.958251e-007, -1.473982e-007, 3.277011e-006, 
    2.672276e-006, 9.396426e-007, -1.337357e-007, 5.8363e-007, 1.911445e-006, 
    2.846991e-006, 3.123783e-006, 1.523149e-006, 6.695591e-007, 
    3.610425e-006, 7.195522e-006, 7.993851e-006, 5.329897e-006, 
    2.819548e-006, 1.005208e-006, -8.703519e-007, -2.133349e-006, 
    -1.762435e-006, -1.310433e-006, -6.895516e-007, 1.265729e-006, 
    1.742566e-006, 1.082819e-006, 2.439443e-006, 4.06963e-006, 2.817935e-006, 
    2.992278e-006, 4.149231e-006, 4.384045e-006, 5.540252e-006, 5.373731e-006,
  4.696227e-006, 5.265698e-006, 4.494563e-006, 5.067013e-006, 6.138158e-006, 
    6.673734e-006, 8.185456e-006, 1.065396e-005, 1.111614e-005, 
    1.013416e-005, 1.070077e-005, 1.176074e-005, 1.375911e-005, 
    1.406496e-005, 1.072871e-005, 6.001443e-006, 3.495068e-006, 
    3.318364e-006, 5.61749e-006, 6.786484e-006, 9.005889e-006, 1.098054e-005, 
    9.416042e-006, 6.199505e-006, 3.054614e-006, 1.789009e-006, 
    2.474339e-006, 2.305584e-006, 8.117386e-007, -6.895534e-007, 
    -3.551319e-006, -4.379202e-006, -2.700588e-006, -1.547112e-006, 
    3.899186e-008, 1.615263e-009, -2.049528e-006, -3.224734e-006, 
    -1.860037e-006, 1.3647e-006, 4.827729e-006, 5.224969e-006, 2.91889e-006, 
    1.588216e-006, 6.011625e-006, 5.340575e-006, 3.325194e-006, 
    3.753848e-007, 1.388789e-006, 4.574533e-006, 4.262105e-006, 
    5.858763e-006, 5.550683e-006, 4.07733e-006, 1.082073e-006, 1.01325e-007, 
    -1.542021e-006, -3.824134e-006, -6.049624e-006, -6.548442e-006, 
    -4.003941e-006, -1.412631e-006, -1.892196e-006, -2.075732e-006, 
    -1.750886e-007, 9.175383e-007, -1.36271e-006, 2.970301e-007, 
    1.784909e-006, 1.070275e-006, -1.086792e-006, -3.735222e-007, 
    1.739711e-006, 1.164899e-006, 5.212674e-006, 9.205196e-006, 
    7.264563e-006, 4.473452e-006, 9.914238e-007, 4.557296e-008, 
    -2.821289e-007, -8.489933e-007, -5.654983e-007, -4.780668e-008, 
    -2.484776e-007, 5.741913e-007, 1.055127e-006, 1.136836e-006, 
    3.130488e-006, 5.319343e-006, 3.398211e-006, 4.541005e-006, 
    5.684171e-006, 6.093705e-006, 5.592781e-006, 4.702062e-006,
  9.19824e-006, 5.533049e-006, 6.113201e-006, 6.883965e-006, 7.133556e-006, 
    8.634728e-006, 1.064179e-005, 1.306881e-005, 1.384442e-005, 
    1.283921e-005, 1.625059e-005, 1.955281e-005, 1.545846e-005, 
    8.870536e-006, 6.247437e-006, 7.321438e-006, 6.589169e-006, 
    4.388516e-006, 3.993884e-006, 5.067266e-006, 5.392732e-006, 
    6.014732e-006, 3.415345e-006, -5.575494e-007, -4.390629e-006, 
    -4.711994e-006, -5.324684e-006, -7.226441e-006, -7.880728e-006, 
    -7.292503e-006, -5.517773e-006, -3.234421e-006, -9.412579e-007, 
    -2.012526e-006, -2.772485e-006, -1.584365e-006, -1.128017e-006, 
    -7.613271e-007, 5.863585e-007, 2.94832e-006, 4.026171e-006, 
    5.825486e-006, 2.268453e-006, 6.160388e-006, 6.671868e-006, 
    7.196515e-006, 5.492941e-006, 2.168988e-006, 3.700579e-006, 
    6.337465e-006, 5.680198e-006, 4.595768e-006, 3.924721e-006, 
    2.882753e-006, 1.6585e-006, 2.580386e-006, 8.032985e-007, -4.662943e-006, 
    -2.617515e-006, -2.241508e-006, 8.010611e-007, -3.437079e-006, 
    -2.663583e-006, -1.919892e-006, -5.854927e-007, -2.22549e-006, 
    -2.203014e-006, 4.02455e-007, -4.651629e-007, -3.296882e-006, 
    -1.111999e-006, 1.620501e-007, 1.661851e-006, 5.820148e-006, 
    5.701062e-006, 5.8152e-007, -3.774963e-006, -5.689762e-007, 
    -2.522029e-007, 1.374632e-006, 1.306584e-006, 2.29838e-006, 
    3.395353e-006, 3.045425e-006, 4.278743e-006, 4.642334e-006, 2.36059e-006, 
    4.32556e-006, 5.386148e-006, 5.302081e-006, 4.599864e-006, 3.9724e-006, 
    4.615013e-006, 3.649293e-006, 4.082423e-006, 8.455168e-006,
  3.013265e-006, 2.111992e-006, 4.207344e-006, 1.822042e-006, 2.062819e-006, 
    4.964941e-006, 7.324417e-006, 6.596991e-006, 4.826859e-006, 
    7.587794e-006, 8.469695e-006, 1.768021e-006, -5.96543e-006, 
    -4.876776e-006, -4.585832e-006, -3.43534e-006, -1.440694e-006, 
    -7.389717e-007, -1.348555e-006, -2.615401e-006, -3.426525e-006, 
    -4.701316e-006, -1.057821e-005, -1.280842e-005, -1.113092e-005, 
    -9.257468e-006, -7.624054e-006, -7.195647e-006, -6.367638e-006, 
    -3.49221e-006, -4.182135e-006, -4.57354e-006, -5.072852e-006, 
    -6.498769e-006, -5.440663e-006, -2.429137e-006, -2.334491e-008, 
    1.31776e-006, 2.130491e-006, 3.462783e-006, 1.558785e-006, 7.910039e-007, 
    2.674758e-006, 7.116792e-006, 5.439546e-006, 5.990143e-006, 7.3007e-006, 
    3.201512e-006, 2.056484e-006, -2.584235e-006, -6.735321e-006, 
    -3.161778e-006, 2.892048e-007, 1.704568e-006, -1.147015e-006, 
    -3.147623e-006, -2.523513e-006, -3.477908e-009, -1.072636e-006, 
    -6.599228e-006, -6.07632e-006, -2.543631e-006, -4.210815e-007, 
    7.758536e-007, -2.387536e-006, 1.608096e-007, 2.75411e-006, 
    3.586461e-006, 3.401437e-006, 5.550555e-006, -1.246735e-007, 
    1.332166e-006, -1.528857e-006, 2.145789e-007, 5.618967e-007, 
    -4.352503e-006, -6.223221e-006, -4.702932e-006, 9.546675e-007, 
    2.363447e-006, 2.458071e-006, 4.956126e-006, 6.015101e-006, 
    1.076013e-005, 1.117897e-005, 9.389467e-006, 8.275234e-006, 
    7.273877e-006, 4.336114e-006, 4.792961e-006, 5.061182e-006, 
    3.588571e-006, 2.881265e-006, 3.054116e-006, 4.118308e-006, 3.841145e-006,
  -1.069158e-006, -1.381586e-006, -4.364549e-006, -4.404534e-006, 
    -2.051393e-006, -2.337869e-006, -1.384193e-006, -2.609069e-006, 
    -1.836195e-006, -2.311916e-006, -9.897973e-006, -1.291521e-005, 
    -1.253299e-005, -1.13635e-005, -8.274365e-006, -6.163616e-006, 
    -6.656473e-006, -6.751965e-006, -8.688743e-006, -8.023902e-006, 
    -9.537489e-006, -1.025485e-005, -8.567547e-006, -5.121157e-006, 
    -5.008405e-006, -5.173186e-006, -3.078829e-006, -2.321105e-006, 
    -1.894807e-006, -1.331171e-006, -2.355624e-006, -6.356837e-006, 
    -5.344922e-006, -4.059571e-006, -2.121677e-006, 1.37712e-007, 
    5.738184e-007, 8.645147e-007, 2.864748e-006, 3.709767e-006, 
    6.064774e-007, 2.334889e-006, 1.097173e-005, 1.413996e-005, 
    6.265691e-006, 3.794332e-006, 5.183101e-007, -4.205976e-006, 
    -7.364404e-006, -1.667428e-005, -1.729553e-005, -8.246177e-006, 
    -3.459056e-006, -6.061793e-006, -6.92283e-006, -3.847479e-006, 
    -1.182034e-006, -4.136811e-006, -3.753725e-006, -5.068381e-006, 
    -4.502512e-006, -5.447655e-007, 2.053501e-006, 2.973029e-006, 
    6.229802e-006, 8.224946e-006, 9.403499e-006, 5.735958e-006, 6.47211e-007, 
    -2.805391e-006, -3.077341e-006, -4.219637e-006, -4.57155e-006, 
    -3.928191e-006, -1.09573e-006, -6.345363e-008, -2.235547e-006, 
    -1.864631e-006, -8.805346e-007, 9.369105e-007, 2.171098e-006, 
    6.850809e-006, 1.580566e-005, 9.281812e-006, 7.446113e-006, 2.56933e-006, 
    -2.65762e-006, -5.469348e-006, -5.404156e-006, -4.570931e-006, 
    -3.456818e-006, -2.900884e-006, -1.480432e-006, -8.637726e-007, 
    -1.804157e-006, -6.755199e-007,
  -4.595891e-006, -5.4614e-006, -6.131207e-006, -3.96582e-006, 
    -2.394617e-006, -1.203641e-006, -2.938509e-006, -1.350418e-006, 
    -1.143664e-006, -4.575402e-006, -1.004959e-005, -7.991617e-006, 
    -8.744995e-006, -1.516727e-005, -1.29121e-005, -7.373093e-006, 
    -6.507462e-006, -8.285044e-006, -6.489952e-006, -7.163857e-006, 
    -5.426133e-006, -1.737475e-006, -1.707922e-006, -2.418583e-006, 
    -3.360219e-007, -3.239747e-007, 1.05761e-006, 1.923243e-006, 
    3.409878e-007, -6.56768e-007, -4.386529e-006, -9.96888e-007, 
    1.309936e-006, 1.153474e-006, 1.951183e-006, 2.619376e-006, 
    1.452615e-006, 5.140901e-007, 2.260878e-006, 3.072867e-006, 
    2.707541e-006, 5.351132e-006, 6.730483e-006, 1.824646e-006, 
    -3.962097e-006, -7.381412e-006, -1.122964e-005, -1.253709e-005, 
    -1.127024e-005, -1.241503e-005, -1.285387e-005, -1.074622e-005, 
    -1.012459e-005, -7.099785e-006, -1.018234e-005, -8.570401e-006, 
    -5.703048e-006, -1.756103e-006, -5.85118e-007, 1.763554e-006, 
    2.311921e-006, 6.80946e-006, 8.159623e-006, 1.090629e-005, 1.095074e-005, 
    1.284617e-005, 1.126925e-005, 7.58854e-006, -2.338489e-006, 
    -6.827588e-006, -8.830801e-006, -9.101257e-006, -4.375601e-006, 
    -1.223385e-006, -1.764919e-006, -1.499678e-006, -1.163408e-006, 
    -9.683263e-007, 1.00943e-006, 6.262217e-007, 6.638715e-006, 
    9.115909e-006, 3.766268e-006, -3.298994e-006, -5.73943e-006, 
    -5.559623e-006, -8.802612e-006, -7.484854e-006, -4.654377e-006, 
    -6.499886e-006, -6.577373e-006, -4.789481e-006, -4.301097e-006, 
    -3.230447e-006, -2.105658e-006, -2.318497e-006,
  -2.968684e-006, -2.332528e-006, -1.99303e-006, -1.587222e-006, 
    -1.315896e-006, -1.658251e-006, -2.099325e-006, -5.690753e-006, 
    -5.424146e-006, -4.922474e-006, -8.774672e-006, -7.179753e-006, 
    -7.758288e-006, -1.573488e-005, -7.970009e-006, -3.424784e-006, 
    -1.018743e-005, -1.166041e-005, -8.434679e-006, -6.681681e-006, 
    -3.65364e-006, -5.601596e-007, -1.983717e-006, -3.71697e-006, 
    -2.140056e-006, 1.351535e-006, 1.455099e-006, 2.18091e-006, 
    1.423557e-006, -1.140312e-006, -1.84017e-006, 4.469111e-007, 
    8.245315e-007, 1.122429e-006, 7.738672e-007, -1.245489e-007, 
    1.174708e-006, 1.070524e-006, 2.224123e-006, 2.931803e-006, 
    5.694727e-006, 4.028654e-006, -3.87927e-006, -6.681557e-006, 
    -1.064974e-005, -7.711229e-006, -9.078532e-006, -5.184611e-006, 
    -7.733703e-006, -1.303144e-005, -1.419956e-005, -1.579238e-005, 
    -1.679944e-005, -1.617484e-005, -1.343675e-005, -8.570401e-006, 
    -5.273767e-006, 1.848613e-006, 2.770499e-006, 6.18659e-006, 
    1.412754e-005, 1.275614e-005, 1.003482e-005, 1.310544e-005, 
    1.002712e-005, 8.703893e-006, 6.876886e-006, 2.863133e-006, 
    -2.491099e-006, -6.173797e-006, -5.709133e-006, -3.900504e-006, 
    -1.848985e-006, -3.311037e-006, -1.739462e-006, -8.313609e-007, 
    8.108714e-007, 1.194825e-006, 7.21092e-007, -3.493453e-006, 
    3.349161e-006, -4.229572e-006, -4.697093e-006, -1.597156e-006, 
    -4.286567e-006, -7.669752e-006, -9.808937e-006, -8.325404e-006, 
    -6.17293e-006, -6.361181e-006, -6.546081e-006, -5.240366e-006, 
    -5.226458e-006, -3.494695e-006, -3.249199e-006, -4.512444e-006,
  -1.24611e-006, -9.886926e-007, -3.422301e-007, -6.304433e-007, 
    -7.138897e-007, -1.566857e-006, -2.594168e-006, -2.468502e-006, 
    -3.503139e-006, -3.271549e-006, -7.442633e-006, -3.673012e-006, 
    -9.814894e-007, -3.705174e-006, -7.164603e-006, -8.943429e-006, 
    -9.427094e-006, -9.074683e-006, -1.035295e-005, -9.440382e-006, 
    -2.837305e-006, -2.106528e-006, -1.906605e-006, -1.184517e-006, 
    1.380593e-006, 1.225621e-006, 1.798197e-006, 1.75722e-006, 8.929519e-007, 
    -1.561642e-006, -3.169477e-006, -2.62633e-006, -1.339118e-006, 
    1.281997e-006, 1.453857e-006, 1.63267e-006, 4.031758e-006, 3.886968e-006, 
    1.496077e-006, 4.766013e-006, 4.40913e-006, -1.232078e-006, 
    -4.394476e-006, -4.951407e-006, -3.557156e-006, -1.600756e-006, 
    -6.250664e-006, -1.17174e-005, -1.692722e-005, -1.907634e-005, 
    -2.025043e-005, -1.498746e-005, -1.133718e-005, -8.923562e-006, 
    -4.409128e-006, 3.819663e-006, 7.862847e-006, 8.372343e-006, 
    8.513282e-006, 1.306894e-005, 1.212048e-005, 1.250729e-005, 
    1.240708e-005, 9.861338e-006, 8.28554e-006, 3.650786e-006, 
    -1.050539e-007, -2.187116e-006, -3.294646e-006, -2.773727e-006, 
    -2.258023e-006, -1.313289e-006, -1.322478e-006, -2.828738e-007, 
    -1.12839e-006, 3.562618e-007, 1.627083e-006, 1.809249e-006, 
    7.939834e-007, -1.650926e-006, -3.059333e-006, -6.610404e-006, 
    -4.292528e-006, -3.747394e-006, -2.355377e-006, -3.130237e-006, 
    -7.951383e-006, -4.031012e-006, -3.023321e-006, -1.634408e-006, 
    -2.71077e-006, -1.977011e-006, -6.665787e-007, -1.340483e-006, 
    -3.130362e-006, -1.779447e-006,
  -5.607808e-007, -8.620323e-007, -5.972881e-007, -2.107273e-007, 
    -4.248073e-007, -1.594797e-006, -1.605973e-006, -1.025945e-006, 
    -1.752376e-006, -9.371588e-007, -1.930321e-006, -1.116346e-006, 
    -9.400146e-007, -2.785897e-006, -6.021932e-006, -9.425106e-006, 
    -6.089111e-006, -7.583822e-006, -9.264675e-006, -3.667672e-006, 
    -4.407011e-007, -2.029046e-007, 3.70419e-007, 1.763292e-007, 
    1.617893e-006, 1.457707e-006, 2.176803e-007, 1.061708e-007, 
    -1.276159e-006, -2.520779e-006, -2.285714e-006, 1.64534e-007, 
    1.480679e-006, 8.369486e-007, 1.165022e-006, 1.301368e-006, 
    2.283851e-006, 1.691406e-006, 2.233933e-006, 1.995266e-006, 
    9.648556e-008, -9.525575e-007, -1.767278e-006, -6.688133e-007, 
    1.875311e-006, -9.981304e-007, -7.504101e-006, -1.337628e-005, 
    -1.334834e-005, -7.515897e-006, -8.888543e-006, -7.200611e-006, 
    -4.917631e-006, 3.995992e-007, 6.387134e-006, 8.591262e-006, 
    5.006295e-006, 3.849713e-006, 7.501993e-006, 9.179239e-006, 
    8.413941e-006, 1.114445e-005, 8.184959e-006, 2.349292e-006, 
    -3.617261e-007, -3.427143e-006, -3.612911e-006, -2.732625e-006, 
    -2.19283e-006, -1.86401e-006, -1.768643e-006, -6.102027e-007, 
    3.864361e-007, -5.643815e-007, -5.924455e-007, 1.151115e-006, 
    1.007815e-006, 8.232892e-007, -3.115583e-007, -2.282983e-006, 
    -3.048529e-006, -4.172326e-006, -2.741565e-006, -3.044804e-006, 
    -3.220886e-006, -1.314282e-006, -1.868979e-006, 1.075989e-006, 
    1.312668e-006, -1.394625e-006, -9.611176e-008, 7.295366e-007, 
    -3.028672e-007, -2.925599e-007, -1.459321e-006, -7.13766e-007,
  -1.806641e-006, -2.353265e-006, -8.085121e-007, -1.228104e-007, 
    -3.490597e-007, -8.496145e-007, -4.200886e-007, -3.052255e-007, 
    -1.172349e-006, 2.454963e-007, -6.618593e-007, 2.399083e-007, 
    -2.8722e-007, -1.253809e-006, -5.214786e-006, -7.7604e-006, 
    -5.250797e-006, -4.517535e-006, -3.540639e-006, -1.486405e-007, 
    2.973278e-006, 2.777078e-006, -3.714122e-007, 1.046186e-006, 
    2.502155e-006, 2.696986e-006, -5.986531e-007, -1.261384e-006, 
    -2.516061e-006, -7.52384e-007, -1.163535e-007, -7.102881e-008, 
    7.787098e-007, 4.0705e-007, 6.421158e-007, 9.545436e-007, 6.043663e-007, 
    1.0026e-006, 7.258104e-007, -9.393934e-007, 1.752123e-007, 4.927315e-007, 
    8.635216e-007, 4.173318e-006, 1.158442e-006, -6.447483e-006, 
    -8.335708e-006, -4.067022e-006, -4.997601e-006, -7.615861e-006, 
    -5.79233e-006, -3.205612e-006, 1.168872e-006, 6.119657e-006, 
    5.64605e-006, 3.801659e-006, 6.819393e-006, 7.314733e-006, 5.958977e-006, 
    4.081925e-006, 4.669775e-006, 1.809125e-006, -2.101685e-006, 
    -2.818058e-006, -4.922226e-006, -3.530706e-006, -3.045798e-006, 
    -2.000109e-006, -2.089639e-006, -2.805267e-006, -8.573143e-007, 
    -2.445031e-007, -5.221614e-007, -1.64099e-006, 2.673519e-007, 
    8.54209e-007, 2.469867e-007, -4.527471e-007, -7.785857e-007, 
    -3.57367e-006, -1.862894e-006, -5.71087e-007, -1.305342e-006, 
    -1.128142e-006, -3.846363e-006, -5.089492e-006, -1.755356e-006, 
    1.948823e-006, 7.232029e-007, 8.296211e-007, 1.196316e-006, 
    -1.924727e-007, -6.474547e-007, -1.062825e-006, -7.104127e-007, 
    -6.390119e-007,
  -1.6282e-006, -1.699602e-006, -7.023414e-007, -2.320856e-007, 
    -1.210719e-007, -5.657474e-007, -9.164214e-008, -3.116827e-008, 
    -7.188569e-007, -3.290643e-008, -7.198496e-007, -6.022492e-008, 
    -5.06267e-007, -1.396859e-006, -3.068893e-006, -2.097586e-006, 
    -4.634257e-007, 8.476272e-007, 2.233808e-006, 2.649798e-006, 
    3.433848e-006, 3.795698e-006, 2.984205e-006, 4.045043e-006, 
    5.206839e-006, 1.499679e-006, -9.451069e-007, -7.78582e-008, 
    2.678609e-006, 4.2667e-006, 6.830942e-007, 9.48583e-007, 5.827596e-007, 
    -4.222102e-009, -2.204131e-007, 4.775823e-007, -3.39995e-007, 
    1.062577e-006, 8.49368e-008, -7.585932e-007, 3.915653e-006, 
    6.045278e-006, 6.138411e-006, 5.481641e-006, -5.37435e-007, 
    -7.055947e-006, -1.005133e-005, -5.7326e-006, -8.389976e-006, 
    -4.181515e-006, -4.818139e-008, 2.155703e-006, 2.782668e-006, 
    3.977988e-006, 5.603706e-006, 6.697825e-006, 6.326165e-006, 
    4.546097e-006, 2.768635e-006, 1.560399e-006, 6.578857e-007, 1.41561e-007, 
    -1.931438e-006, -2.29155e-006, -3.013015e-006, -3.198908e-006, 
    -2.749141e-006, -2.914419e-006, -2.305457e-006, -2.311171e-006, 
    -1.997625e-006, -2.331908e-006, -1.860658e-006, -4.806866e-007, 
    2.827495e-007, 6.978712e-008, -4.557273e-007, -2.160596e-008, 
    -2.682085e-006, -1.303479e-006, -8.311122e-007, -9.924172e-007, 
    -1.438955e-006, -8.89475e-007, -1.735613e-006, -3.488362e-006, 
    -8.676216e-007, 2.958128e-006, 6.571408e-007, -2.976503e-007, 
    -1.22649e-006, -4.466374e-006, -2.430256e-006, -1.768271e-006, 
    -7.387243e-007, -2.232815e-006,
  -2.46341e-006, -1.605724e-006, -1.019487e-007, 1.311675e-006, 
    -1.303852e-008, -1.949569e-008, -6.08464e-009, 2.856056e-008, 
    -7.214641e-008, 1.785656e-007, -6.072196e-008, 7.157523e-007, 
    -1.859541e-006, -1.9261e-006, -1.255174e-006, -1.638879e-006, 
    -1.695504e-006, 6.942682e-007, 3.153333e-006, 3.869334e-006, 
    3.960478e-006, 4.956375e-006, 4.404039e-006, 5.517526e-006, 
    7.434188e-006, 3.366793e-006, 5.120659e-006, 9.778143e-006, 
    1.174087e-005, 1.182742e-005, 1.001283e-005, 6.7655e-006, 5.207085e-006, 
    2.79732e-006, 4.061311e-006, 1.882141e-006, 4.635006e-006, 4.909063e-006, 
    4.102165e-006, 1.507836e-005, 1.604334e-005, 2.159762e-005, 
    1.613572e-005, 1.63056e-006, -6.070233e-006, -5.95512e-006, 
    -2.053157e-005, -1.195992e-005, -9.1662e-006, -1.161818e-005, 
    -5.350015e-006, -4.255646e-006, -2.80614e-006, 2.807876e-006, 
    4.974008e-006, 4.727768e-006, 4.7264e-006, 6.544216e-006, 2.881015e-006, 
    2.159923e-006, 7.407116e-007, -4.856538e-007, -1.168872e-006, 
    -1.778702e-006, -2.475332e-006, -2.98433e-006, -2.461671e-006, 
    -2.421066e-006, -2.197176e-006, -2.830476e-006, -2.083183e-006, 
    -1.598398e-006, -1.706431e-006, -2.749264e-007, 2.04891e-008, 
    3.845744e-007, 1.326574e-006, 4.819281e-007, 1.354765e-007, 
    2.291054e-007, -1.21966e-006, -3.062189e-007, -1.342843e-006, 
    -7.102881e-008, 1.119574e-006, 2.146016e-006, 2.967863e-008, 
    2.760687e-006, -3.710393e-007, -3.540516e-006, -3.875543e-006, 
    -3.574664e-006, -1.449013e-006, 1.754606e-007, -2.031529e-007, 
    -1.974404e-006,
  -1.828e-006, 3.674379e-007, -1.154831e-008, -8.270172e-008, 1.789381e-007, 
    -3.474453e-007, 2.502153e-007, 8.481243e-008, 1.867612e-007, 
    3.856917e-007, 1.507501e-007, -3.116578e-006, -2.479057e-006, 
    -1.153971e-006, -3.200521e-006, -2.712632e-006, -4.23317e-007, 
    4.598747e-006, 7.2406e-006, 7.406496e-006, 5.764388e-006, 3.976125e-006, 
    4.849084e-006, 5.430855e-006, 1.085202e-005, 1.225024e-005, 
    1.972628e-005, 1.760001e-005, 6.760658e-006, 1.305876e-005, 
    1.383523e-005, 9.205316e-006, 7.760524e-006, 7.778778e-006, 
    8.320683e-006, 1.356316e-005, 2.645714e-005, 3.948298e-005, 
    9.325395e-006, 3.748759e-006, 1.925615e-005, 2.798501e-005, 
    3.028313e-005, 7.187569e-006, -1.067798e-006, 3.439185e-006, 
    -7.269649e-006, -8.046132e-006, 2.577646e-006, -2.094821e-007, 
    5.917995e-006, 1.247575e-005, 1.642964e-005, 1.88707e-005, 1.51217e-005, 
    1.360439e-005, 9.846315e-006, 7.637962e-006, 5.2426e-006, 3.857042e-006, 
    1.529853e-006, -1.075368e-007, -1.251201e-006, -1.736482e-006, 
    -2.354135e-006, -1.989553e-006, -2.191588e-006, -2.558281e-006, 
    -1.877298e-006, -1.811484e-006, -1.632174e-006, -1.588837e-006, 
    -6.007654e-007, -1.239277e-007, 1.794596e-006, 2.735108e-006, 
    3.922733e-007, 2.523139e-006, 5.953261e-006, 1.102562e-006, 
    6.519258e-007, 3.195055e-007, 9.067355e-007, 7.399667e-007, 
    3.400693e-006, 4.450728e-006, 5.662514e-008, 6.936498e-007, 
    1.075069e-005, 6.017834e-006, -1.399965e-006, -7.261709e-006, 
    6.218999e-006, 1.665328e-006, 6.152932e-007, -9.821106e-007,
  2.753734e-006, 1.834954e-006, 6.680689e-007, -7.014719e-007, 2.475207e-006, 
    9.385249e-007, 2.949191e-007, 1.983592e-006, 2.402067e-006, 
    1.323471e-006, 2.725919e-006, -1.88003e-006, -3.195679e-006, 
    -1.585111e-006, -1.918649e-006, -1.670422e-006, 2.203014e-006, 
    1.307068e-005, 1.141454e-005, 8.798394e-006, 1.118792e-005, 
    1.222503e-005, 1.581485e-005, 1.908019e-005, 2.05348e-005, 9.725867e-006, 
    1.518292e-005, 8.080653e-006, 4.665055e-006, 1.898395e-005, 8.22631e-006, 
    1.773536e-005, 1.360215e-005, 2.105894e-005, 2.17167e-005, 6.287792e-006, 
    5.057329e-006, 2.726354e-005, 2.999976e-006, 8.419902e-006, 
    3.469512e-005, 6.481874e-006, 1.148619e-005, 1.356825e-005, 
    2.762664e-005, 4.793803e-005, 4.625481e-005, 4.613114e-005, 
    5.388099e-005, 4.835601e-005, 4.560823e-005, 4.571764e-005, 
    3.165292e-005, 2.586283e-005, 1.7903e-005, 1.030502e-005, 5.884096e-006, 
    2.787511e-006, 1.401082e-006, -5.052739e-007, -9.036312e-007, 
    -1.431753e-006, -1.523768e-006, -1.743685e-006, -8.859979e-007, 
    -1.262873e-006, -9.95522e-007, -8.729598e-007, -1.352278e-007, 
    -3.580003e-007, -1.240523e-007, 3.650757e-008, 1.277774e-006, 
    1.549844e-006, 5.701184e-006, 5.8081e-006, 1.457085e-006, 3.922112e-006, 
    1.031794e-005, 8.933248e-007, 3.99823e-006, 2.958999e-006, 1.463791e-006, 
    2.192954e-006, 4.33003e-006, 6.887563e-006, 6.841619e-006, 1.271491e-005, 
    3.222451e-005, 2.309965e-005, -2.727909e-006, 3.368914e-007, 
    1.603812e-005, 6.058068e-006, 4.670272e-006, 3.889576e-006,
  5.156795e-006, 9.774914e-006, 8.237112e-006, 3.790235e-006, 1.096601e-005, 
    1.261185e-005, 8.347135e-006, 7.825343e-006, 4.670521e-006, 
    1.116258e-005, 4.210075e-006, -5.623947e-007, -1.403068e-006, 
    -2.662465e-006, -1.750637e-006, -2.921e-006, 1.461558e-007, 
    6.570048e-006, 7.895134e-006, 5.637608e-006, 7.768347e-006, 
    1.078322e-005, 1.377513e-005, 1.372645e-005, 1.521682e-005, 
    9.040163e-006, 1.002687e-005, 1.054356e-005, 1.255423e-005, 
    2.246089e-005, 3.584846e-006, 2.160582e-005, 1.212967e-005, 9.31236e-006, 
    1.490017e-005, 6.022179e-006, -1.061708e-007, 5.085887e-006, 
    1.713745e-005, 4.299943e-005, 3.707162e-005, 9.602431e-006, 2.30716e-005, 
    2.668623e-005, 2.641678e-005, 1.551856e-005, 1.749396e-005, 
    2.384124e-005, 2.150871e-005, 2.076266e-005, 2.803852e-005, 
    3.218526e-005, 2.810197e-005, 1.896521e-005, 1.438384e-005, 
    8.456906e-006, 6.160637e-006, 3.780921e-006, 1.85656e-006, 8.728352e-007, 
    4.791968e-007, -2.134589e-007, 3.1429e-007, -2.432616e-007, 
    -6.42116e-007, 2.187985e-007, -1.627955e-007, 8.617835e-007, 
    3.688001e-008, 3.253444e-008, 1.488875e-006, 1.823531e-006, 
    2.146387e-006, 5.2955e-006, 6.789713e-006, 1.449001e-005, 6.532169e-006, 
    1.106796e-005, 2.280598e-005, 5.307673e-006, -1.770506e-006, 
    -5.401671e-007, -3.570691e-006, -4.135443e-006, -9.650488e-006, 
    -1.173343e-005, -2.674175e-005, 1.747596e-005, -1.34647e-005, 
    -1.630193e-006, -1.36804e-006, 1.145626e-005, 3.850582e-006, 
    9.837997e-006, 5.170823e-006, 3.979603e-006,
  3.223373e-006, 1.775038e-005, 8.383518e-006, 1.066314e-005, 9.150055e-006, 
    1.782912e-005, 8.117535e-006, -7.456765e-007, 1.462671e-006, 
    8.001552e-006, 3.787871e-006, -1.363704e-006, -5.487352e-007, 
    -1.106659e-006, 1.291682e-006, 1.416978e-006, 8.611758e-006, 
    2.76044e-006, -3.388523e-006, -3.708155e-006, 6.852424e-006, 
    8.93548e-006, 1.289894e-005, 1.342396e-005, 1.256602e-005, 5.773953e-006, 
    4.297992e-006, 1.437714e-005, 4.145011e-006, 1.734748e-006, 
    -1.028602e-005, -8.350857e-006, -5.874412e-006, 4.383306e-006, 
    -3.634887e-006, -7.153183e-006, 5.906077e-006, 1.055276e-005, 
    1.57247e-005, 1.67222e-005, 5.372975e-006, 5.47232e-006, 1.016037e-005, 
    7.852053e-006, 1.967052e-005, 2.003883e-005, 7.666902e-006, 
    -1.236549e-006, 5.218513e-006, 1.209838e-005, 1.348469e-005, 
    1.869723e-005, 2.534216e-005, 2.094855e-005, 2.009298e-005, 
    2.043793e-005, 2.103883e-005, 1.937374e-005, 1.93607e-005, 1.606519e-005, 
    1.191696e-005, 1.026913e-005, 1.314891e-005, 7.535022e-006, 
    9.491418e-006, 8.696319e-006, 2.091427e-005, 1.434286e-005, 
    1.197656e-005, 1.752401e-005, 1.14462e-005, 1.310436e-006, 
    -8.713541e-007, 1.488865e-006, 1.501304e-005, 1.431852e-005, 
    1.093683e-005, 9.721145e-006, -1.047464e-005, -1.610518e-005, 
    -4.730622e-006, -5.902226e-006, -1.361223e-006, -4.8851e-006, 
    -9.06748e-006, -1.610753e-005, -3.362136e-005, -7.652488e-006, 
    -1.465057e-005, -1.071691e-005, 5.075708e-006, 8.42959e-006, 
    -1.983964e-006, -3.244975e-006, 6.221235e-007, -2.988178e-006,
  -6.537266e-006, -2.050401e-006, -4.372741e-006, -2.519537e-006, 
    1.009539e-007, 8.914649e-007, 2.544992e-006, 6.310656e-007, 
    -1.53482e-006, -2.400254e-005, -4.41884e-005, 2.10814e-006, 
    1.486392e-007, 4.7311e-008, 3.453342e-007, 3.394857e-006, 1.180991e-005, 
    9.638941e-006, 7.82236e-006, 9.752308e-006, 8.989002e-006, 9.9957e-006, 
    2.510821e-005, 2.954603e-005, 1.188951e-005, 2.081215e-007, 5.09368e-007, 
    5.964936e-006, -6.417686e-006, -1.236225e-005, -7.346149e-006, 
    -1.682216e-006, -4.667745e-007, 3.525864e-006, -5.911046e-006, 
    -1.550267e-005, 5.675247e-008, 2.994879e-006, 6.023671e-006, 
    8.448958e-006, 6.13444e-006, 1.008448e-007, -1.268162e-005, 
    -9.688229e-007, 8.716561e-006, 8.689858e-006, 1.731139e-006, 
    5.038084e-006, 1.321211e-005, 9.316951e-006, 7.047754e-006, 
    7.375827e-006, 8.21265e-006, 3.545858e-006, 6.302573e-006, 4.923466e-006, 
    1.660366e-006, 6.416936e-006, 1.398585e-005, 1.55069e-005, 1.938579e-005, 
    1.51823e-005, 9.787822e-006, 2.304339e-006, 2.539527e-006, 7.740658e-006, 
    2.47733e-005, -1.030567e-007, -1.681646e-005, -1.286529e-005, 
    -1.666423e-005, -4.701564e-006, -3.201391e-005, -4.903215e-005, 
    -2.341816e-005, -8.734314e-006, -8.47131e-006, -1.824759e-005, 
    -1.499429e-005, -5.694976e-006, -8.515393e-006, -9.747595e-006, 
    -5.881735e-006, -7.882341e-006, -7.102513e-006, -1.599838e-005, 
    -1.160018e-005, -5.362555e-006, -3.302346e-006, -5.787238e-006, 
    -5.979211e-006, -1.160055e-005, -6.076436e-006, -9.662777e-006, 
    -1.028665e-005, -8.019924e-006,
  -3.037356e-006, 5.918264e-007, 2.353016e-006, 4.700076e-006, 2.529599e-006, 
    5.270049e-007, -7.009756e-006, -9.668249e-006, -1.698791e-007, 
    -1.126553e-005, -1.065197e-005, -3.893549e-006, 5.606562e-007, 
    7.400922e-008, 7.265558e-007, -1.698731e-007, 4.22063e-006, 
    1.256578e-005, 1.286144e-005, 1.882314e-005, 2.327722e-005, 
    3.598059e-005, 4.886103e-005, 4.156717e-005, 1.630547e-005, 
    1.509239e-005, -3.904235e-006, -8.864947e-006, -6.975857e-006, 
    2.447487e-007, 1.73416e-005, -4.2381e-007, -1.486093e-005, 3.468616e-006, 
    6.548071e-006, -7.484603e-006, 6.176037e-006, -1.128639e-006, 
    -1.763794e-006, -6.332244e-006, 1.637551e-005, 2.269869e-005, 
    1.811261e-005, 2.648769e-005, 1.651557e-005, 4.141279e-006, 
    1.091015e-006, 1.062428e-005, 1.206212e-005, 7.748233e-006, 
    8.665276e-006, 7.135419e-006, 9.822543e-008, -2.463639e-007, 
    -1.587345e-006, 2.571687e-007, 1.21606e-006, -9.831056e-007, 
    1.541277e-006, 8.760617e-007, 5.070142e-007, 2.520534e-006, 
    2.818815e-007, -2.373876e-006, -2.287954e-006, -5.720183e-006, 
    -8.639196e-006, -1.366423e-005, -2.607852e-005, -2.187912e-005, 
    -3.515545e-005, -2.648694e-005, -2.343841e-005, -2.215008e-005, 
    -1.176186e-005, -9.010608e-006, -4.594525e-006, -6.67125e-006, 
    -7.965665e-006, -9.478877e-006, -1.078757e-005, -7.057935e-006, 
    -5.730242e-006, -5.695099e-006, -4.324815e-006, -4.443775e-006, 
    -1.961489e-006, -2.277518e-006, -2.240142e-006, -1.99005e-006, 
    -3.992642e-006, -7.7681e-006, -8.604549e-006, -1.179129e-005, 
    -7.039682e-006, 1.143788e-006,
  -1.898159e-006, -4.4136e-006, 2.780307e-007, 2.963344e-006, 5.142515e-006, 
    3.279621e-006, 1.854449e-006, 4.017353e-006, 5.451093e-006, 
    2.458319e-006, 9.629875e-007, 8.54209e-007, 8.965526e-008, 1.36507e-006, 
    1.315773e-006, -1.716366e-006, -1.924361e-006, 1.553198e-006, 
    5.837777e-006, 1.700918e-005, 1.598944e-005, 4.032229e-005, 
    4.500635e-005, 5.794936e-006, -2.192712e-006, -3.882e-006, 
    -3.751113e-006, -7.160626e-006, -4.058085e-006, 1.164874e-005, 
    2.390399e-006, -8.533651e-006, -2.274712e-005, -2.54115e-006, 
    4.237772e-006, -1.853332e-006, -6.255257e-006, -5.307542e-006, 
    -7.947529e-006, -1.340471e-005, 1.423595e-005, 1.345836e-005, 
    8.958705e-006, 4.623587e-006, 3.718582e-006, 7.494018e-007, 
    6.378068e-006, 1.198352e-005, 8.149196e-006, -9.985015e-007, 
    -2.405544e-006, -3.639732e-006, -4.273157e-006, -5.872424e-006, 
    -4.313515e-006, -1.806889e-006, -1.83247e-006, -1.436472e-006, 
    -2.75535e-006, -3.087272e-006, -1.5265e-006, -2.305458e-006, 
    -6.256501e-006, -3.748635e-006, -1.023039e-005, -1.243005e-005, 
    -1.430127e-005, -6.128103e-007, 6.693976e-006, -3.70232e-006, 
    -2.483465e-005, -2.153702e-005, -1.450479e-005, -1.899749e-005, 
    -1.210086e-005, -1.187362e-005, -1.063744e-005, -7.238115e-006, 
    -9.156887e-006, -6.01982e-006, -3.575533e-006, -1.078968e-006, 
    -1.689792e-006, -5.317233e-007, -1.628325e-006, -1.158193e-006, 
    -2.098704e-006, -1.718477e-006, -1.647075e-006, -1.047924e-006, 
    -7.676581e-007, 3.659477e-007, -3.169601e-006, -9.550154e-006, 
    -9.811669e-006, 5.324655e-007,
  -6.21254e-007, -3.632158e-007, -5.080054e-007, -1.750885e-008, 
    -9.573995e-008, 7.351235e-008, 1.004587e-007, 1.014893e-006, 
    1.466895e-006, 2.544622e-006, 4.417325e-006, 2.276152e-007, 
    2.694626e-007, 2.462541e-006, 7.047504e-006, 2.419328e-006, 
    -1.027684e-006, -1.266226e-006, 6.99299e-006, 2.802027e-005, 
    3.770118e-005, 3.629451e-005, 1.734135e-005, -6.413837e-006, 
    -1.197059e-005, -9.309879e-006, -2.694127e-006, 8.38314e-007, 
    7.330163e-007, 2.150977e-006, 1.586923e-005, 1.22608e-005, 
    -1.056529e-005, -2.577492e-005, -1.152953e-005, -9.053576e-006, 
    -1.406433e-005, -1.706158e-005, -2.114971e-005, -1.843022e-006, 
    4.747635e-006, 2.976754e-006, 7.326773e-006, 8.160372e-006, 
    8.328505e-006, 8.333594e-006, 5.575272e-006, -4.467438e-009, 
    -1.897417e-006, -5.369136e-006, -6.291766e-006, -2.486135e-006, 
    -2.668425e-006, -2.538536e-006, -1.333405e-006, 6.581286e-008, 
    4.090371e-007, 7.711351e-007, -5.873535e-007, -3.018728e-006, 
    -1.714503e-006, -2.608572e-006, -8.19191e-007, -9.641053e-007, 
    -2.446522e-006, -6.079177e-006, -1.871052e-005, -1.960769e-005, 
    -8.477888e-006, -9.544812e-006, -1.135059e-005, -7.523348e-006, 
    -1.123175e-006, -1.518329e-005, -2.168628e-005, -1.556836e-005, 
    -1.306323e-005, -8.350735e-006, -6.198634e-006, -3.123656e-006, 
    -2.764165e-006, -1.860658e-006, -1.969933e-006, -1.574059e-006, 
    -1.290192e-006, -1.619384e-006, -2.438326e-006, -1.566112e-006, 
    -1.786401e-006, -8.142242e-007, -3.038597e-007, -5.053977e-008, 
    -1.565491e-006, -6.71198e-006, -7.736807e-006, -2.356991e-006,
  -2.323339e-007, -6.530435e-007, -9.726733e-007, -8.319816e-008, 
    -5.352e-008, -5.786617e-008, -5.960466e-009, 2.495944e-008, 
    1.115104e-007, -2.364318e-007, 3.129242e-008, 9.92169e-008, 
    9.189051e-009, 1.230836e-006, 5.436937e-006, 1.166475e-005, 
    1.730944e-005, 7.591148e-006, 1.086431e-005, 2.12241e-005, 2.262046e-005, 
    1.230961e-006, -2.363697e-006, 5.506474e-006, 7.382412e-006, 
    8.149938e-006, 3.490848e-006, -1.127062e-005, -2.505505e-006, 
    5.649901e-006, 3.812711e-006, -2.612916e-006, 1.999215e-007, 
    -1.626338e-005, -2.098642e-005, -1.817247e-005, -1.094105e-005, 
    -2.04208e-005, -1.913719e-005, -5.733345e-006, -8.750088e-006, 
    4.246249e-008, 2.913424e-006, 5.36094e-006, 3.805759e-006, 6.719554e-006, 
    4.416332e-006, -3.82488e-006, -8.320807e-006, -7.395944e-006, 
    -8.110579e-006, -4.627307e-006, -4.933774e-006, -1.591925e-007, 
    9.752803e-007, -1.114357e-006, -7.337585e-007, -6.693108e-007, 
    -4.9149e-007, -1.566236e-006, -1.890088e-006, -9.319438e-007, 
    3.227342e-007, 8.710967e-007, -1.601254e-006, -1.663466e-006, 
    -2.36022e-006, -1.664534e-005, -1.605662e-005, 4.975125e-006, 
    6.818151e-006, -6.981441e-006, -1.387052e-007, -3.162771e-006, 
    -3.537782e-006, -2.530589e-006, -1.705313e-006, -6.06602e-007, 
    -2.242004e-006, -3.111983e-006, -1.927838e-006, -1.342347e-006, 
    -5.191814e-007, -9.089708e-007, -1.031781e-006, -7.769713e-007, 
    -9.077294e-007, -1.475463e-006, -1.680851e-006, -8.708485e-007, 
    -6.28705e-007, -3.171464e-007, -7.273009e-007, -1.725554e-006, 
    -2.221391e-006, -1.635651e-006,
  -1.354391e-006, -4.097819e-007, -6.392598e-007, -1.497567e-007, 
    -2.200405e-007, -1.820425e-007, -6.382664e-008, -2.247592e-008, 
    5.215406e-008, -7.45058e-009, -1.158565e-007, -4.594519e-009, 
    6.581345e-009, -7.450573e-010, 7.649263e-007, 3.055731e-006, 
    4.105394e-006, 5.430728e-006, 1.920648e-005, 1.913719e-005, 
    1.432536e-005, 5.791833e-006, 1.143329e-005, 1.545735e-005, 
    1.059982e-005, 3.917603e-005, 4.544643e-005, 6.579859e-006, 
    -3.703681e-006, 6.013361e-006, 5.278362e-006, -6.92904e-007, 
    -3.172718e-007, -5.540751e-007, -2.000245e-005, -1.699763e-005, 
    -1.313412e-006, -1.837798e-007, -3.092115e-006, -1.439221e-007, 
    -2.664452e-006, 5.507245e-007, -1.668432e-006, -7.042414e-006, 
    2.63999e-006, -1.908964e-006, -1.738594e-006, -7.522602e-006, 
    -7.73805e-006, -5.385156e-006, -3.969048e-006, -2.939876e-006, 
    -1.060218e-006, 1.214568e-006, 5.334623e-007, -1.467761e-007, 
    2.420193e-007, -4.095327e-007, -1.389782e-006, -1.460437e-006, 
    -1.189982e-006, 9.81117e-007, 1.448765e-006, 2.856054e-007, 
    1.135468e-006, -4.508843e-007, -1.361842e-006, -6.420041e-006, 
    3.919013e-007, 1.025337e-005, 7.980068e-006, 1.828248e-006, 
    7.276114e-006, 7.179877e-006, 8.861207e-007, -4.292029e-006, 
    -4.112349e-006, -2.836559e-006, -4.610916e-006, -3.151719e-006, 
    -1.612306e-006, -2.846991e-006, -1.516938e-006, -2.801416e-007, 
    3.32172e-007, -9.67706e-007, -1.119201e-006, -1.01539e-006, 
    -1.557668e-006, -1.516566e-006, -1.445909e-006, -1.001483e-006, 
    -6.916623e-007, -4.708767e-007, -1.262377e-006, -2.969553e-006,
  -3.753727e-006, -2.793223e-006, -1.485273e-006, -6.773819e-007, 
    -5.30233e-007, -7.373591e-007, -4.107754e-007, -1.600633e-007, 
    -1.621743e-007, -2.682208e-008, -2.304713e-007, -3.588696e-008, 
    3.513995e-023, -5.438924e-008, 6.10948e-008, 3.131727e-007, 
    1.216928e-008, 5.81642e-007, 7.578235e-006, 9.55537e-006, 9.336199e-006, 
    2.034604e-005, 3.858902e-006, 2.649178e-006, -4.628298e-006, 
    -1.404936e-006, 9.184208e-006, -7.89389e-006, -6.841583e-008, 
    1.092081e-005, 1.381983e-005, 1.968741e-005, 1.667875e-005, 
    1.242259e-006, -7.189563e-006, -7.232527e-006, -3.295645e-007, 
    5.271037e-006, 4.259346e-008, -4.04194e-007, 1.253064e-006, 
    5.056463e-007, 1.000844e-007, -2.702573e-006, -7.5549e-007, 1.71351e-006, 
    -1.795597e-007, -1.202277e-006, -3.313274e-006, -5.673368e-006, 
    -2.034257e-006, 8.910893e-007, 1.181787e-006, 1.256043e-006, 
    -1.824155e-007, -1.572071e-007, -2.756715e-007, -4.718704e-007, 
    -1.02967e-006, -1.750514e-006, -8.83887e-007, 2.732122e-009, 
    2.30968e-007, 1.599888e-006, 6.439786e-007, 1.632918e-007, 
    -4.000963e-007, 6.424889e-007, 7.779399e-006, 5.477295e-006, 
    2.532576e-006, 1.805648e-006, 8.195457e-009, -1.057113e-006, 
    -3.872065e-006, -4.416208e-006, -8.388732e-006, -1.136686e-005, 
    -1.004152e-005, -7.459521e-006, -7.335594e-006, -6.497278e-006, 
    -2.794091e-006, -1.603861e-006, -8.30616e-007, 3.216164e-007, 
    -4.544836e-008, -7.592143e-007, -1.657754e-007, -8.848806e-007, 
    -9.384007e-007, -1.074746e-006, 3.762543e-007, -4.801899e-007, 
    -4.777064e-007, -5.117183e-006,
  -4.896522e-006, -5.71236e-006, -4.640221e-006, -4.301469e-006, 
    -1.352653e-006, -4.785757e-007, -1.074498e-006, -7.249415e-007, 
    -1.046807e-006, -1.001979e-006, -1.470248e-007, -1.054257e-007, 
    -1.90859e-007, -1.239528e-006, -4.562239e-007, 3.72529e-009, 
    8.195641e-009, 2.508362e-008, -6.300708e-007, -1.193335e-006, 
    1.072139e-006, 4.593285e-007, 2.210254e-008, 1.340483e-006, 
    1.399219e-006, -2.345692e-006, 5.891423e-006, 3.122985e-005, 
    2.312585e-005, 1.384156e-005, 2.246226e-005, 2.58421e-005, 2.213021e-005, 
    1.395084e-005, 7.189312e-006, 4.275764e-006, 5.271162e-006, 
    1.745546e-006, 2.335757e-006, 3.861513e-006, 5.915139e-006, 
    1.142509e-005, 9.591504e-006, 7.959081e-006, 6.347647e-006, 
    4.923097e-006, 5.845601e-006, 4.056593e-006, 1.596163e-006, 
    -1.319374e-006, -1.708294e-006, -2.241507e-006, -7.988265e-007, 
    1.672159e-006, 4.235653e-007, -1.074622e-006, -6.036207e-007, 
    -1.291806e-006, -5.858637e-007, -1.061212e-006, -1.080955e-006, 
    -5.067636e-007, 1.755853e-007, 2.864748e-007, 4.579624e-007, 
    8.350859e-007, 4.677722e-007, 1.33241e-007, 2.603481e-006, 4.389759e-006, 
    2.249952e-006, -1.675635e-006, -2.034381e-006, -6.051123e-007, 
    5.304792e-007, 3.30657e-006, 8.484225e-006, 2.754728e-006, 
    -2.191089e-006, -7.38067e-006, -1.052631e-005, -8.066247e-006, 
    -7.330377e-006, -7.462751e-006, -4.053861e-006, -2.231822e-006, 
    -1.157696e-006, -1.073877e-006, -3.409882e-007, -1.017377e-006, 
    -6.059781e-008, -8.997815e-007, -6.244827e-007, 5.004308e-007, 
    -5.369385e-007, -1.216431e-006,
  -3.937508e-006, -2.370154e-006, -2.608821e-006, -2.923111e-006, 
    -3.048281e-006, -2.172838e-006, -1.747285e-006, -1.962483e-006, 
    -3.516177e-006, -3.027419e-006, -1.359483e-006, -2.135957e-006, 
    -1.832222e-006, -1.62373e-006, -1.212955e-006, -8.087604e-007, 
    -4.060564e-008, 2.793968e-008, 1.676381e-008, -1.723443e-006, 
    -4.506608e-006, -5.061429e-007, -3.041077e-007, 4.502635e-007, 
    -1.076982e-006, -1.204535e-008, -3.353132e-006, -7.421477e-010, 
    1.413177e-005, 1.623097e-005, 1.491085e-005, 1.622624e-005, 
    2.339694e-005, 3.489827e-005, 2.88335e-005, 1.256131e-005, 1.090491e-005, 
    1.854189e-005, 1.078633e-005, 7.07768e-006, 5.912036e-006, 5.746137e-006, 
    5.129848e-006, 6.305676e-006, 8.352723e-006, 1.047763e-005, 
    9.103618e-006, 6.989889e-006, 8.919833e-006, 6.114815e-006, 
    2.316387e-006, 1.223634e-006, -2.061326e-006, 7.947347e-008, 
    1.977011e-006, 1.190728e-006, 3.890445e-007, -4.96706e-007, 
    -7.104131e-007, -5.303573e-007, -7.692724e-007, -7.883955e-007, 
    -5.938111e-007, -2.643714e-007, 3.748885e-007, 1.049538e-006, 
    1.318753e-006, 1.170238e-006, 4.96432e-006, 7.482864e-006, 4.646681e-007, 
    -4.477923e-006, -4.899997e-006, -4.510075e-007, 3.098943e-006, 
    2.421562e-006, 2.489116e-006, 4.807487e-006, -9.562827e-007, 
    -4.825368e-006, -4.671641e-006, -7.302064e-006, -6.078431e-006, 
    -5.615006e-006, -7.265186e-006, -7.09109e-006, -3.28198e-006, 
    -1.787394e-006, -1.015266e-006, -1.376495e-006, -8.319817e-007, 
    -1.289323e-006, -1.443799e-006, -1.370037e-006, -1.658624e-006, 
    -3.136943e-006,
  -5.95438e-006, -2.41821e-006, -3.53468e-006, -4.704173e-006, 
    -3.676862e-006, -4.710008e-006, -4.991516e-006, -3.570567e-006, 
    -3.566841e-006, -2.060583e-006, -2.027552e-006, -5.41235e-006, 
    -5.842497e-006, -1.649931e-006, -7.50646e-007, -5.301088e-007, 
    3.36518e-007, 4.823009e-007, 2.243867e-007, 4.029522e-007, 
    -1.994272e-007, -8.543334e-007, -3.481905e-007, -1.228601e-006, 
    -5.323441e-007, -9.320675e-007, -5.242719e-007, -4.127745e-006, 
    -4.707401e-006, -2.767765e-006, -2.197921e-007, 6.826471e-006, 
    1.515547e-005, 1.561282e-005, 2.583476e-005, 2.343705e-005, 
    1.755779e-005, 1.141143e-005, 6.420538e-006, 6.026028e-006, 
    5.451344e-006, 2.178178e-006, -3.640853e-007, -4.280606e-006, 
    3.13409e-006, 8.75791e-006, 4.624202e-006, 2.944966e-006, 5.596008e-006, 
    5.282713e-006, 4.52002e-006, 6.160262e-006, 2.472101e-006, 3.334755e-006, 
    3.299614e-006, 2.703319e-006, 1.122306e-006, -1.480184e-007, 
    -1.682341e-006, -1.220405e-006, -1.429518e-006, -1.244868e-006, 
    -1.181414e-006, -1.956398e-006, -2.138441e-006, 3.757577e-007, 
    1.610443e-006, 5.011012e-006, 1.10019e-005, 1.124106e-005, 4.054731e-006, 
    -4.166141e-007, 2.103425e-006, 5.049005e-007, -5.152087e-007, 
    4.229441e-007, -2.128381e-006, -2.386545e-006, -5.342935e-006, 
    -8.299946e-006, -1.035631e-005, -1.056405e-005, -8.608898e-006, 
    -6.999077e-006, -5.517528e-006, -4.214048e-006, -3.860146e-006, 
    -4.129608e-006, -2.948444e-006, -1.206249e-006, -1.553322e-006, 
    -1.407042e-006, -1.437217e-006, -3.560508e-006, -2.766276e-006, 
    -5.026783e-006,
  -6.659702e-006, -7.117167e-006, -1.105877e-005, -1.021015e-005, 
    -2.68879e-006, -2.622108e-006, -2.607332e-006, -3.418078e-006, 
    -3.134955e-006, -2.866611e-006, -2.101809e-006, -4.077951e-006, 
    -6.285683e-006, -4.757196e-006, -3.368905e-007, 1.647075e-006, 
    9.218852e-007, 9.69693e-007, 5.698453e-007, 1.147389e-007, 
    -1.023213e-007, 4.343688e-007, -1.323715e-007, 6.52919e-007, 
    1.266722e-006, 2.567967e-007, 1.611559e-006, 3.289182e-006, 3.12974e-006, 
    1.022843e-006, 4.253165e-006, 8.177882e-006, 6.720053e-006, 
    9.435043e-006, 1.202735e-005, 1.308161e-005, 1.329357e-005, 
    1.455732e-005, 9.923551e-006, 6.028265e-006, 7.183105e-006, 
    3.275276e-006, 2.19221e-006, 3.291898e-007, -1.403816e-006, 
    1.016135e-006, 5.915263e-006, 4.547463e-006, 1.532957e-006, 
    -8.854113e-008, 2.685956e-007, 1.205379e-006, 1.709537e-006, 
    3.727029e-006, 1.142669e-006, 1.509612e-006, 2.021343e-006, 
    4.903713e-007, -2.265722e-006, -2.057353e-006, -1.6508e-006, 
    -1.593555e-006, -3.520399e-006, -3.686423e-006, -4.508471e-006, 
    -3.415595e-006, 7.84421e-007, 8.040442e-007, 5.003094e-007, 
    6.406877e-006, 6.493801e-006, 3.512203e-006, -8.925799e-007, 
    -3.331403e-006, -3.181151e-006, -1.840419e-006, 3.273271e-007, 
    4.554822e-007, -3.848218e-007, -4.600486e-006, -1.007827e-005, 
    -1.019215e-005, -5.449605e-006, -4.316866e-006, -4.408881e-006, 
    -3.036361e-006, -1.990546e-006, -6.438549e-007, -1.371403e-006, 
    -1.433493e-006, -2.46639e-006, -2.238651e-006, -2.595659e-006, 
    -3.438195e-006, -4.532809e-006, -6.702543e-006,
  -7.390356e-006, -8.455665e-006, -6.114817e-006, -3.651778e-006, 
    2.210345e-007, 2.430503e-006, 2.252187e-006, -1.978999e-006, 
    -2.468998e-006, -4.121663e-006, -7.29784e-007, 1.794596e-006, 
    6.64344e-007, -3.206233e-007, -7.209683e-007, -9.605037e-007, 
    8.881088e-007, 1.194328e-006, 2.063935e-006, 2.460431e-006, 
    3.020838e-006, 2.267709e-006, 1.96062e-006, 1.519795e-006, 6.432329e-007, 
    -4.405774e-007, 2.153465e-006, 1.568347e-006, 3.65451e-006, 
    6.920098e-006, 7.111828e-006, 5.814432e-006, 6.303937e-006, 
    6.107737e-006, 5.880742e-006, 1.19716e-005, 1.090467e-005, 7.743762e-006, 
    4.268933e-006, 1.088407e-006, 3.52909e-006, 5.332753e-006, 6.896877e-006, 
    5.120659e-006, 2.892191e-006, -1.985703e-006, -2.78217e-006, 
    1.02495e-006, 9.17913e-007, 5.811307e-008, -5.270049e-007, 
    -1.145028e-006, -1.718479e-006, 2.4536e-006, 5.803009e-006, 
    5.779539e-006, 2.393499e-006, -1.599765e-006, -1.255052e-006, 
    -9.554133e-007, -1.523395e-006, -2.157812e-006, -2.938012e-006, 
    -1.643721e-006, -3.287321e-006, -4.491085e-006, -6.722912e-007, 
    4.168596e-007, 7.054459e-007, 1.094366e-006, -8.778006e-007, 
    -1.953791e-006, 4.113936e-007, 2.303495e-007, -1.187498e-006, 
    -2.611428e-006, -1.22028e-006, 3.597379e-007, 5.110229e-006, 
    7.513041e-006, 1.722448e-006, -9.155519e-007, -6.036087e-006, 
    -7.311253e-006, -5.197155e-006, -2.006815e-006, 1.707052e-006, 
    7.901326e-007, 8.20557e-007, 3.909081e-007, -2.024197e-006, 
    -3.286699e-006, -2.247842e-006, -3.144765e-006, -4.758438e-006, 
    -6.436432e-006,
  -6.162863e-007, -1.007815e-006, -1.53954e-006, -2.631545e-006, 
    -2.104043e-006, -2.715737e-006, -1.971175e-006, 6.409973e-007, 
    1.640494e-006, 1.037493e-006, -1.852713e-007, -3.657005e-007, 
    1.337503e-006, 3.316998e-006, 3.764281e-006, 3.050887e-006, 
    2.024572e-006, 2.380957e-006, 2.597396e-006, 1.893564e-006, 
    2.839663e-006, 3.309176e-006, 1.179054e-006, 5.255151e-007, 
    2.089888e-006, 4.972269e-006, 7.974977e-006, 7.695333e-006, 
    3.633773e-006, 4.346668e-006, 8.668874e-006, 3.789864e-006, 
    1.355013e-006, 4.378955e-006, 3.133839e-006, 4.805999e-006, 
    7.453313e-006, 4.952029e-006, 3.779929e-006, 4.291534e-006, 
    4.817297e-006, 4.646057e-006, 5.400303e-006, 4.194306e-006, 
    3.117819e-006, 2.416595e-006, 3.316252e-006, 2.058719e-006, 
    6.000209e-007, -4.485246e-007, -2.38071e-006, -3.335372e-007, 
    -5.553156e-007, 5.479906e-007, 3.034249e-006, 3.104906e-006, 
    6.280825e-007, 1.489247e-006, 1.379351e-006, 9.838477e-007, 
    -1.396487e-006, -2.079953e-006, 1.183278e-006, 3.26286e-006, 
    -1.27442e-006, 5.348265e-007, 1.802046e-006, -6.799892e-007, 
    -1.357248e-006, -1.740937e-007, 1.739336e-006, 4.221871e-006, 
    7.439412e-007, -2.90585e-006, -1.961986e-006, -3.157804e-006, 
    -3.562865e-006, -1.98136e-006, 2.487377e-006, 5.183989e-006, 
    6.793685e-006, 3.772104e-006, 1.336761e-006, -5.761794e-007, 
    -3.165129e-006, -1.35017e-006, 2.426779e-006, 5.389873e-006, 
    3.760182e-006, 3.860892e-006, 3.737583e-006, 8.28506e-007, 7.661583e-008, 
    1.39537e-006, 1.529852e-006, -3.745154e-007,
  8.205589e-007, 1.247476e-006, 6.185237e-007, -3.733114e-006, 
    -3.374493e-006, 2.644956e-007, 1.348059e-006, 9.448577e-007, 
    5.816542e-006, 4.365047e-006, 4.562244e-007, 2.003833e-006, 
    4.046784e-006, 3.515433e-006, 3.725663e-006, 5.727137e-006, 6.08849e-006, 
    4.179155e-006, 3.213932e-006, 1.996508e-006, 1.524266e-006, 
    2.209223e-006, 2.854442e-006, 3.33041e-006, 3.775333e-006, 7.699926e-006, 
    6.186094e-006, 4.846353e-006, 2.764536e-006, 2.137323e-006, 
    3.087025e-006, 4.389261e-006, -1.987941e-006, -2.25765e-006, 
    -7.20247e-008, 3.958121e-006, 2.805638e-006, 1.879658e-006, 
    4.649288e-006, 4.819283e-006, 6.091595e-006, 5.239122e-006, 
    4.804382e-006, 5.055716e-006, 4.555408e-006, 2.904486e-006, 
    3.810226e-006, 2.982344e-006, 2.584729e-006, 2.328678e-006, 
    -6.648406e-007, -7.705148e-007, 1.784429e-007, -5.907077e-007, 
    9.238647e-008, 3.57305e-006, 1.972914e-006, -4.611902e-007, 
    -4.075482e-007, 4.979483e-008, 2.829607e-006, 2.38133e-006, 
    1.365443e-006, 4.383674e-006, 2.721821e-006, 2.968435e-006, 
    2.549838e-006, 3.007675e-006, 7.336836e-006, 6.940092e-006, 
    6.016469e-006, 1.609946e-006, -2.036368e-006, -1.169741e-006, 
    1.057735e-006, 1.852835e-006, 3.666679e-006, 8.598468e-006, 
    5.056585e-006, 6.798655e-007, 4.827354e-006, 3.837051e-006, 
    4.139667e-006, 4.752354e-006, 1.652663e-006, -3.977369e-006, 
    -1.395743e-006, 2.100194e-006, 2.840161e-006, 3.91466e-006, 
    2.562256e-006, 5.944312e-007, -1.277029e-006, -8.141014e-007, 
    2.205372e-006, 2.844879e-006,
  3.192948e-006, 1.491854e-006, -2.100567e-006, -5.54472e-006, 
    -5.835667e-006, -1.115974e-006, -2.529468e-007, 1.999251e-008, 
    3.248442e-007, 1.270697e-006, 7.799517e-007, 1.785407e-006, 
    3.692632e-006, 2.867853e-006, 3.879766e-006, 4.939982e-006, 4.48438e-006, 
    2.475703e-006, 2.11969e-006, 2.032146e-006, 3.280118e-006, 3.521145e-006, 
    2.391886e-006, 1.909833e-006, 4.354242e-006, 5.993992e-006, 
    4.564723e-006, 4.448742e-006, 2.405917e-006, 3.064177e-006, 
    3.234918e-006, 1.261134e-006, 1.271565e-007, 2.200033e-006, 
    2.962724e-006, 2.173208e-006, 1.574554e-007, -3.323705e-006, 
    -1.153599e-006, 8.114424e-006, 1.169108e-005, 8.102879e-006, 
    4.191572e-006, 4.098938e-006, 5.733471e-006, 6.202608e-006, 
    6.041922e-006, 4.067893e-006, 1.29131e-006, 1.762055e-007, 3.04728e-007, 
    1.41648e-006, 2.857298e-006, 3.816189e-006, 3.240009e-006, 5.119171e-006, 
    9.569154e-006, 1.319548e-005, 9.140869e-006, 6.613878e-006, 
    4.699083e-006, 1.756103e-006, 4.068512e-006, 7.727494e-006, 7.29064e-006, 
    4.975746e-006, 2.816691e-006, 1.136834e-006, 2.219653e-006, 
    6.363913e-006, 5.441034e-006, 2.982724e-007, 1.179178e-006, 
    2.664576e-006, 2.377976e-006, 2.430626e-006, 3.16538e-006, 5.104144e-006, 
    8.142119e-006, 1.150593e-005, 9.379411e-006, 3.130608e-006, 4.67375e-006, 
    9.116035e-006, 7.152805e-006, 2.279256e-006, -1.428649e-006, 
    -9.119503e-007, 1.367802e-006, 3.797311e-006, 4.376347e-006, 
    2.421562e-006, 1.370287e-006, -3.992263e-007, 1.646455e-006, 2.715116e-006,
  3.061444e-006, 2.710273e-006, 1.133109e-006, -3.465775e-007, 7.495291e-007, 
    1.035623e-007, 4.04194e-007, 1.876057e-006, 1.222515e-006, 1.085922e-006, 
    8.481238e-007, 1.240272e-006, 2.124532e-006, 3.667672e-006, 
    3.335997e-006, 3.325442e-006, 3.972898e-006, 3.342084e-006, 
    3.167241e-006, 2.649054e-006, 3.747393e-006, 4.041567e-006, 
    2.260505e-006, 3.019224e-006, 2.808869e-006, 7.60705e-007, 
    -9.150554e-007, -2.47173e-006, -2.978244e-006, 9.884443e-007, 
    1.384815e-006, -1.006945e-006, 2.654888e-007, 1.16403e-006, 
    -7.19725e-007, -1.218417e-006, 4.759677e-007, 2.169858e-006, 
    1.286468e-006, 4.021203e-006, 6.527951e-006, 6.411473e-006, 
    6.006659e-006, 4.654254e-006, 3.835063e-006, 4.554911e-006, 
    6.374345e-006, 3.501773e-006, -4.917456e-008, 1.560151e-006, 
    1.408782e-006, 2.970301e-007, 2.948071e-006, 5.148971e-006, 
    5.858266e-006, 7.524464e-006, 8.162608e-006, 6.921713e-006, 
    7.228429e-006, 6.797787e-006, 5.334367e-006, 5.77482e-006, 5.803755e-006, 
    4.139047e-006, 2.93168e-006, 3.164385e-006, 1.096229e-006, 
    -1.046557e-006, 3.957502e-007, 2.11882e-006, 2.639492e-006, 
    2.089143e-006, 2.349789e-006, 5.074218e-006, 5.966052e-006, 
    5.448112e-006, 4.431234e-006, 3.191331e-006, 5.172815e-006, 
    6.936118e-006, 7.707129e-006, 5.993868e-006, 6.083399e-006, 
    7.262703e-006, 7.349377e-006, 4.67437e-006, -3.003948e-006, 
    -3.230323e-006, -8.780517e-007, 2.387291e-006, 3.732244e-006, 
    4.677846e-006, 4.289051e-006, 2.914046e-006, 1.758958e-006, 1.959253e-006,
  9.757769e-007, 7.660437e-007, 1.165768e-006, 9.819869e-007, 2.031152e-006, 
    2.286583e-006, 1.485148e-006, 2.051642e-006, 2.855932e-006, 2.27342e-006, 
    9.689484e-007, 2.016623e-007, -6.33424e-007, 9.85091e-007, 3.69884e-006, 
    3.749753e-006, 3.167615e-006, 3.627687e-006, 3.712501e-006, 
    2.302479e-006, 3.085162e-006, 3.92658e-006, 4.140287e-006, 3.50202e-006, 
    2.650047e-006, 2.85022e-006, 2.800549e-006, 1.370037e-006, 
    -3.787318e-008, 5.412858e-007, -5.518395e-007, -1.089398e-006, 
    -5.751863e-007, 2.007946e-007, 2.276898e-006, 7.953495e-007, 
    1.457334e-006, 2.444038e-006, 3.201018e-006, 6.140272e-006, 
    6.177774e-006, 5.110602e-006, 4.831826e-006, 4.644444e-006, 
    3.953527e-006, 3.799672e-006, 4.084782e-006, 2.67153e-006, 4.656489e-006, 
    6.352366e-006, 6.50088e-006, 4.386281e-006, 2.493212e-006, 2.156446e-006, 
    1.409649e-006, 2.543751e-006, 2.755722e-006, 2.669542e-006, 
    1.700719e-006, 2.934783e-006, 5.141771e-006, 5.357092e-006, 
    4.943834e-006, 4.030268e-006, 2.640983e-006, 3.98235e-007, 
    -6.561477e-007, -2.731877e-007, -3.475698e-007, -1.937151e-007, 
    9.387804e-008, 3.640844e-007, 1.913433e-006, 3.033876e-006, 
    2.522518e-006, 1.791244e-006, 1.290565e-006, 2.146016e-006, 
    5.696216e-006, 7.141506e-006, 3.936763e-006, 2.262865e-006, 
    3.174071e-006, 3.43894e-006, 9.461e-007, -1.992781e-006, -2.976507e-006, 
    -1.090642e-006, 1.281871e-006, 1.128888e-006, 2.960115e-006, 
    4.840518e-006, 3.016367e-006, 1.621122e-006, 1.631429e-006, 1.905238e-006,
  1.057734e-006, 3.116747e-008, -3.964951e-007, 8.82892e-008, 1.113365e-006, 
    2.526988e-006, 2.931928e-006, 2.77621e-006, 3.328299e-006, 2.98818e-006, 
    2.659609e-006, 1.814713e-006, 1.519049e-006, 2.055491e-006, 
    2.793719e-006, 3.318736e-006, 2.666315e-006, 1.299257e-006, 
    2.977749e-007, 1.004339e-006, 2.151107e-006, 2.429634e-006, 
    2.689288e-006, 3.278753e-006, 3.228709e-006, 2.234801e-006, 
    1.245613e-006, 2.183766e-006, 3.081808e-006, 8.682418e-007, 
    -3.190089e-007, 2.63627e-007, 1.050532e-006, 1.443425e-006, 
    1.506135e-006, 1.688798e-006, 1.343712e-006, -3.849436e-008, 
    -1.055872e-006, -5.601596e-007, -2.168126e-007, -4.7311e-008, 
    1.17744e-006, 1.652911e-006, 4.988169e-007, 4.912417e-007, 1.783793e-006, 
    2.679229e-006, 3.227716e-006, 3.218278e-006, 3.138309e-006, 
    2.863507e-006, 2.072751e-006, 2.354508e-006, 2.667432e-006, 
    1.936158e-006, 9.268524e-007, 7.571034e-007, 8.835141e-007, 1.47832e-006, 
    2.184014e-006, 2.6195e-006, 3.177548e-006, 3.390014e-006, 2.697731e-006, 
    2.127762e-006, 1.15186e-006, 4.888825e-007, 1.09151e-006, 1.168872e-006, 
    1.38407e-006, 1.905858e-006, 3.163765e-006, 2.748271e-006, 2.352272e-006, 
    3.556286e-006, 4.080559e-006, 2.236167e-006, 2.715737e-006, 
    3.620734e-006, 2.982468e-006, 2.504016e-006, 2.854317e-006, 
    1.936158e-006, 1.247724e-006, 1.420826e-006, 2.252063e-006, 
    2.473593e-006, 2.262369e-006, 2.591685e-006, 4.136065e-006, 
    3.928692e-006, 3.160784e-006, 3.377099e-006, 3.213932e-006, 1.867115e-006,
  1.224876e-006, 1.348679e-006, 1.693766e-006, 1.341974e-006, 7.984536e-007, 
    8.761881e-007, 7.131448e-007, 4.313888e-007, 3.743917e-007, 
    7.811932e-007, 1.48813e-006, 1.498561e-006, 1.191472e-006, 9.996193e-007, 
    8.24034e-007, 9.017685e-007, 7.003546e-007, 3.065907e-007, 2.041461e-007, 
    -2.468632e-007, -6.314367e-007, -1.35351e-008, 1.021102e-006, 
    1.510854e-006, 1.750762e-006, 1.240273e-006, 1.678864e-007, 
    -5.389256e-007, -3.483146e-007, 1.600629e-007, 1.815461e-007, 
    3.961222e-007, 7.264316e-007, 1.127024e-006, 1.549721e-006, 1.93566e-006, 
    1.498808e-006, 8.142242e-007, 7.305298e-007, 1.447524e-006, 
    1.939635e-006, 2.20413e-006, 2.722442e-006, 3.002212e-006, 2.742931e-006, 
    2.420196e-006, 1.878664e-006, 1.482417e-006, 1.180296e-006, 
    1.050532e-006, 9.992473e-007, 4.816793e-007, 2.863508e-007, 
    5.315987e-007, 8.447714e-007, 9.379037e-007, 9.971359e-007, 
    8.682405e-007, 9.793794e-007, 1.306335e-006, 1.703327e-006, 
    1.914675e-006, 2.017617e-006, 1.800681e-006, 1.541277e-006, 1.51222e-006, 
    1.204014e-006, 1.600882e-006, 2.326941e-006, 2.779439e-006, 
    3.185247e-006, 3.23976e-006, 2.938261e-006, 1.991664e-006, 1.424427e-006, 
    1.432747e-006, 1.554812e-006, 1.46913e-006, 2.183765e-006, 2.851958e-006, 
    3.231565e-006, 2.881885e-006, 2.027055e-006, 1.236052e-006, 
    5.899619e-007, 5.702179e-007, 1.539414e-006, 2.376735e-006, 
    2.751251e-006, 2.984454e-006, 3.054117e-006, 2.856428e-006, 
    2.585228e-006, 2.454346e-006, 2.356371e-006, 1.833837e-006,
  1.686439e-006, 1.503652e-006, 1.302858e-006, 8.615357e-007, 7.960948e-007, 
    6.544092e-007, 3.241003e-007, 2.759198e-007, 6.047389e-007, 
    1.189361e-006, 1.747037e-006, 2.091254e-006, 1.802295e-006, 
    1.138076e-006, 6.966293e-007, 7.782128e-007, 1.139442e-006, 
    1.344705e-006, 1.233071e-006, 1.247351e-006, 1.286716e-006, 
    1.203393e-006, 1.045813e-006, 1.028056e-006, 9.602554e-007, 7.55861e-007, 
    6.649643e-007, 5.880993e-007, 4.661579e-007, 2.067536e-007, 
    -1.482667e-007, -4.58459e-007, -8.220477e-007, -1.015142e-006, 
    -8.286288e-007, -4.860267e-007, 1.138696e-007, 9.206433e-007, 
    1.462673e-006, 1.776591e-006, 2.106776e-006, 2.227724e-006, 
    2.205745e-006, 2.160668e-006, 1.98707e-006, 1.453732e-006, 8.6613e-007, 
    6.182736e-007, 5.746879e-007, 5.080055e-007, 3.819659e-007, 
    2.242623e-007, 4.275389e-007, 7.708868e-007, 8.56568e-007, 1.112496e-006, 
    1.413127e-006, 1.594176e-006, 1.692027e-006, 1.566608e-006, 
    1.128515e-006, 7.309022e-007, 5.818902e-007, 8.292495e-007, 1.16676e-006, 
    1.280134e-006, 1.323099e-006, 1.38916e-006, 1.26784e-006, 6.87688e-007, 
    1.644094e-007, -3.663263e-008, 1.671415e-007, 3.858158e-007, 
    4.481522e-007, 6.95512e-007, 8.365764e-007, 1.030539e-006, 1.02073e-006, 
    7.091712e-007, 4.547333e-007, 6.895511e-007, 8.49242e-007, 7.472931e-007, 
    6.700554e-007, 5.73074e-007, 6.311886e-007, 9.694447e-007, 1.459196e-006, 
    1.700719e-006, 1.722078e-006, 1.554067e-006, 1.279016e-006, 
    1.153971e-006, 1.411016e-006, 1.710653e-006,
  -5.319716e-007, -7.444369e-007, -8.637708e-007, -7.809454e-007, 
    -4.620601e-007, -3.588684e-008, 3.310543e-007, 5.48735e-007, 6.3777e-007, 
    7.539984e-007, 8.939455e-007, 9.96391e-007, 9.899336e-007, 8.537122e-007, 
    7.409603e-007, 7.312747e-007, 7.32889e-007, 7.731219e-007, 8.987886e-007, 
    1.090889e-006, 1.297146e-006, 1.376743e-006, 1.253933e-006, 
    9.699415e-007, 5.756815e-007, 1.656513e-007, -1.0853e-007, 
    -7.313974e-008, 1.157323e-007, 3.3987e-007, 4.266703e-007, 3.527848e-007, 
    2.556799e-007, 1.435483e-007, 1.103936e-007, 2.841152e-007, 
    6.294495e-007, 9.616215e-007, 1.111627e-006, 1.155709e-006, 
    1.228725e-006, 1.375998e-006, 1.519918e-006, 1.675263e-006, 
    1.842032e-006, 1.911447e-006, 1.850227e-006, 1.655022e-006, 
    1.354515e-006, 1.007194e-006, 7.019694e-007, 4.990652e-007, 
    4.287808e-007, 4.307676e-007, 4.054359e-007, 3.301843e-007, 
    3.320474e-007, 4.338722e-007, 6.788719e-007, 1.027932e-006, 1.24375e-006, 
    1.239529e-006, 1.164649e-006, 1.119822e-006, 1.198178e-006, 
    1.320988e-006, 1.349673e-006, 1.319746e-006, 1.273429e-006, 
    1.277029e-006, 1.344209e-006, 1.353522e-006, 1.225249e-006, 
    1.060342e-006, 9.670853e-007, 9.583928e-007, 8.955599e-007, 
    7.310259e-007, 4.842877e-007, 2.899519e-007, 1.763306e-007, 
    8.630241e-008, -8.195457e-009, -1.055514e-008, 9.77268e-008, 
    1.485148e-007, 9.052451e-008, -2.781553e-008, -9.909309e-008, 
    -4.569711e-008, 5.240236e-008, 1.738499e-009, -1.524886e-007, 
    -2.606462e-007, -2.98644e-007, -3.756331e-007,
  -8.821485e-007, -9.155519e-007, -9.454784e-007, -9.575238e-007, 
    -9.361652e-007, -8.794168e-007, -7.866574e-007, -6.678206e-007, 
    -5.407883e-007, -4.138797e-007, -2.976508e-007, -1.899898e-007, 
    -8.493635e-008, 1.105172e-008, 8.679899e-008, 1.283984e-007, 
    1.353524e-007, 1.121311e-007, 6.755181e-008, 2.930528e-008, 
    1.465241e-008, 3.352761e-008, 9.425003e-008, 1.892445e-007, 
    3.077089e-007, 4.333751e-007, 5.621459e-007, 6.812315e-007, 
    7.951012e-007, 9.077285e-007, 1.010299e-006, 1.103307e-006, 
    1.186132e-006, 1.259769e-006, 1.326327e-006, 1.381338e-006, 
    1.422316e-006, 1.446158e-006, 1.445164e-006, 1.42095e-006, 1.382704e-006, 
    1.336634e-006, 1.283363e-006, 1.230464e-006, 1.184146e-006, 
    1.148631e-006, 1.118829e-006, 1.093497e-006, 1.06978e-006, 1.049911e-006, 
    1.022344e-006, 9.863325e-007, 9.561577e-007, 9.495766e-007, 
    9.808691e-007, 1.045441e-006, 1.133357e-006, 1.232699e-006, 
    1.325831e-006, 1.397356e-006, 1.425668e-006, 1.391521e-006, 
    1.281996e-006, 1.115724e-006, 9.049973e-007, 6.639712e-007, 4.02456e-007, 
    1.404433e-007, -1.170984e-007, -3.628438e-007, -5.746883e-007, 
    -7.294116e-007, -8.324787e-007, -8.861221e-007, -8.87364e-007, 
    -8.497386e-007, -7.790827e-007, -6.817281e-007, -5.638844e-007, 
    -4.378458e-007, -3.1131e-007, -1.95826e-007, -9.611222e-008, 
    -3.216155e-008, -7.823019e-009, -2.793968e-008, -8.49368e-008, 
    -1.703702e-007, -2.667311e-007, -3.560135e-007, -4.379699e-007, 
    -5.230308e-007, -6.187706e-007, -7.152557e-007, -7.947287e-007, 
    -8.476277e-007,
  3.599872e-007, 3.23852e-007, 2.902001e-007, 2.638747e-007, 2.437581e-007, 
    2.328306e-007, 2.278636e-007, 2.277394e-007, 2.314647e-007, 2.39412e-007, 
    2.503394e-007, 2.65489e-007, 2.829979e-007, 3.00631e-007, 3.155321e-007, 
    3.254663e-007, 3.283222e-007, 3.234794e-007, 3.124277e-007, 
    2.970298e-007, 2.805144e-007, 2.661099e-007, 2.517055e-007, 
    2.409021e-007, 2.355625e-007, 2.322098e-007, 2.346933e-007, 
    2.432614e-007, 2.572933e-007, 2.769133e-007, 2.987683e-007, 
    3.229827e-007, 3.434718e-007, 3.59118e-007, 3.748884e-007, 3.905346e-007, 
    4.044424e-007, 4.21082e-007, 4.392117e-007, 4.593284e-007, 4.821767e-007, 
    5.053977e-007, 5.226583e-007, 5.312264e-007, 5.284945e-007, 
    5.099922e-007, 4.788241e-007, 4.397083e-007, 3.952533e-007, 
    3.509224e-007, 3.142903e-007, 2.839913e-007, 2.617637e-007, 
    2.443792e-007, 2.336997e-007, 2.31589e-007, 2.360591e-007, 2.45745e-007, 
    2.620122e-007, 2.82377e-007, 3.062189e-007, 3.334135e-007, 3.592422e-007, 
    3.866851e-007, 4.121412e-007, 4.352382e-007, 4.537403e-007, 
    4.721185e-007, 4.899998e-007, 5.152076e-007, 5.391737e-007, 
    5.590418e-007, 5.743154e-007, 5.854913e-007, 5.909553e-007, 
    5.930663e-007, 5.882232e-007, 5.828836e-007, 5.759298e-007, 
    5.667409e-007, 5.554409e-007, 5.473694e-007, 5.461275e-007, 
    5.528329e-007, 5.623947e-007, 5.751849e-007, 5.878508e-007, 
    5.935628e-007, 5.925697e-007, 5.826353e-007, 5.692243e-007, 
    5.502254e-007, 5.217892e-007, 4.834185e-007, 4.411986e-007, 3.993511e-007,
  3.906587e-007, 3.886719e-007, 3.871818e-007, 3.937632e-007, 4.013378e-007, 
    3.987302e-007, 3.92149e-007, 3.861884e-007, 3.576279e-007, 3.209959e-007, 
    3.006309e-007, 3.044804e-007, 3.19009e-007, 3.310541e-007, 3.267079e-007, 
    3.036111e-007, 2.782792e-007, 2.752989e-007, 3.075848e-007, 
    3.580004e-007, 4.102787e-007, 4.431854e-007, 4.423161e-007, 
    4.262974e-007, 4.084159e-007, 3.752609e-007, 3.247212e-007, 
    2.648682e-007, 2.227723e-007, 2.002964e-007, 1.958261e-007, 
    2.074987e-007, 2.142042e-007, 2.240141e-007, 2.245108e-007, 
    2.348174e-007, 2.703319e-007, 3.320475e-007, 4.148732e-007, 
    5.139659e-007, 6.11196e-007, 6.750225e-007, 7.106612e-007, 7.326405e-007, 
    7.405878e-007, 7.23948e-007, 6.893029e-007, 6.518017e-007, 6.326784e-007, 
    6.442269e-007, 6.910414e-007, 7.441888e-007, 8.101263e-007, 
    8.990366e-007, 1.012534e-006, 1.124293e-006, 1.215686e-006, 
    1.265978e-006, 1.230091e-006, 1.107901e-006, 9.473413e-007, 
    7.907549e-007, 6.190191e-007, 4.35859e-007, 2.579143e-007, 1.338619e-007, 
    1.200785e-007, 2.31589e-007, 3.884234e-007, 5.23776e-007, 5.772959e-007, 
    5.648783e-007, 5.369384e-007, 5.595386e-007, 6.135551e-007, 
    6.370244e-007, 6.499392e-007, 7.186086e-007, 8.761886e-007, 
    1.050284e-006, 1.202027e-006, 1.346444e-006, 1.494338e-006, 
    1.590078e-006, 1.570955e-006, 1.444419e-006, 1.258527e-006, 
    1.061211e-006, 8.819006e-007, 7.284184e-007, 5.969159e-007, 4.94967e-007, 
    4.369767e-007, 4.01338e-007, 3.807245e-007, 3.848224e-007,
  5.032867e-007, 4.931043e-007, 5.313506e-007, 5.407881e-007, 5.077571e-007, 
    4.654129e-007, 3.90783e-007, 2.688419e-007, 1.771997e-007, 1.621743e-007, 
    1.834084e-007, 1.881272e-007, 2.113481e-007, 2.445032e-007, 
    2.523263e-007, 2.698351e-007, 2.803902e-007, 2.52823e-007, 2.150734e-007, 
    1.855194e-007, 1.41561e-007, 1.190851e-007, 1.578281e-007, 1.964469e-007, 
    2.222757e-007, 2.502153e-007, 2.795209e-007, 3.015002e-007, 
    3.444652e-007, 4.010896e-007, 4.212062e-007, 3.757576e-007, 
    3.556411e-007, 3.772477e-007, 3.887961e-007, 3.93639e-007, 3.756334e-007, 
    3.788621e-007, 4.065533e-007, 4.077951e-007, 4.425645e-007, 
    5.637606e-007, 7.017205e-007, 7.783374e-007, 7.549922e-007, 
    7.579724e-007, 9.330611e-007, 1.085301e-006, 1.156082e-006, 
    1.149376e-006, 1.090889e-006, 1.098712e-006, 1.22649e-006, 1.656388e-006, 
    2.325823e-006, 2.748644e-006, 2.54636e-006, 1.840666e-006, 9.985019e-007, 
    4.238141e-007, 2.120928e-007, 1.631674e-007, 1.279013e-007, 
    2.194197e-007, 4.1984e-007, 6.21254e-007, 8.415429e-007, 9.689479e-007, 
    1.006946e-006, 9.465966e-007, 8.97795e-007, 9.06984e-007, 9.458513e-007, 
    1.057237e-006, 1.199295e-006, 1.254554e-006, 1.120568e-006, 8.51353e-007, 
    6.334235e-007, 5.349516e-007, 6.021314e-007, 8.055317e-007, 
    1.089896e-006, 1.419211e-006, 1.653656e-006, 1.711647e-006, 1.74207e-006, 
    1.864384e-006, 1.950562e-006, 1.851221e-006, 1.510854e-006, 
    1.087164e-006, 7.759779e-007, 6.136795e-007, 5.85243e-007, 5.671134e-007,
  5.631398e-007, 5.49977e-007, 4.813076e-007, 4.727393e-007, 4.187226e-007, 
    3.237277e-007, 2.786517e-007, 3.304333e-007, 4.197161e-007, 
    4.931043e-007, 5.579244e-007, 5.60532e-007, 5.492319e-007, 4.821767e-007, 
    4.181018e-007, 4.256765e-007, 4.528711e-007, 4.318853e-007, 
    3.813456e-007, 3.914039e-007, 3.347794e-007, 2.236416e-007, 
    1.408159e-007, 4.308913e-008, 4.867718e-008, 5.4265e-008, 7.54992e-008, 
    1.400709e-007, 2.137075e-007, 2.923111e-007, 3.777444e-007, 
    3.863126e-007, 4.116446e-007, 4.994372e-007, 5.808969e-007, 
    6.185223e-007, 6.254762e-007, 7.639329e-007, 9.586414e-007, 
    9.634842e-007, 8.237859e-007, 8.169561e-007, 1.009678e-006, 
    1.265729e-006, 1.501789e-006, 1.81136e-006, 2.251441e-006, 2.662961e-006, 
    2.505009e-006, 1.995762e-006, 1.24077e-006, 8.096295e-007, 8.525949e-007, 
    1.320119e-006, 1.646081e-006, 1.748652e-006, 1.444295e-006, 
    9.895612e-007, 6.38639e-007, 2.358111e-007, -1.549715e-007, 
    -6.372729e-007, -1.42542e-006, -1.863265e-006, -1.649682e-006, 
    -1.202027e-006, -6.660821e-007, -3.085779e-007, -3.664445e-007, 
    -8.929519e-007, -1.299257e-006, -1.148507e-006, -4.061812e-007, 
    4.755957e-007, 1.259893e-006, 1.971051e-006, 2.622231e-006, 
    2.841652e-006, 2.667184e-006, 2.330417e-006, 2.089267e-006, 
    2.073249e-006, 2.05338e-006, 1.865128e-006, 1.873946e-006, 1.91393e-006, 
    1.618266e-006, 1.421322e-006, 1.642729e-006, 1.853704e-006, 
    1.923615e-006, 1.693393e-006, 1.392637e-006, 1.191844e-006, 
    9.655953e-007, 6.783753e-007,
  1.016011e-006, 8.66999e-007, 9.691964e-007, 1.071766e-006, 1.136338e-006, 
    1.105294e-006, 9.674579e-007, 6.889302e-007, 7.467966e-007, 
    9.454786e-007, 1.050283e-006, 1.027311e-006, 6.721666e-007, 
    3.032385e-007, 2.897034e-007, 5.010514e-007, 5.605319e-007, 
    4.418195e-007, 2.85233e-007, 1.899898e-007, 3.300606e-007, 5.17691e-007, 
    4.510086e-007, 2.651166e-007, 6.829623e-009, -1.151116e-007, 
    -1.693766e-007, 1.182159e-007, 5.772956e-007, 7.275491e-007, 
    5.980332e-007, 6.222479e-007, 9.201469e-007, 1.037121e-006, 
    7.951012e-007, 5.866091e-007, 8.688621e-007, 1.393631e-006, 
    1.909336e-006, 2.306452e-006, 2.48154e-006, 2.857049e-006, 3.489107e-006, 
    4.383922e-006, 5.060558e-006, 5.074715e-006, 4.685049e-006, 
    4.211317e-006, 3.965323e-006, 3.506366e-006, 3.441299e-006, 
    3.591179e-006, 4.096702e-006, 5.072727e-006, 5.154932e-006, 
    3.893672e-006, 2.438825e-006, 2.346684e-006, 2.72741e-006, 3.00544e-006, 
    3.056724e-006, 2.942111e-006, 1.912565e-006, 6.639712e-007, 
    -6.618602e-007, -1.65763e-006, -2.143283e-006, -2.340227e-006, 
    -1.963477e-006, -9.58642e-007, -4.764652e-007, 4.979483e-008, 
    1.592313e-006, 2.255167e-006, 2.227227e-006, 2.456084e-006, 
    2.756839e-006, 2.700463e-006, 3.068521e-006, 4.001086e-006, 
    4.351387e-006, 3.641098e-006, 2.736226e-006, 2.76578e-006, 3.384426e-006, 
    4.062554e-006, 3.711259e-006, 2.903864e-006, 1.929949e-006, 
    1.239032e-006, 2.108638e-006, 2.826999e-006, 3.593664e-006, 
    3.255904e-006, 2.301236e-006, 1.528238e-006,
  1.857802e-006, 2.238403e-006, 2.779935e-006, 3.30098e-006, 3.314143e-006, 
    3.24448e-006, 3.115957e-006, 2.683699e-006, 2.089764e-006, 2.577653e-006, 
    2.955646e-006, 3.265092e-006, 3.57839e-006, 3.562371e-006, 2.637257e-006, 
    1.925727e-006, 1.765043e-006, 1.514082e-006, 1.604482e-006, 
    2.139807e-006, 2.310797e-006, 2.184386e-006, 1.431629e-006, 
    7.823019e-009, -1.061584e-006, -1.516938e-006, -1.646827e-006, 
    -1.506011e-006, -9.74288e-007, -2.510842e-007, 5.344546e-007, 
    7.260587e-007, 1.458451e-006, 2.556542e-006, 3.369153e-006, 
    4.837166e-006, 5.829583e-006, 5.715217e-006, 6.472692e-006, 7.13505e-006, 
    7.52161e-006, 7.928411e-006, 7.242088e-006, 6.592274e-006, 7.656465e-006, 
    8.72376e-006, 9.54618e-006, 8.909155e-006, 6.595999e-006, 4.995491e-006, 
    5.508711e-006, 6.209315e-006, 6.310393e-006, 5.570302e-006, 
    5.031874e-006, 3.954396e-006, 3.385295e-006, 3.59801e-006, 3.634393e-006, 
    2.82998e-006, 1.2286e-006, 6.270902e-007, 9.940322e-007, 1.262377e-006, 
    1.575921e-006, 1.871585e-006, 1.667067e-006, 1.907845e-006, 
    1.922995e-006, 2.606958e-006, 2.93764e-006, 2.205993e-006, 9.123232e-007, 
    4.106505e-007, 4.656613e-007, 2.148127e-006, 4.065284e-006, 
    5.424396e-006, 5.919363e-006, 5.702922e-006, 4.761541e-006, 
    3.298001e-006, 2.950182e-006, 3.277014e-006, 3.611297e-006, 
    3.022825e-006, 2.724057e-006, 2.318248e-006, 2.141794e-006, 
    2.026683e-006, 2.396479e-006, 2.919137e-006, 3.389765e-006, 
    2.863382e-006, 2.634525e-006, 2.028421e-006,
  3.418575e-006, 3.329913e-006, 3.21952e-006, 3.309298e-006, 3.052379e-006, 
    3.598381e-006, 3.857042e-006, 3.124276e-006, 3.530955e-006, 
    4.784019e-006, 5.602589e-006, 5.506105e-006, 5.927557e-006, 
    7.395072e-006, 7.574012e-006, 6.81281e-006, 6.800145e-006, 7.46188e-006, 
    8.558358e-006, 9.079402e-006, 7.698934e-006, 5.701929e-006, 
    4.283712e-006, 3.669039e-006, 2.587462e-006, 1.544506e-006, 
    5.725769e-007, -3.000096e-007, -6.308155e-007, -4.965841e-010, 
    1.486515e-006, 1.241391e-006, 9.192772e-007, 1.147266e-006, 
    3.699461e-006, 4.820029e-006, 6.779657e-006, 8.820989e-006, 
    8.159255e-006, 6.534654e-006, 8.04427e-006, 8.647639e-006, 8.000432e-006, 
    1.013465e-005, 1.147625e-005, 9.603176e-006, 8.125602e-006, 
    6.566197e-006, 4.810965e-006, 5.90769e-006, 6.923949e-006, 5.817785e-006, 
    5.279358e-006, 5.942211e-006, 6.605809e-006, 6.777916e-006, 7.29151e-006, 
    6.462757e-006, 5.289663e-006, 3.841145e-006, 3.134211e-006, 
    2.640238e-006, 2.491351e-006, 3.787628e-006, 4.675363e-006, 
    4.903102e-006, 5.010018e-006, 4.761914e-006, 4.078448e-006, 4.51915e-006, 
    5.675975e-006, 5.710746e-006, 5.099302e-006, 5.055468e-006, 
    5.111595e-006, 5.329524e-006, 5.430231e-006, 6.277734e-006, 7.37831e-006, 
    5.733966e-006, 4.75049e-006, 5.03535e-006, 5.35672e-006, 5.738438e-006, 
    5.490333e-006, 4.061436e-006, 3.769621e-006, 3.36518e-006, 3.324946e-006, 
    3.196299e-006, 3.069267e-006, 2.262988e-006, 1.046434e-006, 
    7.800763e-007, 2.122049e-006, 3.214802e-006,
  3.825749e-006, 3.857042e-006, 2.88623e-006, 3.309548e-006, 3.103416e-006, 
    2.148872e-006, 3.685431e-006, 5.51405e-006, 6.215398e-006, 4.832074e-006, 
    3.880261e-006, 4.799291e-006, 5.490332e-006, 7.496899e-006, 
    9.100513e-006, 1.086804e-005, 1.180284e-005, 1.171331e-005, 
    9.542084e-006, 6.836031e-006, 6.148965e-006, 5.322694e-006, 
    5.623946e-006, 6.078806e-006, 7.085873e-006, 7.404264e-006, 6.45804e-006, 
    6.063903e-006, 5.175172e-006, 3.586214e-006, 2.848356e-006, 
    3.157058e-006, 2.624094e-006, 3.112727e-006, 5.660953e-006, 
    6.928294e-006, 5.358334e-006, 6.287173e-006, 6.172681e-006, 
    4.638854e-006, 5.416698e-006, 6.54223e-006, 8.197378e-006, 8.793049e-006, 
    7.779772e-006, 5.496915e-006, 4.410249e-006, 5.941838e-006, 
    4.852687e-006, 4.219015e-006, 4.383797e-006, 3.771856e-006, 
    3.791352e-006, 4.129237e-006, 3.204372e-006, 1.938393e-006, 
    1.859293e-006, 1.654153e-006, 2.809615e-006, 5.336726e-006, 
    4.865229e-006, 4.272288e-006, 3.535548e-006, 2.168863e-006, 
    1.414741e-006, 2.061452e-006, 3.335377e-006, 3.393865e-006, 
    4.747386e-006, 6.527578e-006, 8.723513e-006, 8.129949e-006, 
    6.577746e-006, 7.235756e-006, 8.164594e-006, 6.614127e-006, 
    5.764763e-006, 7.084138e-006, 8.434803e-006, 7.235631e-006, 
    6.555891e-006, 7.066999e-006, 6.769969e-006, 5.842372e-006, 
    5.619104e-006, 5.659833e-006, 5.106256e-006, 4.714106e-006, 
    4.050757e-006, 3.442292e-006, 3.050392e-006, 2.322222e-006, 
    2.417838e-006, 3.745407e-006, 3.243236e-006, 3.4449e-006,
  4.292155e-006, 4.668782e-006, 4.12191e-006, 5.536403e-006, 6.805485e-006, 
    4.788737e-006, 4.911424e-006, 6.540615e-006, 6.675844e-006, 6.51305e-006, 
    6.672492e-006, 8.189803e-006, 1.080272e-005, 1.210533e-005, 
    1.239267e-005, 1.27087e-005, 1.316965e-005, 1.271864e-005, 1.114619e-005, 
    9.13019e-006, 8.59946e-006, 9.067979e-006, 8.776784e-006, 8.590891e-006, 
    1.004338e-005, 1.071965e-005, 9.259211e-006, 8.37172e-006, 7.308276e-006, 
    8.918096e-006, 8.200483e-006, 5.664429e-006, 7.090468e-006, 
    8.110081e-006, 5.295376e-006, 3.107391e-006, 4.552552e-006, 
    6.610033e-006, 4.983443e-006, 3.551197e-006, 5.780161e-006, 5.23093e-006, 
    6.208071e-006, 6.241973e-006, 4.738818e-006, 2.913055e-006, 
    5.066518e-006, 4.970283e-006, 3.820658e-006, 2.122299e-006, 
    2.589697e-006, 4.05858e-006, 3.578638e-006, 2.549465e-006, 3.279747e-006, 
    2.008552e-006, 1.769513e-006, 2.576659e-006, 2.808869e-006, 
    4.055601e-006, 1.816328e-006, 7.467952e-007, 1.05401e-006, 2.437086e-006, 
    3.531079e-006, 4.062678e-006, 4.037965e-006, 4.390378e-006, 
    5.178526e-006, 4.357224e-006, 4.277379e-006, 4.396215e-006, 
    3.998477e-006, 4.026293e-006, 4.892052e-006, 5.283207e-006, 
    5.447491e-006, 6.53751e-006, 5.419923e-006, 2.656134e-006, 1.910701e-006, 
    1.989429e-006, 1.497319e-006, 2.238899e-006, 3.16327e-006, 3.353631e-006, 
    3.744537e-006, 3.923476e-006, 3.094598e-006, 2.026683e-006, 
    2.095972e-006, 3.233677e-006, 3.316874e-006, 2.793224e-006, 
    3.553057e-006, 4.469604e-006,
  5.971764e-006, 6.948037e-006, 6.51926e-006, 5.645677e-006, 6.367018e-006, 
    7.139519e-006, 7.313862e-006, 6.527081e-006, 4.025551e-006, 
    5.019952e-006, 7.591647e-006, 9.923306e-006, 1.193248e-005, 
    1.211539e-005, 1.116929e-005, 9.477633e-006, 8.960442e-006, 
    7.562216e-006, 7.585932e-006, 8.315219e-006, 9.058167e-006, 
    1.025709e-005, 1.13948e-005, 1.079266e-005, 9.141117e-006, 9.75691e-006, 
    1.116283e-005, 1.025299e-005, 8.303796e-006, 7.958337e-006, 
    8.630999e-006, 7.700921e-006, 5.743404e-006, 3.372876e-006, 
    3.554054e-006, 4.512323e-006, 7.47728e-006, 8.226933e-006, 4.018471e-006, 
    2.703815e-006, 3.335128e-006, 5.945314e-006, 7.993229e-006, 
    9.615345e-006, 5.44178e-006, 3.915779e-006, 4.296377e-006, 2.113233e-006, 
    3.194436e-006, 3.026425e-006, 3.703559e-006, 2.383564e-006, 
    -1.141552e-006, -1.412134e-006, -1.448145e-006, -1.478444e-006, 
    2.222012e-006, 4.720066e-006, 3.886224e-006, 2.060955e-006, 
    -8.704774e-007, -1.804281e-006, -1.080582e-006, 1.302735e-006, 
    -3.278255e-007, -4.337489e-007, 1.406297e-006, 1.767403e-006, 
    5.813945e-007, 1.834458e-006, 5.971639e-006, 8.126472e-006, 
    5.857399e-006, 6.221979e-006, 5.957238e-006, 3.897028e-006, 
    3.652276e-006, 3.482279e-006, 2.585226e-006, 2.009165e-007, 
    -1.565366e-006, 1.480304e-006, 2.551948e-006, 1.025201e-006, 
    1.681845e-006, 1.945098e-006, 9.690721e-007, 7.700164e-007, 
    9.602554e-007, 1.975646e-006, 3.021954e-006, 3.819789e-006, 
    4.396339e-006, 4.355237e-006, 6.310765e-006, 6.96741e-006,
  5.511441e-006, 7.02354e-006, 7.035957e-006, 8.002917e-006, 7.251401e-006, 
    6.638591e-006, 5.784132e-006, 6.876016e-006, 6.948536e-006, 
    8.728606e-006, 9.60541e-006, 1.051873e-005, 1.023114e-005, 7.89476e-006, 
    6.799026e-006, 8.940697e-006, 1.055077e-005, 1.032948e-005, 
    9.925539e-006, 1.130067e-005, 1.122678e-005, 9.660547e-006, 
    1.072747e-005, 9.841842e-006, 9.32589e-006, 8.692965e-006, 8.364645e-006, 
    8.993349e-006, 8.767594e-006, 7.60605e-006, 5.334867e-006, 3.690646e-006, 
    2.530218e-006, 3.354377e-006, 6.506965e-006, 6.411348e-006, 
    5.374477e-006, 3.804515e-006, 1.090266e-006, 5.801521e-007, 
    3.916895e-006, 5.339336e-006, 5.47655e-006, 3.323084e-006, 2.132107e-006, 
    3.539026e-007, -2.452471e-007, 1.393755e-006, -1.178683e-006, 
    -1.013403e-006, -2.449997e-007, -3.861878e-007, -3.522386e-006, 
    -1.266102e-006, -3.297626e-006, -2.261997e-006, -6.904211e-007, 
    -8.586794e-007, 2.514944e-006, 1.479561e-006, 9.165451e-007, 
    1.252567e-006, 2.467756e-006, 1.567974e-006, 2.983461e-006, 
    3.236781e-006, 3.242616e-006, 2.936147e-006, 4.61638e-006, 2.639616e-006, 
    2.066419e-006, 2.880395e-006, 4.965685e-006, 3.384925e-006, 
    1.352651e-006, 4.029273e-006, 6.123879e-006, 3.659228e-006, 
    1.809622e-006, -1.743429e-007, -1.94932e-006, -1.432001e-006, 
    5.102411e-007, 8.857496e-007, 9.916712e-007, 1.825889e-006, 
    3.450737e-006, 4.53728e-006, 4.921731e-006, 4.420057e-006, 3.519781e-006, 
    4.642705e-006, 5.220872e-006, 6.142755e-006, 5.125006e-006, 3.687044e-006,
  7.417304e-006, 5.565085e-006, 5.351005e-006, 6.466111e-006, 5.64431e-006, 
    5.142887e-006, 5.962202e-006, 5.602711e-006, 6.558623e-006, 
    6.219992e-006, 6.928545e-006, 7.763507e-006, 6.904575e-006, 
    7.943934e-006, 8.615105e-006, 9.092688e-006, 9.023275e-006, 
    7.282695e-006, 7.308645e-006, 7.320446e-006, 8.479878e-006, 
    7.949395e-006, 7.16274e-006, 5.68293e-006, 5.335238e-006, 5.267189e-006, 
    5.574402e-006, 4.81978e-006, 1.812354e-006, 7.294111e-007, 
    -1.101569e-006, -1.692399e-006, -2.13931e-006, -1.444172e-006, 
    -5.548209e-007, -3.601126e-007, -4.181391e-006, -3.694742e-006, 
    -2.110126e-006, -1.449884e-006, 4.831709e-007, 3.1321e-006, 5.09446e-006, 
    4.186108e-006, 9.415053e-007, 2.134097e-006, -1.692533e-007, 
    -2.135585e-006, -6.635983e-007, 1.615037e-006, 3.848218e-007, 
    -3.717467e-006, -5.896018e-006, -6.184106e-006, -7.553896e-006, 
    -4.560748e-006, -1.177315e-006, -6.896753e-007, 8.811548e-007, 
    7.490307e-007, -9.470932e-007, -1.525877e-006, 5.992752e-007, 
    1.462799e-006, 5.790353e-007, 5.085021e-007, 4.2703e-006, 2.475826e-006, 
    4.495159e-007, 2.650046e-006, 2.38642e-006, 2.672896e-006, 3.535315e-007, 
    -1.455595e-006, 1.543882e-006, 5.578622e-006, 2.498928e-006, 
    -9.648284e-008, -3.207479e-007, 2.646193e-007, 8.439019e-007, 
    -2.284833e-008, 1.319373e-006, 1.569961e-006, 2.890949e-006, 
    4.978105e-006, 6.637349e-006, 6.811817e-006, 7.186085e-006, 
    6.499144e-006, 4.251051e-006, 2.857174e-006, 2.143406e-006, 
    2.870958e-006, 4.060192e-006, 7.266801e-006,
  5.465125e-006, 6.273513e-006, 4.664063e-006, 4.547328e-007, 2.921992e-006, 
    7.103385e-006, 8.057681e-006, 8.944173e-006, 7.538123e-006, 
    9.295343e-006, 9.445224e-006, 1.106275e-005, 9.736916e-006, 
    7.387749e-006, 6.321319e-006, 5.300219e-006, 3.300356e-006, 
    1.801302e-006, 3.032885e-006, 1.950561e-006, 2.829358e-006, 
    2.508736e-006, 2.152472e-006, -1.962853e-006, -4.227459e-006, 
    -7.466351e-006, -9.39754e-006, -9.363517e-006, -9.276468e-006, 
    -8.872896e-006, -8.778525e-006, -6.445995e-006, -6.294498e-006, 
    -7.108598e-006, -8.046005e-006, -8.510302e-006, -7.016955e-006, 
    -5.901853e-006, -4.218891e-006, -2.276523e-006, -1.826509e-006, 
    2.893681e-006, 5.429238e-006, 3.571557e-006, 1.848613e-006, 
    1.341599e-006, 1.833465e-006, 4.376099e-006, 5.184982e-006, 
    2.570079e-006, -2.840035e-006, -4.862497e-006, -5.243346e-006, 
    -4.442285e-006, -3.906836e-006, -2.313529e-006, -3.901245e-006, 
    -4.340334e-006, -2.125278e-006, 8.088864e-007, -1.156703e-006, 
    2.723209e-007, 2.1905e-007, 5.734473e-007, 7.723756e-007, -5.47243e-007, 
    1.945842e-006, 4.114212e-006, 2.550336e-006, 2.308436e-006, 
    1.562265e-006, -3.448367e-007, 1.760571e-006, -2.426386e-007, 
    -8.806601e-007, -2.036741e-006, -3.356487e-006, -2.038974e-006, 
    -7.686522e-007, 3.029778e-006, 1.617273e-006, 2.173583e-006, 
    4.213056e-006, 2.559274e-006, 5.742782e-006, 9.759391e-006, 
    9.307514e-006, 6.971135e-006, 5.437312e-006, 1.69126e-007, 5.476177e-007, 
    1.691158e-006, -6.340451e-007, -6.545342e-007, 2.822406e-006, 
    3.506244e-006,
  1.185013e-006, 1.503526e-006, 1.246233e-006, 1.53333e-006, 2.512212e-006, 
    3.732121e-006, 4.936755e-006, 4.24795e-006, 4.346544e-006, 5.262966e-006, 
    5.287056e-006, 2.73039e-006, -2.51544e-006, -4.678346e-006, 
    -3.823887e-006, -4.364178e-006, -5.00977e-006, -2.577654e-006, 
    -8.713469e-007, -6.556511e-007, -5.007785e-006, -6.852297e-006, 
    -7.930399e-006, -8.435423e-006, -9.566422e-006, -8.902327e-006, 
    -8.154535e-006, -8.303425e-006, -8.004779e-006, -5.430977e-006, 
    -4.86349e-006, -7.623681e-006, -9.566918e-006, -8.928899e-006, 
    -1.052283e-005, -9.616464e-006, -6.250168e-006, -4.540387e-006, 
    -4.865728e-006, -3.243113e-006, -1.848241e-006, 1.656264e-006, 
    6.417558e-006, 9.526811e-006, 5.391488e-006, 2.755969e-006, 
    5.245085e-006, 6.235266e-006, 6.576131e-006, 3.212193e-006, 
    -4.102909e-006, -8.431576e-006, -7.354469e-006, -7.613995e-006, 
    -3.69189e-006, -5.907317e-006, -7.057315e-006, -1.555931e-006, 
    2.926827e-007, 1.852957e-006, 1.687557e-006, 1.472235e-006, 
    2.806337e-008, 2.145272e-006, 3.04915e-006, 2.321478e-006, 1.034638e-006, 
    2.675006e-006, 1.446777e-006, 1.568471e-006, 4.844118e-006, 
    5.825983e-006, 3.767509e-006, 1.435477e-006, -1.40605e-006, 
    -2.078959e-006, -5.960963e-006, -6.832059e-006, -1.818686e-006, 
    2.432986e-006, 2.499793e-006, 4.434462e-006, 4.055599e-006, 
    4.947557e-006, 5.857644e-006, 4.042064e-006, 4.686914e-006, 
    4.177542e-006, 2.127141e-006, 2.564266e-007, -8.961797e-007, 
    -2.137822e-006, -4.071735e-007, -2.674788e-007, -1.793105e-006, 
    -8.158531e-008,
  -8.795414e-007, -1.087785e-006, -1.085675e-006, -2.172962e-006, 
    -1.381462e-006, -1.236913e-010, -2.74802e-007, -3.522873e-007, 
    -1.118705e-006, -2.044564e-006, -1.111639e-005, -1.303901e-005, 
    -1.080818e-005, -9.635836e-006, -8.283803e-006, -6.293629e-006, 
    -4.030391e-006, -2.707167e-006, -3.402929e-006, -6.03286e-006, 
    -8.410962e-006, -8.217743e-006, -6.400795e-006, -5.114326e-006, 
    -4.683187e-006, -4.376099e-006, -5.546584e-006, -4.788984e-006, 
    -3.550202e-006, -4.058456e-006, -5.985425e-006, -8.835892e-006, 
    -7.72501e-006, -7.29151e-006, -5.904958e-006, -4.070003e-006, 
    -3.642464e-006, -1.447523e-006, -7.482868e-007, 1.274422e-006, 
    3.242865e-006, 4.793579e-006, 1.057858e-005, 1.25392e-005, 1.010758e-005, 
    7.56979e-006, 6.9987e-006, 2.334265e-006, -2.75001e-006, -6.140272e-006, 
    -8.086117e-006, -9.969248e-006, -9.824707e-006, -7.800882e-006, 
    -1.158652e-005, -6.577498e-006, -4.576519e-006, 4.872709e-007, 
    4.534548e-006, 5.99238e-006, 6.849317e-006, 1.006362e-005, 6.426992e-006, 
    4.905836e-006, 6.525468e-006, 6.707385e-006, 5.455691e-006, 
    4.036599e-006, -3.609428e-006, 1.143788e-006, 4.659221e-006, 
    2.50799e-006, 1.610068e-006, 6.105729e-007, -7.116541e-007, 
    -8.600455e-007, -4.170462e-006, -5.966549e-006, 1.950812e-007, 
    3.52909e-006, 8.914612e-007, -1.809623e-006, 1.34396e-006, 3.489356e-006, 
    3.496436e-006, 1.979388e-007, -2.360717e-006, -4.209829e-006, 
    -3.820907e-006, -2.860277e-006, -1.956276e-006, -2.674384e-006, 
    -3.851575e-006, -2.937517e-006, -3.642466e-006, -1.053388e-006,
  -2.194941e-006, -1.785656e-006, -1.345823e-006, -6.880609e-007, 
    8.592997e-008, -1.743438e-007, -1.637141e-006, 1.396984e-007, 
    1.895428e-006, -1.782801e-006, -6.424387e-006, -5.975116e-006, 
    -5.2616e-006, -8.91586e-006, -8.488447e-006, -4.396961e-006, 
    -4.836791e-006, -5.627548e-006, -2.534316e-006, -7.177387e-007, 
    -3.004321e-006, -5.053971e-007, -9.727974e-007, -1.870964e-006, 
    -8.411698e-007, -9.962669e-007, -2.690653e-006, -2.847115e-006, 
    -2.725174e-006, -4.449115e-006, -8.410463e-006, -5.955746e-006, 
    -2.881016e-006, -1.953169e-006, -2.029786e-006, -1.140808e-006, 
    -4.687663e-007, 1.544878e-006, 3.177301e-006, 2.694627e-006, 
    1.842653e-006, 3.123532e-006, 5.017344e-006, 2.287081e-006, 
    9.783871e-007, 1.154094e-006, 1.425047e-006, -1.428154e-006, 
    -7.179879e-006, -8.011237e-006, -4.649908e-006, -4.31513e-006, 
    -5.125999e-006, -6.070608e-006, -9.455038e-006, -6.275746e-006, 
    -2.998986e-006, 3.031517e-006, 8.510302e-006, 9.917345e-006, 
    1.381698e-005, 1.015912e-005, 8.075061e-006, 1.009094e-005, 
    8.384755e-006, 8.280324e-006, 6.841372e-006, 2.528603e-006, 
    2.009423e-006, 3.710516e-006, 2.506502e-006, 1.462549e-006, 
    1.166387e-006, -1.641114e-006, -2.701084e-006, -3.924842e-006, 
    -4.271542e-006, -2.156446e-006, -6.819769e-007, -3.897274e-006, 
    -3.434967e-006, -2.899764e-006, -4.047652e-006, -2.565979e-006, 
    -2.826378e-006, -2.02718e-006, -3.411746e-006, -6.087868e-006, 
    -4.742295e-006, -6.15418e-006, -4.322454e-006, -4.549325e-006, 
    -4.482021e-006, -3.328299e-006, -1.986447e-006, -1.743809e-006,
  -1.423929e-006, -1.914426e-006, -6.958844e-007, -2.391635e-007, 
    -5.616496e-007, -1.29876e-006, -9.00277e-008, -4.009653e-007, 
    1.238162e-006, -4.240994e-006, -7.341925e-006, -6.876514e-006, 
    -4.900372e-006, -7.748604e-006, -5.732105e-006, -3.45471e-006, 
    -1.170984e-006, 2.260382e-006, 3.234172e-006, -3.407404e-007, 
    -3.182142e-006, -2.506625e-006, -1.823032e-006, -6.793689e-007, 
    9.713076e-007, -1.26573e-006, -3.449122e-006, -4.30035e-006, 
    -3.599375e-006, -5.361687e-006, -6.447733e-006, -2.617761e-006, 
    -1.438956e-006, 6.397563e-007, 2.198542e-006, 3.60782e-006, 
    3.662581e-006, 3.532817e-006, 3.928567e-006, 5.513057e-006, 
    6.738181e-006, 3.966565e-006, -1.667191e-006, -1.795714e-006, 
    -2.818431e-006, -1.16378e-006, -4.004316e-006, -5.260234e-006, 
    -1.640368e-006, 1.707671e-006, 2.130124e-006, -2.828365e-006, 
    -7.833169e-006, -1.046459e-005, -9.705251e-006, -6.26122e-006, 
    -2.04593e-006, 9.891886e-006, 1.851867e-005, 1.746081e-005, 
    1.265643e-005, 1.326911e-005, 1.22613e-005, 9.32589e-006, 3.005069e-006, 
    5.655733e-006, 6.250291e-006, 4.834183e-006, 1.272932e-006, 
    9.957694e-007, -1.034015e-006, -1.604731e-006, -1.645833e-006, 
    -2.313902e-006, -2.454966e-006, -1.347189e-006, -1.028056e-006, 
    4.244348e-007, 1.245489e-007, -6.428981e-006, -6.683791e-006, 
    -1.179464e-005, -1.349275e-005, -1.056045e-005, -1.085302e-006, 
    -2.103299e-006, -5.023057e-006, -2.633905e-006, -1.302609e-006, 
    -1.152729e-006, -2.82824e-006, -3.283968e-006, -1.537179e-006, 
    -2.165511e-006, -1.43225e-006, -1.6621e-006,
  -6.91165e-007, -5.833799e-007, 7.064396e-007, -4.433093e-008, 
    -2.286087e-007, 1.45285e-008, -1.497569e-007, -1.783793e-006, 
    -1.75101e-006, -2.16191e-006, -3.977989e-006, -2.917895e-006, 
    -2.472599e-006, -7.440398e-006, -1.004711e-005, -6.509821e-006, 
    -2.170727e-006, 6.793689e-007, 7.326398e-007, 1.620625e-006, 
    -5.304564e-006, -2.882132e-006, -6.172813e-007, -1.617893e-006, 
    -4.635379e-006, -5.332505e-006, -1.418963e-006, -6.361552e-007, 
    -1.258775e-006, -4.043306e-006, -2.809365e-006, 1.032402e-006, 
    2.826378e-006, 5.51045e-006, 5.459785e-006, 3.40119e-006, 5.656853e-006, 
    6.882598e-006, 5.021071e-006, 5.358954e-006, 6.223718e-006, 
    3.422549e-006, 2.276525e-006, 4.072612e-006, 2.058347e-006, 
    -3.124896e-006, -5.48698e-006, -4.984811e-006, -1.234066e-006, 
    1.28361e-006, -6.172813e-007, -3.20586e-006, -6.753828e-006, 
    -4.375477e-006, 1.315151e-006, 8.911142e-006, 1.697329e-005, 
    1.662337e-005, 1.347971e-005, 1.215575e-005, 1.004425e-005, 
    4.584963e-006, 2.426281e-006, 2.490853e-006, 3.742054e-006, 
    1.943732e-006, 2.533072e-006, 9.859596e-007, -1.87233e-006, 
    -1.795342e-006, -1.984959e-006, -1.933922e-006, -1.770134e-006, 
    -1.837561e-006, -7.37359e-007, 2.646198e-007, 1.882141e-006, 
    1.558041e-006, 1.860286e-006, -3.8784e-006, -8.998563e-006, 
    -1.019475e-005, -6.14586e-006, -5.08378e-006, -3.091245e-006, 
    -3.444776e-006, -3.566468e-006, -4.947178e-007, -1.531094e-006, 
    -1.693144e-006, -1.593678e-006, -1.252692e-006, -3.080071e-006, 
    -2.299124e-006, -9.037549e-007, -1.19855e-006,
  -5.671136e-007, 1.353524e-007, -3.460796e-007, -1.401951e-007, 
    -5.215406e-008, 2.310923e-007, -2.127141e-007, -7.364898e-007, 
    -1.117587e-006, -3.09435e-006, -3.21207e-006, -2.246225e-006, 
    -4.324938e-006, -6.104012e-006, -4.660586e-006, 1.490116e-008, 
    4.834201e-007, -1.396611e-006, -3.669782e-006, -2.701952e-006, 
    -6.614864e-007, -9.801242e-007, -8.260213e-007, -3.380454e-006, 
    -5.770847e-006, -1.779448e-006, 2.715742e-007, -9.985015e-007, 
    -1.147639e-006, -1.978626e-006, 5.998959e-007, 3.562868e-006, 
    4.311775e-006, 4.300351e-006, 4.103159e-006, 5.239496e-006, 
    6.343673e-006, 3.966316e-006, 2.79285e-006, 3.393119e-006, 1.849482e-006, 
    2.174079e-006, 1.890585e-006, 2.167498e-006, -2.213692e-006, 
    -4.787122e-006, -4.050011e-006, -2.584233e-006, -1.463417e-006, 
    -1.014769e-006, -4.214296e-006, -4.46886e-006, -4.854304e-006, 
    -1.977012e-006, 7.924933e-006, 1.216742e-005, 9.803845e-006, 
    8.520732e-006, 5.602713e-006, 4.92682e-006, 3.972029e-006, 1.24996e-006, 
    -7.505223e-007, -1.723318e-006, -6.817208e-008, -5.621469e-007, 
    -1.836568e-006, -1.415486e-006, -6.788723e-007, -1.334151e-006, 
    -2.082189e-006, -8.322295e-007, -1.442309e-006, -1.483909e-007, 
    8.692382e-009, 1.883258e-006, 2.162034e-006, 1.317635e-006, 
    1.434486e-006, -5.522494e-006, -5.995234e-006, -4.362563e-006, 
    -2.570699e-006, -2.387414e-006, -3.581494e-006, -2.552692e-006, 
    -2.136578e-006, -8.694769e-010, 6.711734e-007, 7.587187e-008, 
    -1.335517e-006, -1.329059e-006, -1.275167e-006, -9.946507e-008, 
    -3.279501e-007, -1.045564e-007,
  -1.245489e-006, -6.32554e-007, -1.298886e-007, 4.234413e-008, 1.73226e-007, 
    2.539407e-007, -2.859781e-007, 6.755198e-008, -1.060838e-006, 
    -1.114358e-006, -1.754487e-006, -1.959751e-006, -1.640245e-006, 
    -1.985331e-006, -4.091238e-006, -2.281122e-007, -1.126031e-006, 
    -2.484023e-006, 6.279588e-007, 1.507502e-006, 2.108762e-006, 
    2.334764e-006, -7.713834e-007, -1.696126e-006, -1.047675e-006, 
    -7.135168e-007, -4.079193e-007, -3.211198e-007, -1.376868e-006, 
    -1.662721e-006, 2.048537e-006, 2.641728e-006, 1.2589e-006, 1.187126e-006, 
    1.402324e-006, 2.545615e-006, 8.92828e-007, 1.127273e-006, 1.428152e-006, 
    -1.074995e-006, 5.029142e-007, 2.630179e-006, 8.910893e-007, 
    -2.523139e-006, -4.084656e-006, -2.660727e-006, -4.686415e-006, 
    -4.947557e-006, -4.298241e-006, -6.175536e-006, -8.250523e-006, 
    -6.061544e-006, -2.846369e-006, 2.360219e-006, 7.884455e-006, 
    7.731096e-006, 5.920232e-006, 3.320227e-006, 2.106404e-006, 
    2.454593e-006, 1.711399e-006, 5.74315e-007, -2.734487e-006, 
    -1.341974e-006, -2.639741e-006, -2.089019e-006, -2.606958e-006, 
    -2.721946e-006, -2.272179e-006, -2.642597e-006, -8.665029e-007, 
    -1.298015e-006, -7.952253e-007, -1.188369e-007, -5.568068e-007, 
    1.417597e-006, 9.407601e-007, 1.420205e-006, -5.410486e-006, 
    -9.546429e-006, -3.061444e-006, -9.981295e-007, -1.465033e-006, 
    -9.309501e-007, -3.677234e-006, -4.070997e-006, -4.759677e-007, 
    2.628937e-006, 1.503278e-006, 7.229555e-007, -1.149998e-006, 
    4.637986e-007, 8.717143e-008, 1.850221e-007, -1.049662e-006, 
    -1.995513e-007,
  -1.531467e-006, -1.158441e-006, -4.969537e-007, -6.183983e-008, 
    2.570454e-008, 2.001723e-007, 1.322477e-007, 6.978712e-008, 
    -5.215407e-007, -8.307397e-007, -1.952673e-006, -1.331542e-006, 
    -1.915296e-006, -2.361337e-006, -4.659842e-006, -1.909708e-006, 
    -8.6402e-007, 1.244993e-006, 6.357581e-006, 7.268165e-006, 4.47755e-006, 
    2.305955e-006, 2.102306e-006, 7.27674e-007, -8.481256e-007, 
    9.084742e-007, 7.680301e-007, 8.78299e-007, -1.139319e-006, 
    -1.478195e-006, 1.482914e-006, 2.285217e-006, 1.785035e-006, 
    1.115849e-006, 1.616776e-007, 7.733704e-007, 7.240724e-007, 
    1.794349e-007, -3.355244e-007, -1.45038e-007, 2.627447e-006, 
    2.149864e-006, 9.216365e-007, 1.601875e-007, -1.814838e-006, 
    -7.540733e-006, -8.131812e-006, -7.887806e-006, -9.66241e-006, 
    -9.877234e-006, -8.586794e-006, -7.353103e-006, -1.852959e-006, 
    1.21879e-006, 5.566577e-006, 4.999838e-006, 4.483016e-006, 3.214304e-006, 
    2.144774e-006, 1.260638e-006, -1.188368e-006, -1.589954e-006, 
    -2.39859e-006, -1.825889e-006, -3.38989e-006, -2.527733e-006, 
    -2.939875e-006, -2.675753e-006, -2.441307e-006, -2.082934e-006, 
    -1.899153e-006, -1.516069e-006, -6.896753e-007, 2.498425e-007, 
    1.310309e-006, 1.363829e-006, 2.152845e-006, -6.047412e-008, 
    -1.055077e-005, -2.676621e-006, -1.016383e-006, -4.778306e-007, 
    -8.465101e-007, -3.285705e-007, -1.630187e-006, -3.095716e-006, 
    1.738841e-006, 8.353345e-007, 1.962111e-006, 9.570285e-007, 
    5.496058e-007, 6.571418e-007, 4.204603e-007, -4.543608e-007, 
    -1.68408e-006, -1.250953e-006,
  -2.244239e-006, -1.376867e-006, -1.054754e-006, 2.120933e-007, 
    2.71822e-007, 1.68259e-007, 1.54972e-007, 2.607703e-008, 7.83553e-008, 
    -8.602935e-007, -1.089026e-006, -2.955024e-006, -3.433476e-006, 
    -3.272544e-006, -2.975514e-006, -1.583869e-006, -5.734455e-007, 
    1.772121e-006, 7.459146e-006, 1.00142e-005, 6.011252e-006, 3.788991e-006, 
    5.039075e-006, 2.938757e-006, 3.809728e-007, 2.601493e-006, 
    1.524388e-006, 2.253056e-006, 4.762412e-006, 5.775318e-006, 
    6.056453e-006, 2.868598e-006, 3.394857e-006, 2.33377e-006, 3.481905e-006, 
    2.901877e-006, 3.283346e-006, 1.490985e-006, -8.637708e-007, 
    7.633134e-007, 2.966572e-007, 5.258869e-006, 6.386637e-006, 
    7.943563e-007, -1.879533e-006, -1.618229e-005, -1.812155e-005, 
    -1.484317e-005, -1.553595e-005, -1.720128e-005, -1.182383e-005, 
    -3.6786e-006, 3.873061e-006, 8.052586e-006, 1.122455e-005, 1.138697e-005, 
    7.846951e-006, 3.290301e-006, 4.200883e-007, -6.085884e-007, 
    -2.269695e-006, -1.921256e-006, -1.44653e-006, -1.626586e-006, 
    -1.78044e-006, -2.175818e-006, -2.60075e-006, -2.053752e-006, 
    -2.420818e-006, -1.672407e-006, -1.831725e-006, -9.288392e-007, 
    -1.122057e-006, 1.216307e-006, 2.130369e-006, 6.862481e-006, 
    -5.050995e-006, -5.994861e-006, -7.852911e-007, -1.210347e-006, 
    -5.272528e-007, -4.65413e-007, -4.778306e-007, -1.894931e-007, 
    -2.45745e-007, 4.023332e-008, 1.430262e-006, 2.117083e-006, 
    1.184146e-006, 2.707038e-007, 2.168117e-007, 1.028056e-006, 
    9.951491e-007, -2.148871e-006, -2.124533e-006, -2.281119e-006,
  -1.712888e-006, -8.153415e-007, -1.507998e-006, -1.112621e-007, 
    6.263454e-007, 1.559158e-006, 7.535018e-007, 7.214658e-008, 1.58449e-007, 
    -4.849086e-007, -1.46913e-006, -3.462409e-006, -2.636512e-006, 
    -2.209594e-006, -3.803645e-006, -5.936994e-006, -3.654013e-006, 
    -1.609198e-006, 6.500632e-007, 1.827502e-006, -1.160181e-006, 
    -1.238041e-006, 2.308065e-006, 5.323564e-006, 1.036388e-005, 
    8.373461e-006, 8.631747e-006, 9.935473e-006, 4.460414e-006, 7.32541e-006, 
    7.292629e-006, 1.682092e-006, 1.923616e-006, 3.469114e-006, 
    2.762799e-006, 4.60185e-006, 2.021789e-005, 1.15931e-005, -8.141495e-006, 
    -4.849955e-006, -1.646204e-006, -2.006818e-006, -1.480939e-005, 
    -1.765701e-005, -1.140821e-005, -2.165673e-005, -1.614355e-005, 
    -1.276608e-005, -8.465067e-007, 5.767994e-006, 1.542233e-005, 
    1.81963e-005, 2.427846e-005, 2.036566e-005, 1.504235e-005, 1.103456e-005, 
    4.837166e-006, 1.705936e-006, -7.83677e-007, -1.400957e-006, 
    -1.698981e-006, -1.33204e-006, -2.315267e-006, -2.059713e-006, 
    -2.632166e-006, -1.935537e-006, -1.802172e-006, -1.632546e-006, 
    -1.683583e-006, -1.816203e-006, -1.580765e-006, -1.376122e-006, 
    4.488975e-007, 1.90114e-007, 1.597901e-006, 6.166969e-006, 
    -3.480664e-007, 6.309401e-007, 4.111851e-006, 7.335098e-007, 
    6.705523e-008, -1.000489e-006, -5.642573e-007, -6.946424e-007, 
    -9.446094e-007, -5.37932e-007, -3.211198e-007, -1.201033e-006, 
    -5.446373e-007, 1.180048e-006, 2.388531e-006, 5.04367e-006, 
    5.068382e-006, -2.718216e-007, -1.784539e-006, -2.243743e-006,
  1.270572e-006, 3.981095e-007, 1.062329e-006, 1.597405e-006, 3.226846e-006, 
    7.819011e-006, 1.039815e-005, 5.702426e-006, 3.542131e-006, 
    2.690032e-006, 1.402696e-006, -1.179924e-006, -3.390139e-006, 
    -3.349284e-006, -6.481384e-006, -9.34874e-006, -8.451068e-006, 
    -4.678095e-006, -4.521633e-006, 5.510956e-007, 4.862002e-006, 
    5.848582e-006, 8.481118e-006, 9.631367e-006, 1.742728e-005, 
    1.309849e-005, 1.473402e-005, 9.683272e-006, 7.086246e-006, 
    1.414282e-005, 9.979308e-006, 1.488228e-005, 1.619504e-006, 
    6.053222e-006, 1.399368e-005, 4.961465e-006, 1.164898e-005, 
    -4.034613e-006, -7.553772e-006, 1.928958e-006, 1.420441e-005, 
    2.471977e-006, -9.549534e-006, 5.461523e-006, 2.211394e-005, 
    2.636301e-005, 2.915313e-005, 3.053211e-005, 3.368656e-005, 
    3.426969e-005, 3.127183e-005, 2.562938e-005, 1.769314e-005, 
    9.289135e-006, 4.842009e-006, 1.024455e-006, 1.132489e-007, 
    -8.263933e-007, -1.434609e-006, -1.676505e-006, -9.554128e-007, 
    -1.115103e-006, -1.37339e-006, -1.289944e-006, -1.40965e-006, 
    -1.183152e-006, -1.347065e-006, -1.289944e-006, -1.042585e-006, 
    -9.526807e-007, -5.486113e-007, 2.472348e-007, 1.654525e-006, 
    2.675752e-006, 2.894558e-007, 3.911182e-006, 2.454966e-006, 
    4.833069e-006, 9.209787e-006, 4.099682e-006, 2.275408e-006, 
    -1.384317e-006, -3.176307e-006, -2.737716e-006, -1.462673e-006, 
    -2.859036e-006, -7.90904e-006, -5.913278e-006, 5.779912e-006, 
    1.083898e-005, 1.501913e-005, 1.929912e-005, 1.779075e-005, 9.44386e-006, 
    4.945323e-006, 2.578397e-006,
  1.540681e-005, 1.502161e-005, 1.27852e-005, 1.314891e-005, 1.088207e-005, 
    1.220455e-005, 4.881498e-006, 3.306937e-006, 6.188449e-006, 
    1.122207e-005, 2.595534e-006, -1.688053e-006, -1.308695e-006, 
    -3.380204e-006, -4.738569e-006, -4.623209e-006, -2.132852e-006, 
    2.731758e-008, 5.134643e-007, 1.252687e-006, 3.216664e-006, 6.79717e-006, 
    1.290727e-005, 1.088605e-005, 1.272162e-005, 5.838396e-006, 
    8.792056e-006, 8.547431e-006, 1.728224e-005, 2.153416e-005, 
    1.138933e-005, 2.221999e-005, 6.172777e-007, 4.993999e-006, 
    1.259371e-005, 8.432318e-006, 7.848321e-006, -4.791094e-006, 
    -1.825269e-006, 1.413164e-005, 4.027781e-006, -1.367182e-006, 
    2.412242e-006, 1.4098e-005, 3.401762e-005, 4.993279e-005, 6.156565e-005, 
    6.777645e-005, 6.118081e-005, 5.654432e-005, 4.186928e-005, 
    3.174009e-005, 2.233461e-005, 1.305764e-005, 7.344534e-006, 
    1.829862e-006, 1.169617e-006, 5.111099e-007, 1.188369e-007, 
    -3.440925e-007, -5.173185e-007, -7.426988e-007, -7.376075e-007, 
    -1.072387e-006, -1.004835e-006, -6.118166e-007, -4.61067e-007, 
    -3.932664e-007, -6.072241e-008, 1.52861e-007, 1.771252e-006, 
    3.495936e-006, 6.05161e-006, 1.240224e-005, 4.127622e-006, 
    -2.302848e-006, 2.102552e-006, 5.391114e-006, 1.951033e-005, 
    2.045346e-005, 8.386851e-007, -3.405163e-006, -9.913493e-006, 
    -1.248357e-005, -1.034898e-005, -1.934891e-005, -2.407419e-005, 
    4.52486e-006, 2.195872e-005, 2.569556e-005, 2.867294e-005, 2.8382e-005, 
    2.583129e-005, 1.817222e-005, 1.570632e-005, 1.242198e-005,
  1.130638e-005, 2.031799e-005, 1.134388e-005, 1.87284e-005, 1.42516e-005, 
    3.227964e-006, -4.236397e-006, -6.142262e-006, 5.188085e-006, 
    8.015704e-006, -4.946189e-006, -1.854698e-006, -3.992268e-007, 
    -2.206117e-006, -2.237906e-006, 1.756223e-006, 4.961345e-006, 
    2.439694e-006, 3.429006e-006, 2.776091e-006, 8.459887e-006, 
    5.273396e-006, 8.084506e-006, 1.380468e-005, 1.694101e-005, 
    9.455282e-006, 3.164634e-006, 9.160241e-006, 1.919779e-005, 2.45663e-005, 
    9.407602e-006, 7.60195e-006, 1.311886e-005, 5.415583e-006, 1.057859e-006, 
    3.401685e-006, 4.109366e-006, 5.643815e-007, 5.551847e-007, 
    -1.050669e-005, -7.028386e-006, -1.798211e-005, 1.207367e-005, 
    4.173381e-005, 3.520822e-005, 3.305624e-005, 2.766339e-005, 
    3.211287e-005, 2.992091e-005, 2.94303e-005, 3.155731e-005, 2.660044e-005, 
    3.048914e-005, 3.036782e-005, 2.398764e-005, 1.866544e-005, 
    1.609934e-005, 8.663908e-006, 5.949161e-006, 4.909685e-006, 
    3.986557e-006, 6.710243e-006, 7.374832e-006, 6.255383e-006, 
    6.880984e-006, 8.38712e-006, 1.433802e-005, 1.4661e-005, 1.391173e-005, 
    2.197201e-005, 1.331668e-005, -8.769348e-007, -3.499168e-006, 
    9.554875e-006, 1.527194e-005, -1.422875e-005, -2.51086e-007, 
    5.665919e-006, 8.389979e-006, -6.309405e-006, -3.315259e-006, 
    -5.151331e-006, -1.909335e-006, -5.974991e-006, -2.109061e-005, 
    -7.644296e-006, -1.070475e-005, -2.109009e-006, 1.548244e-005, 
    1.06583e-005, 1.407639e-005, 6.073475e-006, -3.161651e-006, 
    9.993746e-007, 4.155307e-006, 2.07503e-007,
  -4.892354e-008, 3.67537e-006, 6.770715e-006, 1.457644e-005, -4.018293e-007, 
    -8.409224e-006, -8.893257e-006, -5.265327e-006, -6.345537e-006, 
    -5.606809e-006, -2.662788e-005, 1.206619e-006, -5.152078e-007, 
    3.452101e-008, -2.941738e-007, 5.123516e-006, 1.328935e-005, 
    1.081601e-005, 1.176111e-005, 1.377426e-005, 5.13556e-006, 1.45665e-005, 
    1.2984e-005, 7.787472e-006, 2.704932e-006, 7.951756e-006, 8.119016e-006, 
    1.319609e-005, 2.269336e-005, 2.303396e-005, 1.247227e-005, 
    2.617438e-005, 1.67371e-005, 4.907488e-007, -5.253038e-006, 
    -6.543996e-008, 2.987435e-006, -3.201021e-006, -5.148475e-006, 
    -1.105157e-005, 7.909417e-006, 4.815935e-006, 2.606498e-005, 
    3.702628e-005, 2.435421e-005, 1.615187e-005, 1.470682e-005, 1.45295e-005, 
    1.398523e-005, 1.091015e-006, -6.03497e-006, -8.426483e-006, 
    -1.635031e-006, 3.325942e-006, -3.43733e-006, -4.125177e-007, 
    -7.75115e-007, 1.271816e-006, 1.850276e-008, -1.093894e-005, 
    -4.064292e-006, 1.275279e-005, 1.582479e-005, -2.387416e-006, 
    1.109715e-005, 1.225242e-006, 7.513911e-006, 1.134252e-005, 
    6.078932e-006, -7.358074e-006, -1.842964e-005, -8.150688e-006, 
    -3.49262e-005, -5.427661e-005, -3.447607e-005, -1.740654e-005, 
    -8.446223e-006, -1.294563e-005, -1.293185e-005, -9.888907e-006, 
    -7.9448e-006, -8.127217e-006, -2.686182e-006, -5.096321e-006, 
    -6.834543e-006, 2.135956e-006, -5.132704e-006, -3.141537e-006, 
    -3.035366e-006, -8.110583e-006, -8.659932e-006, -1.300077e-005, 
    -2.242476e-005, -2.003796e-005, -1.100277e-005, -7.695198e-007,
  -2.582892e-007, 5.498281e-006, 1.046372e-005, 1.367318e-005, 9.621428e-006, 
    1.084307e-006, -8.444611e-006, -1.02022e-005, -2.737339e-006, 
    2.11125e-006, -9.402258e-006, -8.447591e-006, -1.629069e-006, 
    -1.140808e-006, -2.818804e-007, -4.085405e-008, 6.000822e-006, 
    1.30775e-005, 1.195831e-005, 8.106232e-006, 5.087626e-006, 1.639302e-005, 
    1.883594e-005, 1.09495e-005, -6.645925e-006, 1.199741e-005, 
    3.323717e-005, 3.091407e-005, 3.98395e-005, 3.341176e-005, 2.708609e-005, 
    3.766801e-005, 1.729267e-005, 1.04061e-005, 1.041466e-006, 
    -1.361346e-005, -4.590678e-006, -1.232205e-006, -2.187859e-006, 
    -3.478919e-006, 1.340049e-005, 1.359954e-005, 2.160308e-005, 
    1.462115e-005, 1.031297e-005, 1.40698e-005, 1.209739e-005, 1.36435e-005, 
    1.310942e-005, -7.721246e-007, 1.666696e-006, 9.148316e-006, 
    3.763045e-006, -3.037225e-006, 2.803899e-006, 3.61403e-006, 6.41284e-006, 
    3.44155e-006, -5.468351e-006, 1.168624e-006, 8.259089e-006, 
    -2.051518e-006, -4.172703e-006, -9.437776e-006, 1.347435e-006, 
    -1.736356e-006, -5.962698e-006, -2.265107e-006, -5.85652e-006, 
    -1.730124e-005, -1.049961e-005, -3.386637e-005, -4.376807e-005, 
    -4.110821e-005, -1.999761e-005, -1.222591e-005, -7.277231e-006, 
    -6.042048e-006, -6.552786e-006, -1.044273e-005, -1.469192e-005, 
    -9.483596e-006, -1.199916e-005, -7.479637e-006, -5.642822e-006, 
    -6.435191e-006, -6.285807e-006, -5.494307e-006, -4.550318e-006, 
    -4.536286e-006, -4.70976e-006, -8.676947e-006, -3.669786e-006, 
    -4.445264e-006, 2.030654e-006, 3.247835e-006,
  7.496154e-006, 4.211812e-006, 3.387529e-006, 5.961955e-006, 6.48126e-006, 
    2.159054e-006, -2.223996e-007, -2.290557e-006, -1.615657e-006, 
    -2.422556e-006, -5.235648e-006, 6.919106e-007, 1.989181e-006, 
    3.247832e-006, 1.034265e-006, 1.41561e-007, -3.234793e-007, 
    2.008552e-006, 8.95212e-006, 1.259495e-005, 6.223221e-006, 1.171753e-005, 
    9.198113e-006, 5.793583e-006, 2.925706e-006, 1.156765e-005, 
    1.696497e-005, 1.830695e-005, 1.888399e-005, 2.669767e-005, 
    -9.293726e-006, 8.525079e-006, -1.009282e-005, 7.13468e-006, 
    1.280889e-006, -8.415431e-006, -6.816037e-006, 4.493071e-006, 
    1.268858e-005, 9.094052e-006, 1.709511e-005, 8.493902e-006, 
    1.318082e-005, 7.622191e-006, 1.18232e-005, -9.519354e-007, 
    2.569948e-006, 6.527829e-006, 6.593764e-006, 3.835186e-006, 
    2.937391e-006, 2.951674e-007, -3.717345e-006, -3.147248e-006, 
    -1.969313e-006, -2.231822e-006, -4.080062e-006, -8.037314e-006, 
    -7.442757e-006, -3.468867e-006, -3.036981e-006, -7.275865e-006, 
    -6.354972e-006, -4.091486e-006, -2.747649e-006, 2.781177e-006, 
    1.14236e-005, 9.889896e-006, 1.429928e-005, 3.562993e-006, 
    -1.903139e-005, -4.249935e-005, -3.149062e-005, -2.148363e-005, 
    -9.523705e-006, -8.199735e-006, -6.034101e-006, -7.164726e-006, 
    -9.273985e-006, -9.073317e-006, -8.351604e-006, -8.377061e-006, 
    -5.914891e-006, -4.046286e-006, -3.857538e-006, -2.752866e-006, 
    -2.632911e-006, -2.586469e-006, -2.445778e-006, -1.596659e-006, 
    -1.777957e-006, -2.387042e-006, -8.049979e-006, -7.689745e-006, 
    2.192086e-006, 6.790586e-006,
  1.026442e-006, 2.780312e-007, 5.478661e-007, 4.193435e-007, 7.862846e-007, 
    9.97757e-007, 5.16822e-007, 1.077478e-006, 1.099954e-006, 1.55891e-006, 
    -2.796824e-006, 2.191713e-007, 2.559274e-007, 3.216291e-006, 
    3.313646e-006, 1.262625e-006, 1.690164e-006, 3.055483e-006, 
    5.284325e-006, 2.285714e-005, 2.295984e-005, 2.119889e-005, 9.92306e-006, 
    -1.968445e-006, 6.848451e-006, 9.622177e-006, 8.509305e-006, 
    1.095534e-005, -3.135945e-006, 1.637141e-006, -7.626775e-006, 
    1.21098e-005, -7.472554e-006, -1.591667e-005, -5.418689e-006, 
    -4.596761e-006, -1.147389e-006, 1.554191e-005, 2.361846e-005, 
    2.721101e-005, 2.459063e-005, 9.794283e-006, 2.038112e-006, 
    3.192617e-007, -6.345035e-006, -1.652661e-006, -1.426415e-006, 
    -1.198823e-005, -1.557407e-005, -1.002091e-005, -7.272261e-006, 
    -7.503604e-006, -3.850955e-006, -1.872952e-006, -1.679859e-006, 
    -3.783662e-007, -5.467485e-006, -6.987403e-006, -5.054349e-006, 
    -4.347414e-006, -3.270432e-006, -2.782171e-006, -2.486259e-006, 
    -1.541152e-006, -1.2815e-006, -4.34816e-006, -1.733427e-005, 
    2.825262e-006, -6.65088e-007, -3.376615e-005, -1.99544e-005, 
    -1.452752e-005, -5.086139e-006, -9.656946e-006, -1.771437e-005, 
    -1.356155e-005, -1.355323e-005, -9.139254e-006, -8.172667e-006, 
    -8.097912e-006, -8.835147e-006, -5.024547e-006, -2.560268e-006, 
    -2.090384e-006, -1.525134e-006, -1.293172e-006, -1.746416e-006, 
    -1.182655e-006, -1.455471e-006, -9.669611e-007, -7.092954e-007, 
    -4.333755e-007, -2.1182e-006, -4.389385e-006, -1.906355e-006, 
    9.059904e-007,
  5.292395e-007, -8.02055e-007, -2.520781e-007, -8.891026e-008, 
    -2.99265e-008, -4.457931e-008, -1.937151e-008, -2.011657e-008, 
    7.947285e-009, 1.033147e-007, 4.433096e-008, 7.972123e-008, 
    1.318753e-007, 1.904492e-006, 3.21058e-006, 3.951664e-006, 1.971374e-005, 
    1.32747e-005, 1.097557e-005, 1.628784e-005, 1.478717e-005, 6.814054e-006, 
    6.799026e-006, 6.472816e-006, 2.058099e-006, 2.78902e-007, 1.210061e-005, 
    4.937247e-007, 6.220944e-008, 1.523273e-006, 5.515292e-006, 
    2.350287e-006, 2.315763e-006, -1.427288e-006, 1.985536e-007, 
    6.248556e-006, 2.66383e-006, 6.188326e-006, 1.206112e-005, 1.043094e-005, 
    9.174888e-006, 1.454355e-006, -4.474321e-006, -6.189315e-006, 
    -7.564326e-006, -2.176566e-006, -2.743051e-006, -6.859376e-006, 
    -1.331779e-005, -1.063136e-005, -1.488986e-005, -1.577151e-005, 
    -9.362275e-006, -2.70543e-006, -2.064557e-006, -4.49419e-006, 
    -2.201895e-006, -3.665189e-006, -3.871446e-006, -1.805151e-006, 
    -1.80838e-006, -2.104665e-006, -2.015381e-007, -9.586415e-008, 
    -6.075948e-007, 3.892928e-007, -1.270957e-005, -1.376234e-005, 
    -1.142807e-005, -3.327801e-006, -1.156077e-007, -7.427981e-006, 
    -5.679576e-006, -7.56482e-006, -8.26679e-006, -3.949302e-006, 
    -6.086626e-006, -3.055109e-006, -6.673983e-006, -8.186822e-006, 
    -6.295367e-006, -3.765275e-006, -1.674643e-006, -4.96706e-007, 
    -5.447619e-007, -8.482493e-007, -9.725491e-007, -1.318132e-006, 
    -1.427407e-006, -1.396736e-006, -1.314903e-006, -7.029623e-007, 
    -1.038114e-006, -1.146272e-006, -8.477521e-007, 3.018727e-007,
  -2.120932e-007, 3.474454e-007, 2.055119e-007, 1.69004e-007, -4.993131e-007, 
    -3.357729e-007, -8.990367e-008, -2.880891e-008, -1.812975e-008, 
    -4.967053e-010, 5.30233e-008, 1.642853e-007, 9.660919e-008, 
    1.105169e-008, 1.396984e-007, 1.556302e-006, 2.790491e-006, 
    2.303471e-006, 1.189522e-005, 1.517832e-005, 1.459755e-005, 
    1.392203e-005, 1.273639e-005, 1.748887e-005, 2.989909e-006, 
    6.348266e-006, 3.108146e-005, 1.136884e-005, -4.842877e-008, 
    -9.462237e-007, -1.988436e-006, -3.827859e-006, -4.818066e-007, 
    6.431714e-006, 2.499422e-006, 1.449385e-006, 4.434336e-006, 
    7.809824e-006, 4.815807e-006, 7.020932e-006, 1.413512e-005, 
    3.318117e-006, -2.293909e-006, -8.239473e-006, -1.394874e-006, 
    3.806377e-006, 4.630787e-006, -2.596535e-007, -5.986542e-006, 
    -9.073565e-006, -8.390471e-006, -1.262948e-005, -9.963785e-006, 
    -8.928146e-008, 2.007928e-007, 2.893285e-008, -3.829475e-006, 
    -4.152209e-006, -2.299125e-006, -1.575425e-006, -8.549541e-007, 
    -1.634161e-006, -2.169363e-007, 5.030383e-007, -8.245343e-008, 
    -1.555309e-006, -7.516766e-006, -9.153908e-006, 2.565359e-006, 
    4.280483e-006, 8.465226e-006, 7.122762e-007, 4.649657e-006, 
    5.126498e-006, -2.81657e-006, -7.339815e-006, -8.641557e-006, 
    -4.846603e-006, -4.141653e-006, -8.080031e-006, -8.51949e-006, 
    -6.006782e-006, -1.806393e-006, -1.087908e-006, -1.143788e-006, 
    -3.09944e-007, -1.05556e-008, -1.3041e-006, -1.657754e-006, 
    -1.17893e-006, -1.672779e-006, 5.451329e-008, -2.955396e-007, 
    -1.17359e-006, -1.2363e-006, -3.0001e-007,
  -3.282602e-006, -2.465894e-006, -1.813099e-006, -8.353343e-007, 
    -7.04204e-007, -7.222097e-007, -2.474835e-007, -7.947286e-008, 
    -1.130005e-007, -1.498809e-007, -4.470344e-009, 3.700455e-008, 
    3.259913e-023, 7.450573e-010, 3.526608e-007, 4.464139e-007, 
    1.270324e-007, 1.385808e-007, 1.627827e-006, 5.494308e-006, 
    5.381306e-006, 1.465889e-005, 3.84028e-006, 3.80762e-006, 5.983187e-006, 
    1.403503e-005, 3.348167e-005, 5.761423e-006, 4.357717e-006, 
    2.017245e-006, 2.12677e-006, 2.859408e-006, 2.300738e-006, 2.755225e-006, 
    6.816412e-006, 3.803398e-006, 2.991907e-006, -2.421439e-006, 
    3.132594e-006, 3.290799e-006, 9.742751e-006, 2.049779e-006, 
    1.145527e-006, 1.404558e-006, 6.042297e-006, 1.173926e-005, 
    8.441757e-006, 5.635247e-006, 1.649933e-006, -4.821146e-006, 
    -2.465895e-006, -7.450581e-008, -4.267931e-007, -3.448501e-006, 
    -7.631879e-007, 2.703318e-007, -4.121421e-007, -9.529285e-007, 
    -6.948903e-007, -1.634781e-006, -8.232892e-007, -2.458683e-008, 
    9.309499e-007, 1.561642e-006, -4.333754e-007, -2.987186e-006, 
    -5.818159e-006, -2.58175e-006, 5.517776e-006, 3.882498e-006, 
    7.238114e-006, 5.215778e-006, 8.751949e-007, 6.968785e-007, 
    1.730397e-006, 1.483932e-007, -6.582588e-006, -7.639326e-006, 
    -6.850685e-006, -7.411712e-006, -7.297594e-006, -7.817522e-006, 
    -5.954505e-006, -2.891321e-006, -1.402447e-006, -1.123547e-006, 
    -4.978228e-007, -1.096104e-006, -9.2561e-007, -1.859044e-006, 
    -1.174584e-006, -8.648881e-007, 1.023462e-006, -4.863987e-007, 
    -9.66092e-007, -3.550574e-006,
  -5.313258e-006, -5.730862e-006, -6.317471e-006, -4.312396e-006, 
    -1.989677e-006, -1.089399e-006, -9.858359e-007, -7.521361e-007, 
    -1.73226e-006, -7.869055e-007, 1.117588e-009, 1.862645e-009, 
    -4.731119e-008, -7.015967e-008, 2.563e-007, 8.50608e-008, 6.842117e-008, 
    3.961225e-008, -5.566826e-007, -1.350666e-006, 5.281219e-007, 
    2.001349e-006, 2.170354e-006, 3.284588e-006, 2.64918e-006, 3.189594e-006, 
    1.882509e-007, -1.0591e-005, -2.513829e-006, 4.940477e-006, 
    1.570533e-005, 1.245638e-005, 6.551671e-006, 6.327282e-006, 
    9.943795e-006, 8.985277e-006, 7.227187e-006, 4.271293e-006, 
    1.015862e-005, 9.348614e-006, 1.182606e-005, 6.107861e-006, 
    -4.929825e-008, 8.592997e-007, -1.674518e-006, 2.517923e-006, 
    6.051238e-006, 6.15865e-006, 2.073739e-007, -4.630547e-007, 
    -1.521166e-007, 2.077843e-006, 1.438708e-006, -1.490241e-006, 
    -4.487738e-007, 6.66827e-007, -1.22438e-007, -9.164214e-007, 
    -1.267592e-006, -1.139318e-006, -9.090945e-007, -1.378385e-008, 
    2.411505e-007, 1.029422e-007, 8.034209e-008, -1.165147e-006, 
    -1.533578e-006, -1.016258e-006, 2.530714e-007, 3.621479e-006, 
    7.678693e-006, 5.538264e-006, 2.342835e-006, 4.608433e-006, 
    1.129496e-005, 1.042386e-005, 7.465107e-006, -1.101071e-006, 
    -4.433594e-006, -6.593389e-006, -5.942584e-006, -5.873047e-006, 
    -6.747245e-006, -4.200514e-006, -3.305325e-006, -2.16576e-006, 
    6.762639e-007, -7.325166e-007, -1.531342e-006, -1.576791e-006, 
    -6.991127e-007, -1.026814e-006, 2.179295e-007, 9.513149e-007, 
    -8.769334e-007, -2.89691e-006,
  -2.979612e-006, -1.59579e-006, 2.935531e-007, -2.86971e-007, 
    -2.435098e-006, -3.069267e-006, -2.720704e-006, -1.189609e-006, 
    -1.931935e-006, -1.31391e-006, -3.064672e-007, -1.773237e-007, 
    -6.771336e-007, -6.765129e-007, -2.910693e-007, 1.291434e-007, 
    -2.644958e-008, 5.923211e-008, 4.271666e-008, -9.972601e-007, 
    -1.60262e-006, 1.858921e-007, 6.704281e-007, 8.780512e-007, 
    -5.509701e-007, -4.284084e-007, -4.839399e-006, -1.735973e-005, 
    -1.191186e-005, -4.701316e-006, -4.600981e-006, 3.139052e-006, 
    1.016185e-005, 9.126466e-006, 1.91917e-005, 1.556004e-005, 6.300957e-006, 
    8.864328e-006, 1.791989e-005, 1.790424e-005, 1.52157e-005, 1.223335e-005, 
    7.633493e-006, 3.108506e-006, -1.105163e-007, 1.932185e-007, 
    1.851717e-006, 2.321725e-006, 9.570285e-007, 8.687384e-007, 
    1.426779e-007, -5.832571e-007, 1.214941e-006, -9.58642e-007, 
    2.122173e-006, 7.4543e-007, -4.061812e-007, -1.214941e-006, 
    -1.938517e-006, -1.252194e-006, -1.188492e-006, -7.381041e-007, 
    -1.701216e-007, -1.054257e-007, 3.187606e-007, -5.493562e-007, 
    -1.37873e-006, -1.049911e-006, 1.408036e-006, 7.049865e-006, 
    9.976451e-006, 9.363393e-006, 4.400063e-006, 4.252295e-006, 
    5.339334e-006, 6.122889e-006, 6.326536e-006, 5.179147e-006, 
    1.150616e-006, -4.015365e-006, -6.245573e-006, -6.877879e-006, 
    -3.624955e-006, -8.347124e-007, -1.954162e-006, -5.712112e-006, 
    -3.554548e-006, -7.491553e-007, -6.999817e-007, -1.196811e-006, 
    -1.401454e-006, -1.639128e-006, -1.650552e-006, -8.008133e-007, 
    -9.718041e-007, -8.877369e-007,
  -5.28271e-006, -2.515937e-006, -2.124657e-006, -2.159799e-006, 
    -3.565476e-006, -5.910918e-006, -7.20496e-006, -2.518048e-006, 
    -2.840286e-006, -2.751996e-006, -3.373002e-006, -5.901107e-006, 
    -2.384186e-006, 3.387531e-007, 1.423806e-006, 1.301244e-006, 
    1.223634e-006, 1.405677e-007, -8.121131e-008, -2.207855e-007, 
    -5.010515e-007, -4.548583e-007, -9.747828e-008, 2.991408e-007, 
    -1.362214e-007, -3.664445e-007, 2.359352e-007, -2.748769e-006, 
    -2.882505e-006, -3.09994e-006, -3.701945e-006, -7.821123e-006, 
    -7.800136e-006, -2.642351e-006, 4.69424e-006, 1.007244e-005, 
    8.470193e-006, 6.685532e-006, 3.415222e-006, 1.202846e-005, 
    1.490315e-005, 1.861466e-005, 1.523706e-005, 1.480282e-005, 1.04893e-005, 
    3.446516e-006, 2.351029e-006, 3.169105e-006, 2.939127e-006, 
    2.131987e-006, 4.487854e-006, 3.409881e-006, -4.476569e-007, 
    2.853323e-006, 4.807114e-006, 3.886098e-006, 1.008933e-006, 
    -5.898373e-007, -1.123672e-006, -1.92523e-006, -1.746292e-006, 
    -7.413328e-007, -1.112744e-006, -5.30978e-007, 4.950912e-007, 
    2.272179e-006, 1.834333e-006, 3.387035e-006, 8.961435e-006, 
    7.793305e-006, 5.233289e-006, 3.884485e-006, 2.318e-006, 1.644716e-006, 
    1.671413e-006, 3.155568e-006, 2.462417e-006, -2.898896e-006, 
    -6.45034e-006, -7.852042e-006, -9.446094e-006, -9.445101e-006, 
    -9.03271e-006, -7.820378e-006, -5.333375e-006, -3.895038e-006, 
    -3.914287e-006, -2.848854e-006, -1.523147e-006, -1.983345e-006, 
    -2.373383e-006, -9.605037e-007, -1.899401e-006, -3.188104e-006, 
    -2.042329e-006, -9.297082e-007,
  -7.275739e-006, -5.668154e-006, -9.887666e-006, -6.201863e-006, 
    -1.720959e-006, -4.115702e-006, -3.205862e-006, -2.549837e-006, 
    -3.559763e-006, -4.002824e-006, -2.820045e-006, -3.121172e-006, 
    -2.45894e-006, 6.606206e-008, 1.464536e-006, 1.145154e-006, 1.11945e-006, 
    1.502782e-006, 4.849087e-007, -7.388496e-008, -3.694247e-007, 
    -6.135554e-007, -8.265179e-007, -6.556547e-008, 2.291054e-007, 
    8.357074e-008, -9.696932e-007, -2.776578e-007, -1.349799e-007, 
    -5.44389e-007, -5.654983e-007, 7.23081e-007, -4.808851e-006, 
    -3.469115e-006, 1.357257e-007, 4.645808e-006, 6.162998e-006, 
    3.862257e-006, 3.594534e-006, 3.569075e-006, 3.685054e-006, 
    6.978462e-006, 7.396688e-006, 5.276004e-006, 6.190563e-006, 
    4.003818e-006, 3.145633e-006, 5.597001e-006, 4.774953e-006, 
    3.608689e-006, 4.654878e-006, 4.379326e-006, 5.295624e-006, 
    5.517282e-006, 4.058829e-006, 3.957997e-006, 3.431613e-006, 
    1.705439e-006, 2.102306e-006, 1.311054e-006, -3.593668e-007, 
    -6.253522e-007, -4.374733e-007, -7.974604e-007, -1.587843e-006, 
    -1.87134e-007, 2.356246e-006, 4.342075e-006, 7.448967e-006, 
    4.190581e-006, 2.341345e-006, 7.105355e-007, -2.259016e-006, 
    -3.057843e-006, -2.518047e-006, -2.174329e-007, -1.932203e-007, 
    -4.19778e-006, -4.899997e-006, -6.936491e-006, -7.846207e-006, 
    -6.326536e-006, -5.637108e-006, -6.121023e-006, -7.507204e-006, 
    -4.608059e-006, -2.047047e-006, -1.317883e-006, -4.830454e-007, 
    -1.12007e-006, -2.111618e-006, -4.686417e-007, -3.634641e-007, 
    -1.858423e-006, -1.200165e-006, -3.54958e-006,
  -4.314879e-006, -8.578847e-006, -9.452673e-006, -9.655923e-007, 
    2.71524e-006, -6.680784e-008, -1.7073e-006, -2.677366e-006, 
    -1.708791e-006, -3.125022e-006, -2.464031e-006, -1.685196e-006, 
    1.654025e-007, 2.312412e-006, 4.074226e-006, 2.519414e-006, 
    1.483038e-006, 1.552577e-006, 4.726148e-007, -8.999059e-007, 
    -5.622705e-007, -6.083396e-007, -4.068015e-007, -1.681224e-006, 
    -1.422936e-006, -9.926662e-007, 8.256484e-007, 3.860519e-006, 
    3.253794e-006, -9.443611e-007, 6.165355e-007, 5.926922e-007, 
    3.987923e-006, 3.406531e-006, 4.258627e-006, 8.949268e-006, 
    1.017812e-005, 4.693993e-006, 4.878144e-006, 3.662954e-006, 
    -2.282359e-007, -2.804027e-006, 1.97229e-006, 3.317618e-006, 
    3.197041e-006, 2.014265e-006, 2.032521e-006, 2.398341e-006, 
    4.646929e-006, 3.275025e-006, 2.49048e-006, 3.797435e-006, 4.344929e-006, 
    5.83666e-006, 4.985806e-006, 1.73698e-006, 1.125038e-006, -4.98816e-007, 
    5.795318e-007, 7.227063e-007, -2.806373e-007, -4.990634e-007, 
    -2.976522e-007, -3.808116e-006, -5.094831e-006, -3.001715e-006, 
    -1.694883e-006, -1.400957e-006, 8.15342e-007, -3.909081e-007, 
    -7.910021e-007, 1.803055e-007, 3.481282e-006, 3.020339e-006, 
    2.499175e-006, 2.592787e-007, -1.288827e-006, -1.671415e-006, 
    -5.31847e-007, -3.511585e-006, -2.538662e-006, 3.430247e-006, 
    2.809244e-006, -1.949593e-008, -9.395189e-007, -3.719702e-006, 
    -6.239861e-007, 2.021588e-007, 1.596905e-006, 3.034875e-007, 
    9.352952e-007, 5.780421e-007, -5.351994e-007, -2.504621e-007, 
    3.671894e-007, -2.056237e-006,
  -2.821907e-006, -2.106404e-006, -1.506383e-006, -2.610177e-007, 
    -1.721073e-007, -5.114834e-007, 1.817445e-006, 3.378962e-006, 
    4.423286e-006, 2.400204e-006, 2.753859e-006, 1.436099e-006, 
    1.118829e-006, 2.374873e-006, 4.338845e-006, 4.475689e-006, 
    3.240382e-006, 3.15259e-006, 2.284223e-006, 1.193086e-006, 6.869432e-007, 
    1.495082e-007, 9.571522e-007, 5.751845e-007, 4.58087e-007, 2.319613e-006, 
    3.85195e-006, 2.981349e-006, 1.746168e-006, 1.158565e-006, 3.886844e-006, 
    5.356844e-006, 4.183377e-006, 3.108256e-006, 6.053473e-006, 
    6.784125e-006, 3.278255e-006, 4.153451e-006, 5.468602e-006, 
    3.345809e-006, -7.549897e-008, -2.511713e-006, 1.588214e-006, 
    6.525468e-006, 7.136912e-006, 5.046031e-006, 2.909699e-006, 
    4.394105e-006, 4.714477e-006, 3.425283e-006, 5.695947e-007, 
    2.143286e-006, 4.681322e-006, 7.262079e-006, 7.441142e-006, 
    2.749141e-006, 1.915545e-006, 2.114599e-006, 1.395867e-006, 
    2.353885e-006, 2.275656e-006, 4.560501e-006, 6.881975e-006, 
    5.166854e-006, -7.612107e-008, -1.422937e-006, -1.818313e-006, 
    -3.659972e-006, -2.781426e-006, -6.864466e-007, -2.684319e-006, 
    -2.586345e-006, 1.934171e-006, 5.00406e-006, 3.227964e-006, 
    2.950927e-006, 3.178542e-006, 5.706024e-006, 5.06391e-006, 3.473833e-006, 
    3.056102e-006, 3.398334e-006, 6.460647e-006, 8.236368e-006, 
    8.221345e-006, 5.43557e-006, 1.235803e-006, -1.03948e-006, 
    -3.842033e-007, 9.586402e-007, 1.483906e-006, 2.305955e-006, 
    2.364441e-006, 1.976763e-006, 2.819796e-006, 4.147478e-008,
  5.977854e-007, 1.249462e-006, -1.496448e-006, -3.076964e-006, 
    -2.887349e-006, 4.366048e-007, 2.85295e-006, 3.819663e-006, 
    4.363184e-006, 3.924843e-006, 2.931181e-006, 5.23217e-006, 7.217501e-006, 
    5.346163e-006, 4.074847e-006, 4.472087e-006, 4.041816e-006, 
    4.835551e-006, 2.951672e-006, 2.959743e-006, 3.97116e-006, 3.007551e-006, 
    2.573679e-006, 1.982599e-006, 1.022965e-006, 2.394368e-006, 
    2.376612e-006, 2.973278e-006, 3.181645e-006, 2.7402e-006, 1.764918e-006, 
    6.612143e-006, 3.188848e-006, 1.134475e-006, 1.480281e-005, 
    1.936406e-005, 3.942721e-006, -1.396611e-006, 2.007806e-006, 
    2.189976e-006, 1.731267e-006, 2.359475e-006, 4.325186e-006, 
    7.676459e-006, 5.17927e-006, 3.692383e-006, 5.574897e-006, 5.910422e-006, 
    7.295484e-006, 5.196282e-006, 3.967682e-006, 5.788852e-006, 
    6.827588e-006, 4.980217e-006, 5.66716e-006, 5.832688e-006, 3.349654e-006, 
    3.709894e-006, 1.894063e-006, 3.86437e-007, 1.77895e-006, 3.915033e-006, 
    1.687804e-006, 4.339963e-006, 4.679088e-006, 2.173459e-006, 
    1.059224e-006, 1.053761e-006, 1.718601e-006, 1.803166e-006, 
    3.175934e-006, 1.891827e-006, -7.988256e-007, 4.416943e-007, 
    1.34421e-006, 1.21606e-006, 3.395602e-006, 5.829706e-006, 9.274854e-006, 
    7.160505e-006, 6.60134e-006, 2.911313e-006, 2.880271e-006, 5.051867e-006, 
    4.041318e-006, 5.915141e-006, 4.937252e-006, 8.111201e-007, 
    -6.099544e-007, -9.29831e-007, -2.767883e-007, 3.642072e-007, 
    2.801915e-006, 5.281217e-006, 2.878656e-006, 1.865874e-006,
  1.874814e-006, 9.674586e-007, 3.085906e-006, 3.659352e-006, 3.455578e-006, 
    3.081932e-006, 3.269439e-006, 1.253313e-006, 1.306957e-006, 
    2.691522e-006, 4.66307e-006, 2.731631e-006, 3.148987e-006, 3.51034e-006, 
    2.510846e-006, 2.03152e-007, -5.677339e-007, -9.387804e-008, 
    1.571203e-006, 2.185131e-006, 2.216051e-006, 1.92138e-006, 2.903987e-006, 
    3.419693e-006, 3.66134e-006, 3.435338e-006, 4.334499e-006, 3.240259e-006, 
    3.400817e-006, 1.983966e-006, -8.073948e-007, -4.41074e-007, 
    1.691278e-007, 2.258022e-006, 4.500896e-006, 5.780284e-006, 
    6.223223e-006, 7.930646e-006, 1.140038e-005, 9.174521e-006, 
    6.614253e-006, 4.78824e-006, 3.995374e-006, 4.88721e-006, 5.535161e-006, 
    4.483387e-006, 4.617497e-006, 6.374468e-006, 7.663419e-006, 
    7.131572e-006, 3.51866e-006, 3.085037e-006, 2.300243e-006, 3.040333e-006, 
    5.299597e-006, 8.949264e-006, 9.992222e-006, 1.136288e-005, 
    8.184961e-006, 7.241841e-006, 2.253924e-006, 9.889409e-007, 
    6.029986e-007, 1.117711e-006, 1.786773e-006, 2.397721e-006, 
    2.038231e-006, 2.005323e-006, 1.024207e-006, -6.75147e-007, 
    6.465852e-007, 8.761881e-007, -1.058479e-006, -8.614115e-007, 
    9.93412e-007, 1.929948e-006, 3.315508e-006, 4.836917e-006, 5.266567e-006, 
    7.317587e-006, 5.983065e-006, 3.798803e-006, 6.667524e-006, 
    8.088848e-006, 4.95687e-006, 9.232757e-006, 1.135916e-005, 6.870803e-006, 
    2.375491e-007, -1.153101e-006, -1.375005e-006, 5.464244e-009, 
    1.838927e-006, 3.306321e-006, 4.50996e-006, 3.748262e-006,
  3.179412e-006, 2.871082e-006, 1.512964e-006, 1.486638e-006, 1.47745e-006, 
    -6.495666e-007, -2.609317e-006, -3.70419e-007, 1.628696e-006, 
    2.573679e-006, 1.772742e-006, 2.599507e-006, 3.950547e-006, 
    3.597761e-006, 3.202011e-006, 1.395245e-006, 7.015969e-007, 
    7.585932e-007, 2.337869e-006, 3.119434e-006, 2.098829e-006, 
    2.188359e-006, 2.770871e-006, 2.546236e-006, 2.712011e-006, 
    4.254653e-006, 4.633641e-006, 2.724802e-006, 1.946588e-006, 1.31006e-006, 
    1.688551e-006, 2.919385e-006, 3.04915e-006, 2.783537e-006, 2.009545e-006, 
    1.757964e-006, 2.147877e-006, 2.936769e-006, 3.815441e-006, 
    8.529176e-006, 9.654961e-006, 7.536883e-006, 6.144741e-006, 3.78862e-006, 
    4.099433e-006, 5.456061e-006, 7.139892e-006, 6.785243e-006, 
    4.995614e-006, 4.114707e-006, 2.557535e-006, 3.866975e-006, 
    5.325675e-006, 4.678343e-006, 1.554439e-006, 1.127893e-006, 
    3.116702e-006, 2.579389e-006, 1.575674e-006, 2.693881e-006, 
    4.734844e-006, 4.771848e-006, 2.332652e-006, 9.809928e-007, 
    7.306535e-007, 1.829118e-006, 3.252302e-006, 4.545227e-006, 
    4.096455e-006, 2.284349e-006, 1.936282e-006, 2.221515e-006, 
    9.395189e-007, 5.708389e-007, 1.065557e-006, 1.625469e-006, 4.75496e-006, 
    5.806362e-006, 5.23068e-006, 4.592786e-006, 3.318488e-006, 4.528089e-006, 
    8.472428e-006, 1.208124e-005, 1.04143e-005, 1.027125e-005, 1.100972e-005, 
    8.636713e-006, 5.762653e-006, 3.25938e-006, 3.920619e-006, 2.311543e-006, 
    3.787318e-008, -4.115209e-007, 6.915379e-007, 2.350906e-006,
  -4.955873e-007, -5.01921e-007, -7.191047e-007, -4.193435e-007, 
    1.231829e-007, -2.272373e-008, -9.39146e-007, -2.974011e-007, 
    8.725874e-007, 1.334027e-006, 5.912043e-007, 7.990748e-007, 
    2.540523e-006, 2.422929e-006, 1.166016e-006, 8.62653e-007, 2.441302e-007, 
    1.500795e-006, 3.016243e-006, 3.592298e-006, 3.569573e-006, 
    3.007675e-006, 2.948567e-006, 3.94322e-006, 4.88249e-006, 5.874659e-006, 
    6.100536e-006, 5.333373e-006, 2.86686e-006, 1.788139e-006, 4.425638e-007, 
    -8.600455e-007, -1.047303e-006, 9.55537e-007, 1.91306e-006, 
    1.433616e-006, 8.439019e-007, -1.086047e-006, -1.567229e-006, 
    1.18589e-007, 3.043066e-006, 4.891803e-006, 5.765756e-006, 5.124633e-006, 
    4.019961e-006, 3.298869e-006, 3.375485e-006, 5.296743e-006, 
    6.445869e-006, 5.346661e-006, 3.865857e-006, 3.394609e-006, 
    2.209593e-006, 2.156943e-006, 2.516184e-006, 3.904104e-006, 
    4.310408e-006, 4.949545e-006, 3.89268e-006, 3.719951e-006, 4.571677e-006, 
    3.580749e-006, 1.008684e-006, 4.77582e-007, 1.104673e-006, 3.024315e-006, 
    2.464031e-006, 4.51133e-007, -3.834566e-007, -1.175958e-007, 
    7.376093e-008, -1.095484e-006, -2.934659e-006, -2.903367e-006, 
    -5.681068e-007, 1.076981e-006, 2.524009e-006, 3.949181e-006, 
    5.18076e-006, 4.710505e-006, 3.283719e-006, 1.746043e-006, 1.052271e-006, 
    8.113675e-007, 3.725041e-006, 6.699438e-006, 6.299591e-006, 
    4.789357e-006, 3.658857e-006, 4.968791e-006, 6.707385e-006, 
    6.390364e-006, 2.702698e-006, -8.025509e-007, -9.48211e-007, 
    -6.534165e-007,
  -7.441886e-007, -1.66272e-007, -1.155709e-006, -1.300872e-006, 
    -7.835524e-007, 1.62423e-007, 2.090136e-006, 3.153707e-006, 
    2.763421e-006, 1.53929e-006, 9.67706e-007, 1.252815e-006, 1.040474e-006, 
    1.449138e-006, 2.105037e-006, 2.248462e-006, 2.352396e-006, 
    3.264099e-006, 3.908202e-006, 3.668914e-006, 2.727534e-006, 2.72033e-006, 
    3.105278e-006, 3.965695e-006, 3.559763e-006, 3.140172e-006, 
    2.803406e-006, 1.86637e-006, 1.794225e-006, 7.182352e-007, 
    -3.501737e-008, -6.08713e-007, -1.091262e-006, -9.557853e-007, 
    9.275936e-008, 6.699311e-007, -4.281601e-007, -1.12926e-006, 
    -7.269282e-007, -3.644582e-007, -4.457979e-008, -1.153594e-007, 
    5.494803e-007, 9.172909e-007, 5.725778e-007, 1.581386e-006, 
    2.799928e-006, 2.980356e-006, 2.897531e-006, 2.246474e-006, 
    1.610443e-006, 1.24139e-006, 6.920345e-007, 1.074373e-006, 2.008428e-006, 
    1.984835e-006, 1.973162e-006, 2.708286e-006, 2.821038e-006, 
    2.621363e-006, 1.938641e-006, 1.349425e-006, 1.419957e-006, 
    1.540408e-006, 1.190976e-006, 1.482169e-006, 1.774728e-006, 
    1.719594e-006, 6.740293e-007, -1.830358e-007, 5.027905e-007, 
    1.424674e-006, 2.223253e-006, 2.377853e-006, 1.486763e-006, 
    1.627704e-006, 2.728402e-006, 5.470962e-006, 6.316603e-006, 
    4.308422e-006, 2.562751e-006, 1.434485e-006, 1.198177e-006, 
    1.033644e-006, 8.732081e-007, 1.647944e-006, 2.082189e-006, 
    5.884713e-007, -6.154178e-007, -1.343712e-006, -1.122554e-006, 
    -7.150074e-007, -2.474826e-007, 3.866853e-007, -3.424784e-007, 
    -1.422564e-006,
  3.612286e-007, -1.99303e-007, -2.173056e-008, 1.768276e-007, 2.104789e-007, 
    2.565484e-007, 3.341584e-007, 1.412257e-006, 2.410387e-006, 
    2.216175e-006, 1.756101e-006, 1.432871e-006, 1.354888e-006, 
    1.027435e-006, 6.782511e-007, 5.587935e-007, 9.650985e-007, 
    1.543387e-006, 2.347679e-006, 2.945339e-006, 2.564987e-006, 
    2.076229e-006, 2.341717e-006, 2.175445e-006, 1.290192e-006, 
    5.720804e-007, 6.383907e-007, 8.330999e-007, 5.426509e-007, 
    -2.53196e-007, -2.545612e-007, 4.888825e-007, 8.36204e-007, 
    7.516392e-007, 6.083401e-007, 1.351907e-006, 1.900146e-006, 
    1.421323e-006, 1.247103e-006, 1.092007e-006, 7.707631e-007, 
    8.980433e-007, 1.074623e-006, 1.2363e-006, 1.549845e-006, 1.956274e-006, 
    2.593175e-006, 2.673516e-006, 2.530838e-006, 2.396107e-006, 
    2.520532e-006, 2.102181e-006, 1.592065e-006, 1.201654e-006, 
    9.169189e-007, 8.011857e-007, 1.072512e-006, 1.68408e-006, 1.81372e-006, 
    2.015009e-006, 2.039721e-006, 1.790002e-006, 1.614789e-006, 
    2.052263e-006, 2.792726e-006, 2.653152e-006, 1.936654e-006, 
    1.262998e-006, 1.09089e-006, 2.040342e-006, 2.738957e-006, 2.4649e-006, 
    2.130246e-006, 1.983593e-006, 1.644839e-006, 1.467268e-006, 
    1.827627e-006, 2.121926e-006, 1.667564e-006, 9.578962e-007, 
    7.531298e-007, 8.569409e-007, 1.0478e-006, 1.021971e-006, 7.094195e-007, 
    4.429371e-007, 5.046527e-007, 1.5758e-007, -6.557752e-007, 
    -1.090144e-006, -8.60914e-007, -3.97612e-007, 7.624385e-008, 
    2.947945e-007, 6.880618e-007, 9.925416e-007,
  8.200604e-007, 1.123175e-006, 1.703079e-006, 2.145767e-006, 2.242749e-006, 
    2.302726e-006, 2.393499e-006, 2.399335e-006, 2.246598e-006, 
    2.016872e-006, 1.908342e-006, 1.599144e-006, 1.098836e-006, 
    6.965056e-007, 6.181499e-007, 4.171079e-007, 4.008416e-007, 
    5.786615e-007, 8.641427e-007, 1.319747e-006, 1.756101e-006, 
    1.805524e-006, 1.362711e-006, 7.209683e-007, 3.752612e-007, 
    1.242997e-007, -1.822909e-007, -1.043081e-007, 3.560135e-007, 
    9.239961e-007, 1.226987e-006, 1.262749e-006, 1.095359e-006, 9.20023e-007, 
    9.735422e-007, 1.020109e-006, 1.340981e-006, 1.760945e-006, 
    2.061575e-006, 2.223502e-006, 2.142663e-006, 1.961987e-006, 
    1.874194e-006, 1.944104e-006, 2.124906e-006, 1.999363e-006, 1.66744e-006, 
    1.607586e-006, 2.088645e-006, 2.645204e-006, 3.112232e-006, 3.60844e-006, 
    3.933534e-006, 4.036972e-006, 4.097944e-006, 3.975754e-006, 
    3.512328e-006, 2.987186e-006, 2.511715e-006, 2.18985e-006, 2.062817e-006, 
    1.850475e-006, 1.636397e-006, 1.723196e-006, 2.062693e-006, 2.29838e-006, 
    2.454842e-006, 2.303472e-006, 1.821791e-006, 1.356875e-006, 
    1.120568e-006, 9.072319e-007, 8.321058e-007, 1.008809e-006, 
    1.307577e-006, 1.702954e-006, 1.937399e-006, 2.218037e-006, 
    2.586221e-006, 2.70692e-006, 2.316262e-006, 1.790002e-006, 1.366809e-006, 
    9.377795e-007, 1.145651e-006, 1.698608e-006, 1.986946e-006, 
    1.606469e-006, 1.074126e-006, 6.857017e-007, 2.630054e-007, 
    7.525068e-008, 4.839158e-007, 9.472169e-007, 9.798759e-007, 8.62281e-007,
  7.381041e-007, 1.094366e-006, 1.445661e-006, 1.614044e-006, 1.542643e-006, 
    1.274546e-006, 9.249893e-007, 5.139659e-007, 9.648511e-008, 
    -9.362884e-008, 2.70702e-008, 2.60522e-007, 4.475314e-007, 4.973263e-007, 
    4.102785e-007, 3.212444e-007, 2.889587e-007, 3.300606e-007, 
    3.546479e-007, 2.653651e-007, 9.822361e-008, -1.291392e-008, 
    -5.091351e-009, 1.285225e-007, 2.723182e-007, 2.7741e-007, 1.38084e-007, 
    -1.153603e-007, -3.968671e-007, -5.171942e-007, -3.13793e-007, 
    1.830358e-007, 8.779271e-007, 1.560524e-006, 1.977383e-006, 
    2.070268e-006, 1.942119e-006, 1.706555e-006, 1.521905e-006, 
    1.494462e-006, 1.639376e-006, 1.837438e-006, 1.84315e-006, 1.619012e-006, 
    1.338869e-006, 1.176695e-006, 1.121312e-006, 1.116966e-006, 
    1.165022e-006, 1.364326e-006, 1.776219e-006, 2.311419e-006, 
    2.803529e-006, 3.049523e-006, 3.019471e-006, 2.914543e-006, 
    2.852827e-006, 2.744049e-006, 2.513454e-006, 2.26299e-006, 2.064804e-006, 
    2.031526e-006, 2.191092e-006, 2.41672e-006, 2.622604e-006, 2.818802e-006, 
    2.926961e-006, 2.924973e-006, 2.847488e-006, 2.776831e-006, 
    2.675007e-006, 2.509231e-006, 2.251938e-006, 1.862273e-006, 
    1.422688e-006, 9.560335e-007, 5.299844e-007, 1.703697e-007, 
    -8.580582e-008, -2.885854e-007, -4.426888e-007, -5.016723e-007, 
    -4.315129e-007, -2.303468e-007, 7.152585e-008, 4.857775e-007, 
    8.949387e-007, 1.21519e-006, 1.473849e-006, 1.581013e-006, 1.531218e-006, 
    1.362463e-006, 1.037245e-006, 6.674481e-007, 4.785761e-007, 5.318479e-007,
  3.991036e-007, 3.814703e-007, 3.896648e-007, 4.294025e-007, 4.832946e-007, 
    5.2837e-007, 5.396705e-007, 5.128486e-007, 4.513813e-007, 3.675623e-007, 
    2.761681e-007, 1.90611e-007, 1.352282e-007, 1.308827e-007, 1.708668e-007, 
    2.415227e-007, 3.226096e-007, 3.840773e-007, 4.091612e-007, 
    3.932664e-007, 3.42478e-007, 2.59156e-007, 1.549724e-007, 3.501737e-008, 
    -8.667575e-008, -2.156949e-007, -3.417335e-007, -4.480289e-007, 
    -5.155807e-007, -5.256379e-007, -4.717458e-007, -3.606083e-007, 
    -2.119687e-007, -5.538277e-008, 8.692314e-008, 2.017869e-007, 
    2.858542e-007, 3.387531e-007, 3.628429e-007, 3.576283e-007, 
    3.234795e-007, 2.644956e-007, 1.916042e-007, 1.221897e-007, 
    6.941445e-008, 3.563855e-008, 2.35932e-008, 2.930574e-008, 4.346157e-008, 
    6.134314e-008, 7.587187e-008, 8.977986e-008, 1.009553e-007, 9.48703e-008, 
    5.43896e-008, -2.173056e-008, -1.260387e-007, -2.356865e-007, 
    -3.265841e-007, -3.905343e-007, -4.351141e-007, -4.610665e-007, 
    -4.559761e-007, -4.123895e-007, -3.293162e-007, -2.169363e-007, 
    -8.84138e-008, 4.221965e-008, 1.646576e-007, 2.55307e-007, 2.895795e-007, 
    2.6611e-007, 1.971921e-007, 9.760333e-008, -3.079549e-008, -1.81918e-007, 
    -3.46452e-007, -5.055226e-007, -6.239861e-007, -6.884338e-007, 
    -6.947666e-007, -6.474552e-007, -5.658721e-007, -4.600729e-007, 
    -3.403675e-007, -2.168117e-007, -8.940697e-008, 2.210345e-008, 
    1.112621e-007, 1.829112e-007, 2.476072e-007, 3.054738e-007, 
    3.530331e-007, 3.936393e-007, 4.198409e-007, 4.209578e-007,
  -1.122555e-007, -1.324961e-007, -1.46528e-007, -1.524886e-007, 
    -1.522402e-007, -1.423061e-007, -1.216927e-007, -9.07728e-008, 
    -5.30232e-008, -1.266608e-008, 3.402431e-008, 8.083884e-008, 
    1.290192e-007, 1.739712e-007, 2.194197e-007, 2.620121e-007, 3.0001e-007, 
    3.33786e-007, 3.624707e-007, 3.865609e-007, 4.04194e-007, 4.145006e-007, 
    4.200887e-007, 4.209578e-007, 4.162391e-007, 4.046907e-007, 
    3.914038e-007, 3.786137e-007, 3.669411e-007, 3.534058e-007, 
    3.417333e-007, 3.301849e-007, 3.186366e-007, 3.106892e-007, 
    3.019968e-007, 2.883374e-007, 2.72567e-007, 2.519538e-007, 2.298505e-007, 
    2.0427e-007, 1.817941e-007, 1.616776e-007, 1.425545e-007, 1.236796e-007, 
    1.076609e-007, 9.561586e-008, 9.474661e-008, 1.024456e-007, 
    1.134972e-007, 1.312544e-007, 1.593182e-007, 1.925976e-007, 
    2.287329e-007, 2.715735e-007, 3.201267e-007, 3.7166e-007, 4.255523e-007, 
    4.770857e-007, 5.289912e-007, 5.844979e-007, 6.371488e-007, 
    6.868195e-007, 7.345031e-007, 7.748604e-007, 8.096297e-007, 
    8.385628e-007, 8.509805e-007, 8.553268e-007, 8.504837e-007, 
    8.374452e-007, 8.229167e-007, 8.086363e-007, 7.993233e-007, 
    7.919966e-007, 7.830561e-007, 7.746119e-007, 7.645538e-007, 
    7.520118e-007, 7.349997e-007, 7.141382e-007, 6.886821e-007, 
    6.541609e-007, 6.080916e-007, 5.512188e-007, 4.892549e-007, 
    4.218271e-007, 3.529092e-007, 2.84364e-007, 2.1557e-007, 1.50626e-007, 
    9.35047e-008, 4.656613e-008, 4.718686e-009, -3.265836e-008, 
    -6.270898e-008, -8.90343e-008,
  -9.9217e-008, -8.046629e-008, -4.02332e-008, 1.154831e-008, 4.333754e-008, 
    4.358594e-008, 2.967806e-008, 2.22276e-008, 2.02408e-008, 2.297259e-008, 
    4.197153e-008, 7.276731e-008, 9.983779e-008, 1.292676e-007, 
    1.595666e-007, 1.80304e-007, 2.01414e-007, 2.266219e-007, 2.613912e-007, 
    2.918144e-007, 3.134211e-007, 3.094474e-007, 2.974023e-007, 
    3.099442e-007, 3.525366e-007, 3.983577e-007, 4.250556e-007, 
    4.275392e-007, 4.102786e-007, 3.706664e-007, 3.178914e-007, 
    2.599011e-007, 2.212822e-007, 2.118448e-007, 2.170602e-007, 
    2.252559e-007, 2.369285e-007, 2.584109e-007, 2.843639e-007, 
    3.011276e-007, 3.063431e-007, 3.123035e-007, 3.517915e-007, 
    4.054358e-007, 4.008411e-007, 3.381322e-007, 2.775342e-007, 
    2.613913e-007, 2.709528e-007, 2.80266e-007, 2.786519e-007, 3.452101e-007, 
    5.075087e-007, 7.116548e-007, 8.907168e-007, 9.87947e-007, 9.807447e-007, 
    9.361654e-007, 9.114544e-007, 8.712213e-007, 7.624426e-007, 
    5.599111e-007, 3.53406e-007, 2.006689e-007, 1.251697e-007, 1.424303e-007, 
    1.888723e-007, 2.277395e-007, 2.313404e-007, 2.279878e-007, 2.83743e-007, 
    4.017106e-007, 5.314748e-007, 6.242344e-007, 6.763887e-007, 
    6.798655e-007, 6.599976e-007, 6.334235e-007, 5.397947e-007, 
    4.167359e-007, 3.231066e-007, 2.489737e-007, 1.322478e-007, 
    -6.072241e-008, -2.702077e-007, -4.690141e-007, -6.434821e-007, 
    -7.127724e-007, -6.854534e-007, -5.698453e-007, -4.044425e-007, 
    -2.50091e-007, -1.486392e-007, -9.921678e-008, -9.064888e-008, 
    -9.896848e-008,
  -1.945841e-007, -6.792447e-008, 2.396609e-008, 3.837044e-008, 
    3.414846e-008, 8.717177e-008, 1.451621e-007, 1.73226e-007, 1.800557e-007, 
    1.636644e-007, 1.73971e-007, 1.902382e-007, 2.138317e-007, 2.63378e-007, 
    3.498047e-007, 3.986061e-007, 3.955017e-007, 3.552685e-007, 
    3.006309e-007, 2.447516e-007, 1.862645e-007, 1.35973e-007, 1.213203e-007, 
    1.423061e-007, 1.990547e-007, 2.782792e-007, 3.37263e-007, 3.476937e-007, 
    3.180157e-007, 2.590318e-007, 2.381702e-007, 2.375493e-007, 
    2.499669e-007, 2.707044e-007, 2.935529e-007, 3.186365e-007, 
    3.535301e-007, 4.169842e-007, 4.649162e-007, 4.827977e-007, 
    5.030385e-007, 5.345792e-007, 5.736947e-007, 6.797413e-007, 7.915e-007, 
    8.853774e-007, 9.493281e-007, 1.024703e-006, 1.065557e-006, 
    9.339306e-007, 7.893891e-007, 8.148454e-007, 1.121933e-006, 
    1.492848e-006, 1.809374e-006, 2.006193e-006, 1.991665e-006, 
    1.819308e-006, 1.594548e-006, 1.390278e-006, 1.00856e-006, 6.66827e-007, 
    4.609424e-007, 4.089129e-007, 4.332514e-007, 6.38142e-007, 1.086667e-006, 
    1.575798e-006, 1.892075e-006, 1.883258e-006, 1.633167e-006, 
    1.375129e-006, 1.23841e-006, 1.207864e-006, 1.13137e-006, 1.017253e-006, 
    1.044696e-006, 1.120816e-006, 1.115104e-006, 9.227542e-007, 
    5.335855e-007, 2.266215e-007, 1.10269e-007, -1.287708e-007, 
    -4.940975e-007, -8.698553e-007, -1.164402e-006, -1.259893e-006, 
    -1.314283e-006, -1.161546e-006, -8.594243e-007, -6.544092e-007, 
    -6.097061e-007, -5.571792e-007, -4.321337e-007, -3.123034e-007,
  1.511227e-007, 1.286467e-007, 9.35047e-008, 1.31627e-007, 1.591941e-007, 
    1.347313e-007, 1.559655e-007, 2.279878e-007, 2.546857e-007, 
    3.111859e-007, 3.97116e-007, 4.177292e-007, 3.807247e-007, 4.081676e-007, 
    5.748122e-007, 6.016344e-007, 4.568448e-007, 3.427267e-007, 
    3.259629e-007, 3.28074e-007, 2.296021e-007, 1.459073e-007, 2.063811e-007, 
    2.594044e-007, 2.399088e-007, 2.476077e-007, 2.795209e-007, 
    3.467003e-007, 4.066775e-007, 2.966573e-007, 1.68259e-007, 1.127521e-007, 
    1.130005e-007, 1.158566e-007, 1.526128e-007, 2.207855e-007, 
    2.725671e-007, 3.188849e-007, 3.855675e-007, 2.951671e-007, 
    1.107653e-007, -7.388496e-008, -1.439205e-007, 1.082819e-007, 
    6.010134e-007, 1.12628e-006, 1.337876e-006, 1.471862e-006, 1.358241e-006, 
    1.188368e-006, 1.213327e-006, 1.102065e-006, 7.957219e-007, 
    1.003717e-006, 1.569093e-006, 1.820549e-006, 1.89878e-006, 1.936033e-006, 
    1.85892e-006, 1.806146e-006, 1.729776e-006, 1.493469e-006, 9.833529e-007, 
    1.477702e-007, -4.199646e-007, -4.477797e-007, -1.395747e-007, 
    5.469965e-007, 1.374508e-006, 1.662102e-006, 1.683955e-006, 
    1.822536e-006, 1.92585e-006, 1.89518e-006, 2.304712e-006, 3.045549e-006, 
    3.454586e-006, 3.309176e-006, 2.979114e-006, 2.673764e-006, 
    2.430006e-006, 2.056857e-006, 1.583372e-006, 1.378854e-006, 
    1.242633e-006, 1.00558e-006, 6.545333e-007, 3.912792e-007, 7.448762e-010, 
    -5.832562e-007, -5.928177e-007, -9.36293e-008, 3.254663e-007, 
    5.425263e-007, 4.255523e-007, 2.325824e-007,
  -3.539026e-008, -1.055514e-008, 1.117587e-008, -6.134314e-008, 
    -9.437395e-008, -9.524319e-008, 6.146729e-008, 4.675239e-007, 
    8.848806e-007, 1.028553e-006, 1.100078e-006, 1.004214e-006, 8.36576e-007, 
    6.057323e-007, 5.993993e-007, 5.905827e-007, 5.255143e-007, 4.69635e-007, 
    4.156182e-007, 3.352762e-007, 3.29564e-007, 3.219893e-007, 4.819283e-007, 
    8.031725e-007, 8.277595e-007, 6.268422e-007, 5.31599e-007, 4.974504e-007, 
    4.924834e-007, 5.806485e-007, 5.564343e-007, 7.482865e-007, 
    9.095916e-007, 8.599211e-007, 8.061529e-007, 7.465483e-007, 
    5.374354e-007, 4.450478e-007, 5.451338e-007, 3.227342e-007, 
    -1.045564e-007, -2.447514e-007, -5.873517e-008, 4.454205e-007, 
    1.095608e-006, 1.155709e-006, 5.021693e-007, 3.003825e-007, 
    1.492227e-006, 2.328431e-006, 2.69711e-006, 2.776334e-006, 3.290176e-006, 
    4.097943e-006, 3.820285e-006, 2.863135e-006, 2.277145e-006, 
    2.943848e-006, 3.781046e-006, 4.287808e-006, 4.538646e-006, 3.6786e-006, 
    2.555922e-006, 2.034258e-006, 2.445156e-006, 2.072131e-006, 
    1.228849e-006, 4.195917e-007, 7.723775e-007, 1.892447e-006, 
    2.326691e-006, 2.542635e-006, 2.150362e-006, 1.591445e-006, 
    2.287328e-006, 2.642721e-006, 2.075981e-006, 1.688053e-006, 1.88686e-006, 
    2.030903e-006, 1.540408e-006, 1.222268e-006, 1.371279e-006, 
    1.224503e-006, 1.003593e-006, 1.049787e-006, 1.17893e-006, 1.150866e-006, 
    5.185602e-007, -5.662423e-008, -8.294955e-008, 1.502531e-007, 
    5.086258e-007, 3.204987e-007, 7.202289e-008, -1.887474e-008,
  1.087412e-006, 1.903002e-006, 2.242376e-006, 2.032394e-006, 1.571203e-006, 
    8.642673e-007, 6.347891e-007, 8.816523e-007, 1.508618e-006, 
    2.172341e-006, 2.26361e-006, 2.845253e-006, 3.448502e-006, 3.538281e-006, 
    3.236532e-006, 2.771616e-006, 2.423425e-006, 2.171844e-006, 
    2.279629e-006, 2.188732e-006, 2.226233e-006, 2.362579e-006, 
    2.446522e-006, 2.423922e-006, 1.628076e-006, 1.098836e-006, 
    1.828869e-006, 2.215181e-006, 2.187615e-006, 2.245481e-006, 
    1.733129e-006, 1.493966e-006, 1.567354e-006, 1.789754e-006, 
    2.203013e-006, 3.37561e-006, 3.596769e-006, 2.58585e-006, 1.488874e-006, 
    1.661479e-006, 2.86003e-006, 3.168236e-006, 2.683822e-006, 1.650676e-006, 
    1.173217e-006, 2.342958e-006, 2.694504e-006, 3.980473e-006, 5.72813e-006, 
    7.023042e-006, 6.312008e-006, 5.172193e-006, 4.535788e-006, 
    4.823009e-006, 4.822388e-006, 4.846974e-006, 4.166862e-006, 
    4.371008e-006, 5.238378e-006, 5.107746e-006, 3.887589e-006, 
    2.906595e-006, 2.68221e-006, 2.066915e-006, 1.985332e-006, 1.727665e-006, 
    1.397108e-006, 1.474594e-006, 1.555929e-006, 2.25318e-006, 2.549837e-006, 
    2.539903e-006, 2.430504e-006, 2.412125e-006, 2.571194e-006, 
    2.194072e-006, 2.430132e-006, 2.213194e-006, 1.504397e-006, 
    5.492329e-007, -3.830846e-007, -4.258e-007, -1.676381e-008, 
    1.239277e-007, 3.27329e-007, 8.674961e-007, 2.040962e-006, 3.386413e-006, 
    3.408144e-006, 2.389774e-006, 2.242004e-006, 3.390636e-006, 
    3.837298e-006, 3.071254e-006, 1.798446e-006, 8.900961e-007,
  2.99886e-006, 3.955636e-006, 3.743793e-006, 3.691392e-006, 2.54127e-006, 
    1.2779e-006, 2.01476e-006, 3.272668e-006, 4.098936e-006, 4.214546e-006, 
    4.349153e-006, 5.497162e-006, 6.049375e-006, 6.289283e-006, 
    6.439537e-006, 5.758057e-006, 6.438047e-006, 8.550287e-006, 
    9.773672e-006, 9.136896e-006, 7.456664e-006, 6.045152e-006, 
    5.049879e-006, 4.352381e-006, 3.597389e-006, 3.710513e-006, 
    3.792966e-006, 2.817065e-006, 3.265838e-006, 4.686042e-006, 
    5.099302e-006, 5.499523e-006, 6.193794e-006, 5.706277e-006, 
    5.655238e-006, 5.934016e-006, 5.942209e-006, 7.852292e-006, 
    8.025145e-006, 6.872664e-006, 6.48933e-006, 7.167831e-006, 6.512306e-006, 
    8.17987e-006, 1.005059e-005, 9.762496e-006, 9.190911e-006, 9.40847e-006, 
    9.396299e-006, 8.979689e-006, 6.184602e-006, 3.584475e-006, 
    3.233179e-006, 3.947318e-006, 4.48587e-006, 4.717707e-006, 4.94284e-006, 
    4.79867e-006, 4.642705e-006, 4.086767e-006, 3.758198e-006, 4.486491e-006, 
    2.879897e-006, 2.77584e-006, 3.034249e-006, 3.568208e-006, 4.201506e-006, 
    4.128616e-006, 4.902235e-006, 5.38888e-006, 3.993138e-006, 4.063175e-006, 
    4.8168e-006, 3.850957e-006, 2.693385e-006, 2.029539e-006, 1.838307e-006, 
    2.80651e-006, 3.918136e-006, 3.459305e-006, 3.842761e-006, 4.118682e-006, 
    2.884493e-006, 2.041956e-006, 2.255787e-006, 2.876917e-006, 
    3.612415e-006, 3.258016e-006, 2.440437e-006, 1.593058e-006, 
    2.408897e-006, 3.736093e-006, 3.25938e-006, 1.798943e-006, 8.856259e-007, 
    1.921132e-006,
  3.096461e-006, 1.596411e-006, 9.501973e-007, 1.076235e-006, 1.124416e-006, 
    2.182274e-006, 3.090501e-006, 3.216415e-006, 4.061063e-006, 
    4.865105e-006, 4.875536e-006, 4.567331e-006, 5.830327e-006, 
    7.572398e-006, 7.975723e-006, 8.238852e-006, 7.915372e-006, 
    7.505094e-006, 6.644426e-006, 5.08676e-006, 4.370015e-006, 5.356222e-006, 
    7.666897e-006, 7.812307e-006, 8.150189e-006, 8.388733e-006, 
    9.246667e-006, 9.045751e-006, 8.044764e-006, 7.464363e-006, 
    7.484728e-006, 7.732709e-006, 7.785111e-006, 9.277464e-006, 
    8.932999e-006, 7.828947e-006, 8.395191e-006, 9.302421e-006, 
    9.068102e-006, 8.073697e-006, 9.467329e-006, 1.025498e-005, 
    8.443121e-006, 9.696558e-006, 1.177576e-005, 1.22259e-005, 8.951003e-006, 
    7.29772e-006, 5.649277e-006, 3.66196e-006, 4.738073e-006, 5.364169e-006, 
    5.513057e-006, 4.173442e-006, 3.397216e-006, 2.89691e-006, 2.958377e-006, 
    4.010275e-006, 4.353125e-006, 4.65326e-006, 5.179892e-006, 5.958105e-006, 
    5.392232e-006, 4.828971e-006, 4.185364e-006, 4.380694e-006, 
    5.470714e-006, 5.780656e-006, 6.535152e-006, 5.072976e-006, 
    3.226474e-006, 4.769861e-006, 5.773081e-006, 5.501881e-006, 
    5.539878e-006, 5.257129e-006, 6.044904e-006, 6.497776e-006, 
    4.625694e-006, 4.238511e-006, 4.389138e-006, 3.75261e-006, 4.120295e-006, 
    2.360221e-006, 2.557039e-006, 3.847232e-006, 4.285946e-006, 
    5.094085e-006, 5.201003e-006, 5.086138e-006, 5.147358e-006, 
    5.713106e-006, 5.048141e-006, 3.140916e-006, 2.754106e-006, 3.263354e-006,
  2.713128e-006, 3.618003e-006, 4.848092e-006, 4.293894e-006, 3.8332e-006, 
    5.293141e-006, 6.454562e-006, 6.475797e-006, 6.418924e-006, 
    7.268412e-006, 7.876008e-006, 7.005285e-006, 7.297844e-006, 
    6.957849e-006, 7.169694e-006, 7.722403e-006, 7.968398e-006, 
    7.505218e-006, 7.354467e-006, 7.686143e-006, 8.794541e-006, 
    1.135481e-005, 1.244483e-005, 1.165581e-005, 1.065346e-005, 
    1.072263e-005, 9.812788e-006, 9.515259e-006, 9.65347e-006, 8.509433e-006, 
    5.604699e-006, 4.310163e-006, 5.872673e-006, 8.157887e-006, 
    7.798646e-006, 8.434554e-006, 9.628635e-006, 9.44448e-006, 7.53763e-006, 
    8.980183e-006, 1.081477e-005, 9.541709e-006, 8.63634e-006, 8.420895e-006, 
    7.019315e-006, 5.842743e-006, 7.026891e-006, 6.402033e-006, 4.21293e-006, 
    2.768138e-006, 2.403309e-006, 3.641595e-006, 3.534431e-006, 
    4.738942e-006, 3.439685e-006, 7.99695e-007, 2.114475e-006, 2.75088e-006, 
    2.941117e-006, 3.171959e-006, 3.3658e-006, 2.337869e-006, 1.445909e-006, 
    1.872952e-006, 3.178789e-006, 4.480284e-006, 3.344192e-006, 
    5.160764e-007, 1.484777e-006, 3.439683e-006, 5.096073e-006, 
    4.591047e-006, 4.052494e-006, 4.58248e-006, 4.876158e-006, 3.482402e-006, 
    4.179899e-006, 5.19678e-006, 4.30147e-006, 4.986301e-006, 4.500027e-006, 
    3.499164e-006, 3.082554e-006, 3.17643e-006, 3.563488e-006, 3.470481e-006, 
    3.08392e-006, 1.579152e-006, 2.072627e-006, 2.927705e-006, 2.835815e-006, 
    3.477186e-006, 3.537662e-006, 4.14153e-006, 3.650412e-006, 3.335748e-006,
  4.284953e-006, 5.679578e-006, 6.204597e-006, 5.159527e-006, 5.77333e-006, 
    7.672235e-006, 7.682667e-006, 6.356833e-006, 5.748871e-006, 
    6.797536e-006, 6.812686e-006, 7.314857e-006, 7.997203e-006, 9.48136e-006, 
    1.020406e-005, 1.004698e-005, 1.028789e-005, 1.068674e-005, 
    1.101283e-005, 1.073666e-005, 9.939446e-006, 8.749465e-006, 
    8.947649e-006, 8.396431e-006, 6.762024e-006, 6.488339e-006, 7.66317e-006, 
    8.744868e-006, 8.055071e-006, 6.615617e-006, 6.095692e-006, 
    6.488586e-006, 6.76289e-006, 6.659207e-006, 6.68069e-006, 6.763388e-006, 
    6.691738e-006, 4.450605e-006, 4.099062e-006, 4.734844e-006, 
    7.113566e-006, 5.82449e-006, 4.970902e-006, 7.569293e-006, 5.291276e-006, 
    3.406778e-006, 4.323449e-006, 6.00169e-006, 3.323828e-006, 2.329798e-006, 
    2.401943e-006, 3.231316e-006, 8.25401e-007, -1.022965e-006, 
    -2.006442e-006, -2.337993e-006, -1.493841e-006, -9.453543e-007, 
    -1.584242e-006, -9.196501e-007, -2.48474e-009, -2.471097e-008, 
    -3.352761e-008, -3.974492e-009, -6.283317e-007, -8.239113e-007, 
    5.915772e-007, 1.267592e-006, 2.643714e-006, 3.294646e-006, 
    3.996365e-006, 5.155802e-006, 5.690503e-006, 4.464884e-006, 
    3.215297e-006, 3.021087e-006, 4.624573e-006, 4.383301e-006, 
    3.233801e-006, 1.660734e-006, 1.268834e-006, 1.755854e-006, 
    1.825641e-006, 2.320236e-006, 1.841909e-006, 2.763421e-006, 
    4.144013e-006, 4.635129e-006, 4.612159e-006, 4.559755e-006, 4.82723e-006, 
    5.504489e-006, 7.513414e-006, 6.46909e-006, 5.788977e-006, 4.3042e-006,
  4.083786e-006, 3.548339e-006, 4.025675e-006, 5.429982e-006, 5.7254e-006, 
    4.909685e-006, 4.721433e-006, 4.767131e-006, 6.172806e-006, 
    5.133825e-006, 5.157417e-006, 7.476036e-006, 8.287279e-006, 
    7.008635e-006, 6.416314e-006, 7.958337e-006, 9.645519e-006, 
    9.836131e-006, 9.20122e-006, 7.904942e-006, 6.453072e-006, 6.657468e-006, 
    8.60095e-006, 7.835402e-006, 5.650025e-006, 5.427872e-006, 4.517162e-006, 
    5.403283e-006, 6.436432e-006, 6.15741e-006, 6.348018e-006, 7.721039e-006, 
    4.644691e-006, 1.729903e-006, 2.231573e-006, 1.729899e-006, 
    7.039562e-007, 3.228706e-008, -6.013834e-007, -3.784917e-007, 
    1.945344e-006, 1.539789e-006, -3.198784e-007, -5.985203e-008, 
    2.451241e-006, 1.652166e-006, 9.338073e-007, 2.067165e-006, 
    1.031533e-006, 6.527953e-007, -2.978617e-006, -3.424038e-006, 
    -2.303721e-006, -2.753859e-006, -3.222502e-006, -1.34272e-006, 
    -1.301989e-006, -1.374259e-006, -2.854938e-006, -4.398335e-007, 
    -1.759206e-006, -3.568332e-006, -2.347926e-006, -1.314529e-006, 
    -2.509356e-006, -2.609193e-006, -1.195822e-007, 1.13137e-006, 
    8.348361e-007, 6.526716e-007, 9.730466e-007, 2.103921e-006, 
    4.654139e-007, -1.553199e-006, -1.687433e-006, 1.118704e-006, 
    3.897399e-006, 2.178178e-006, -5.262591e-007, -1.178061e-006, 
    -1.496822e-006, -2.392382e-006, -2.346933e-006, -1.614168e-006, 
    7.399667e-007, 4.786998e-007, 1.601751e-006, 4.8322e-006, 4.680083e-006, 
    4.752601e-006, 5.227203e-006, 6.729859e-006, 7.245937e-006, 
    6.901226e-006, 5.617863e-006, 5.226582e-006,
  3.804515e-006, 4.99512e-006, 5.203608e-006, 5.287427e-006, 2.662215e-006, 
    1.938886e-006, 2.821285e-006, 4.948302e-006, 5.524855e-006, 
    6.245325e-006, 6.253396e-006, 6.238497e-006, 7.350867e-006, 
    7.494909e-006, 6.099544e-006, 5.60383e-006, 6.653991e-006, 5.620594e-006, 
    5.951028e-006, 5.90707e-006, 6.226946e-006, 7.185216e-006, 6.810202e-006, 
    4.662572e-006, 4.400685e-006, 4.662696e-006, 2.902372e-006, 
    2.513327e-006, 4.824375e-006, 4.31612e-006, 1.40518e-006, -1.139939e-006, 
    -2.978122e-006, -4.075839e-006, -4.709142e-006, -5.362432e-006, 
    -6.230795e-006, -5.499769e-006, -5.062051e-006, -6.596245e-006, 
    -6.96443e-006, -1.286095e-006, -1.007102e-007, -7.96219e-007, 
    -7.947529e-008, -2.604353e-006, -2.148003e-006, 1.046683e-006, 
    7.189919e-008, -1.390776e-006, 9.859596e-007, -1.20091e-006, 
    -5.46885e-006, -2.64508e-006, -1.195818e-006, 2.142539e-006, 
    3.380082e-007, -3.977384e-007, -4.482021e-006, -2.126893e-006, 
    -3.043562e-006, -4.771477e-006, -2.159801e-006, -1.841534e-006, 
    -2.291177e-006, 9.884388e-008, -3.710375e-007, -8.742027e-007, 
    -1.678616e-006, -3.701822e-006, -1.379474e-006, -3.677604e-006, 
    -5.394719e-006, -2.704561e-006, -7.475392e-007, 8.553288e-007, 
    -1.045068e-006, -5.152571e-006, -2.383316e-006, -1.49409e-006, 
    -2.604351e-006, -2.594043e-006, -1.331173e-007, 5.41906e-007, 
    -8.774314e-007, 9.48583e-007, 2.972658e-006, 6.021557e-006, 
    7.535768e-006, 1.020245e-005, 1.255026e-005, 9.366373e-006, 
    7.400664e-006, 6.224342e-006, 4.29327e-006, 3.045177e-006,
  2.22884e-006, 1.654527e-006, 1.771623e-006, -2.085912e-006, -8.131065e-007, 
    2.012652e-006, 3.385543e-006, 6.578739e-006, 6.920845e-006, 
    7.097298e-006, 6.547323e-006, 4.025052e-006, 2.239769e-006, 
    -1.366439e-006, 2.880879e-007, 2.413988e-006, 3.012021e-006, 
    1.829616e-006, 1.745047e-006, 2.694254e-006, 3.227964e-006, 
    2.584235e-006, -8.419156e-007, -7.071867e-007, -1.868233e-006, 
    -4.155314e-006, -6.264945e-006, -6.829698e-006, -7.633618e-006, 
    -7.698562e-006, -7.914256e-006, -8.144356e-006, -8.736177e-006, 
    -8.825089e-006, -8.941939e-006, -8.126844e-006, -7.034467e-006, 
    -8.184586e-006, -8.193278e-006, -5.937865e-006, -4.369393e-006, 
    -1.638631e-006, -2.473589e-007, 4.351132e-007, -9.528048e-007, 
    -1.372398e-006, -1.770881e-006, -1.519049e-006, -1.632174e-006, 
    -1.819681e-006, 7.064373e-007, -2.475703e-006, -2.075856e-006, 
    3.208715e-007, 1.463421e-006, -2.163142e-007, -1.346569e-006, 
    -5.041064e-006, -6.197517e-006, -1.756722e-006, -2.310924e-006, 
    -3.270059e-006, -1.023211e-006, -3.419318e-006, -4.731241e-006, 
    -3.851332e-006, -3.152836e-006, -3.052133e-006, -9.206451e-007, 
    3.202509e-006, 7.40074e-008, -1.097345e-006, 2.315763e-006, 
    1.169989e-006, -1.552577e-006, -5.428246e-006, -9.053078e-006, 
    -5.787238e-006, -1.752998e-006, -5.469965e-007, -8.787956e-007, 
    -6.581104e-009, -1.934046e-006, -2.222385e-006, -1.626708e-006, 
    4.000834e-006, 8.355826e-006, 1.199854e-005, 1.257782e-005, 
    1.228005e-005, 8.54929e-006, 3.443904e-006, 1.509485e-006, 2.261258e-007, 
    1.595654e-007, 1.102559e-006,
  -5.472699e-006, -5.783513e-006, -4.44899e-006, -3.295267e-006, 
    -1.729777e-006, -1.816699e-006, 1.159187e-006, 3.804887e-006, 
    6.048134e-006, 3.038967e-006, -2.738958e-006, -4.746518e-006, 
    -5.457303e-006, -8.179486e-007, 5.99648e-007, -1.546618e-006, 
    -4.198773e-006, -6.473314e-006, -7.044398e-006, -6.79617e-006, 
    -8.051096e-006, -8.189803e-006, -8.488943e-006, -9.219597e-006, 
    -8.846571e-006, -9.040907e-006, -8.929024e-006, -8.853649e-006, 
    -8.599336e-006, -7.255252e-006, -6.220242e-006, -6.877508e-006, 
    -9.675574e-006, -9.838986e-006, -9.578343e-006, -7.729232e-006, 
    -5.156422e-006, -4.720563e-006, -5.090236e-006, -1.540035e-006, 
    1.114855e-006, 2.702698e-006, 3.727153e-006, 2.847859e-006, 
    1.322976e-006, 1.974331e-008, -1.663961e-006, 2.481102e-009, 
    2.786765e-006, -1.442681e-006, -4.443402e-006, -2.672277e-006, 
    -2.313904e-006, -2.060457e-006, -1.216682e-006, -4.502137e-006, 
    -7.669874e-006, -6.987775e-006, -4.92893e-006, -9.017676e-007, 
    -3.686298e-006, -6.682672e-006, -5.198643e-006, -8.828938e-007, 
    2.120436e-006, 5.199254e-007, 1.672903e-006, 6.068869e-006, 
    4.908445e-006, 3.392499e-006, 2.148747e-006, 8.787974e-007, 
    2.980232e-007, -2.762899e-007, -1.279263e-006, -4.17543e-006, 
    -5.491449e-006, -4.794199e-006, 5.309776e-007, -3.890455e-007, 
    -7.746121e-007, -1.570706e-006, -2.660479e-006, -1.021352e-006, 
    5.445007e-006, 8.053954e-006, 9.608888e-006, 1.088381e-005, 
    4.719572e-006, 1.683085e-006, -8.451425e-007, -2.834324e-006, 
    -1.230837e-006, -9.608739e-007, -1.12268e-006, -3.931051e-006,
  -6.404396e-006, -5.881737e-006, -5.081793e-006, -4.504869e-006, 
    -2.91864e-006, -2.209345e-006, -9.433679e-007, -1.759206e-006, 
    -2.96856e-006, -5.238751e-006, -1.06146e-005, -9.162726e-006, 
    -6.789962e-006, -5.033116e-006, -5.220993e-006, -2.892068e-006, 
    -4.248943e-006, -8.649007e-006, -9.309129e-006, -1.052668e-005, 
    -1.124293e-005, -6.105999e-006, -5.782645e-006, -4.737328e-006, 
    -4.922227e-006, -5.208824e-006, -4.163137e-006, -4.348904e-006, 
    -3.119185e-006, -2.548471e-006, -5.581478e-006, -8.563573e-006, 
    -6.552786e-006, -4.700943e-006, -1.760573e-006, 2.359347e-007, 
    2.099946e-006, 2.721076e-006, 2.531708e-006, 4.975995e-006, 
    5.624444e-006, 7.708246e-006, 1.068016e-005, 7.681299e-006, 
    4.446756e-006, 1.670545e-006, 5.571819e-007, 3.038585e-007, 
    -1.949196e-006, -4.407888e-006, -2.685189e-006, -4.879385e-006, 
    -5.129848e-006, -7.219984e-006, -5.065896e-006, -4.808106e-006, 
    -6.068127e-006, -2.815326e-006, -2.930563e-006, -2.293909e-006, 
    -7.961193e-006, -6.760532e-006, 1.333654e-006, 4.932161e-006, 
    2.922243e-006, 5.155678e-006, 6.136797e-006, 6.912647e-006, 
    3.084664e-006, 2.361834e-006, 2.454843e-006, 2.306948e-006, 
    1.939883e-006, -4.546109e-007, -1.912314e-006, -1.0853e-006, 
    -3.024192e-006, -2.019605e-006, 1.282121e-006, 7.980816e-007, 
    -1.248469e-006, -3.423789e-006, -6.339178e-007, 4.858772e-006, 
    6.493556e-006, 7.535764e-006, 7.5344e-006, 3.293157e-006, -1.822038e-006, 
    -5.023554e-006, -8.595733e-006, -1.025274e-005, -1.224702e-005, 
    -1.049836e-005, -1.06809e-005, -8.388361e-006,
  -4.340956e-006, -3.984198e-006, -3.093605e-006, -2.193575e-006, 
    -1.593431e-006, -1.182656e-006, -1.87767e-006, -6.409486e-006, 
    -8.302306e-006, -9.252875e-006, -8.742012e-006, -6.316603e-006, 
    -3.803149e-006, -2.04059e-006, -5.849943e-007, -9.027608e-007, 
    -3.996864e-006, -5.968907e-006, -5.09595e-006, -5.371372e-006, 
    -4.996111e-006, -3.687913e-006, -2.670165e-006, 5.96543e-007, 
    7.438157e-007, 9.064934e-009, -6.506889e-008, -3.83332e-007, 
    -3.454588e-007, -7.612007e-007, -4.811337e-006, -3.784894e-006, 
    -2.94795e-007, 2.413243e-006, 3.221135e-006, 4.22659e-006, 4.912913e-006, 
    5.289788e-006, 6.283944e-006, 6.415198e-006, 8.472553e-006, 
    1.083861e-005, 8.470688e-006, 4.85045e-006, 2.939501e-006, 2.059587e-006, 
    9.374089e-007, -1.03315e-006, -3.818423e-006, 9.443611e-007, 
    2.806759e-006, 4.432102e-006, 2.084671e-006, -1.31478e-006, 
    -3.420562e-006, -6.337094e-006, -7.105122e-006, -3.104407e-006, 
    3.176428e-007, -4.135291e-008, 2.19432e-006, 7.337952e-006, 8.40053e-006, 
    7.277726e-006, 6.404269e-006, 8.997944e-006, 6.700928e-006, 
    5.147111e-006, 2.689289e-006, 1.366061e-006, -2.471481e-006, 
    -1.96807e-006, -2.93925e-007, -3.096957e-007, -4.282847e-007, 
    -5.44017e-007, -3.103169e-007, 8.001925e-007, 2.239271e-006, 
    -7.849176e-007, -4.137804e-006, -1.523767e-006, 3.18835e-006, 
    5.979589e-006, 5.991635e-006, 2.269073e-006, -3.174693e-006, 
    -6.958842e-006, -7.510309e-006, -8.805591e-006, -7.132689e-006, 
    -7.102763e-006, -6.504481e-006, -5.067388e-006, -4.912417e-006, 
    -4.75968e-006,
  -1.831353e-006, -1.230091e-006, -7.287908e-007, -3.373871e-007, 
    -6.325542e-007, -3.53406e-007, -1.691405e-006, -2.675752e-006, 
    -5.897629e-006, -7.132316e-006, -5.456308e-006, -2.785027e-006, 
    -3.812214e-006, -3.852198e-006, -3.148119e-006, -2.024322e-006, 
    -2.441928e-006, -1.737973e-006, -2.27665e-006, -3.020589e-006, 
    -4.883856e-006, -2.874682e-006, -1.33241e-007, 2.650047e-006, 
    2.449255e-006, 2.267212e-006, 1.680354e-006, 1.192466e-006, 
    -1.886237e-007, -1.501292e-006, -1.982724e-006, 4.226963e-007, 
    2.799804e-006, 4.292776e-006, 3.659725e-006, 6.189942e-006, 
    4.933278e-006, 3.349905e-006, 5.682434e-006, 5.414337e-006, 
    7.313986e-006, 8.454299e-006, 3.385669e-006, 2.872446e-006, 
    5.091351e-009, 2.377605e-006, -3.439709e-008, 9.750329e-007, 
    3.456822e-006, 7.219489e-006, 8.186449e-006, 6.247188e-006, 
    -6.027512e-007, -3.965197e-006, -2.529348e-006, 2.076478e-006, 
    5.35947e-007, 3.065539e-006, 7.576498e-006, 8.785228e-006, 8.640563e-006, 
    6.773571e-006, 7.262206e-006, 6.907059e-006, 7.60518e-006, 5.19057e-006, 
    2.214685e-006, 1.03439e-006, 2.47981e-007, -8.836396e-007, 
    -2.952911e-007, 4.325066e-007, 3.069636e-007, 3.439686e-007, 
    7.748604e-007, 4.73236e-007, 1.310309e-006, 1.585856e-006, 1.580641e-006, 
    -2.070268e-006, -3.548586e-006, -6.55825e-006, -3.469489e-006, 
    -4.45023e-006, -5.536651e-006, -7.463123e-006, -9.63869e-006, 
    -8.411458e-006, -7.134304e-006, -5.779043e-006, -1.565119e-006, 
    -2.953783e-006, -3.941109e-006, -2.655635e-006, -1.33502e-006, 
    -2.376859e-006,
  1.683838e-007, -8.046618e-008, -2.369284e-007, -1.461555e-007, 
    -1.018242e-008, 1.16353e-007, -2.52699e-007, -1.852711e-006, 
    -9.775158e-007, -2.255166e-006, -1.799315e-006, -1.810739e-006, 
    -2.317131e-006, -5.524482e-006, -4.508843e-006, -3.190711e-006, 
    6.382652e-008, -8.948155e-007, -2.928822e-006, -2.460555e-006, 
    -3.568952e-006, -3.265466e-006, 3.977375e-007, 1.311302e-006, 
    1.138448e-006, 2.512088e-007, 3.666928e-007, 1.990547e-007, 
    -2.632537e-007, -5.625188e-007, 5.18188e-007, 1.472483e-006, 
    2.378225e-006, 1.72928e-006, 3.427764e-006, 5.114327e-006, 5.681688e-006, 
    6.859997e-006, 4.391745e-006, 6.816412e-006, 9.64726e-006, 6.296858e-006, 
    9.090945e-007, 1.250828e-006, -1.205628e-006, -4.672756e-006, 
    -5.675356e-006, -6.51454e-006, -1.2286e-006, 4.379079e-006, 
    2.542387e-006, -7.624476e-008, -2.932298e-006, 2.759076e-006, 
    2.988054e-006, 9.22133e-007, -1.279004e-007, 5.811202e-006, 
    8.882209e-006, 8.120387e-006, 3.885976e-006, 7.462999e-006, 5.74924e-006, 
    3.537534e-006, 1.932929e-006, -1.341105e-006, -2.463908e-006, 
    -1.011044e-006, -1.101072e-006, -2.679726e-007, -2.967772e-008, 
    -3.936384e-008, 4.547337e-007, 3.317991e-007, 7.562335e-008, 
    4.841636e-007, 3.849482e-008, 1.438831e-006, 3.024191e-006, 
    -2.752369e-006, -6.44823e-006, -8.652236e-006, -6.868566e-006, 
    -6.105131e-006, -6.347149e-006, -4.978603e-006, -7.514904e-006, 
    -3.025929e-006, -2.68432e-006, -1.150991e-006, -1.775722e-006, 
    -1.540035e-006, -1.126527e-006, -2.697107e-007, -4.569665e-008, 
    5.460033e-007,
  -8.215511e-007, -6.073465e-007, -4.197136e-008, 3.77496e-008, 
    -1.533577e-007, -6.974983e-007, -1.629939e-006, -1.636396e-006, 
    -1.572818e-006, -2.329548e-006, -5.235279e-007, -3.07833e-007, 
    -2.371024e-006, -6.109601e-006, -2.790615e-006, -6.42116e-007, 
    8.145971e-007, -2.047916e-006, -2.648681e-006, -2.932672e-006, 
    -2.167374e-006, -2.232691e-007, 1.711026e-006, 5.668653e-007, 
    -2.694651e-008, -1.85395e-007, -1.310061e-006, -1.85805e-006, 
    -1.370037e-006, 7.096678e-007, 9.427467e-007, 8.987884e-007, 
    1.136834e-006, 2.867729e-006, 5.406762e-006, 6.354476e-006, 
    5.144253e-006, 4.567454e-006, 5.11917e-006, 5.50809e-006, 2.221763e-006, 
    -5.149595e-007, -1.016136e-006, 4.334997e-007, -1.734745e-006, 
    -3.827612e-006, -3.787751e-006, -5.255764e-006, -5.739306e-006, 
    -3.775087e-006, -1.246604e-006, -2.513578e-006, -3.459925e-006, 
    -4.114334e-006, -1.980243e-006, -3.05387e-006, 8.431562e-007, 
    6.706019e-006, 3.933286e-006, -1.174336e-006, 1.681843e-006, 
    4.798174e-006, 1.621867e-006, -1.147639e-006, -1.544009e-006, 
    -2.492468e-006, -1.8357e-006, -1.975894e-006, -9.735431e-007, 
    -1.058479e-006, -1.283114e-006, -4.009653e-007, -7.167459e-007, 
    2.550582e-007, 1.88003e-007, 6.205091e-007, 1.663218e-006, 1.980985e-006, 
    4.540632e-006, -9.401887e-006, -8.078292e-006, -8.987884e-006, 
    -7.22309e-006, -6.319831e-006, -8.29262e-006, -4.211441e-006, 
    -1.723568e-006, 1.281624e-006, 8.776778e-007, 8.717234e-008, 
    1.101444e-007, -2.669731e-008, -7.949766e-007, -7.065591e-008, 
    -9.144351e-007, -6.364035e-007,
  -7.639328e-007, -5.776683e-007, -3.656994e-007, 2.268702e-007, 
    -2.807626e-007, -1.235058e-006, -3.778686e-007, -6.916628e-008, 
    -6.102026e-007, -1.03203e-006, -9.803723e-007, -6.869432e-007, 
    -9.494524e-007, -1.78193e-006, -3.191326e-007, -1.177068e-006, 
    -7.32889e-007, -1.119202e-006, -2.316758e-006, -3.167738e-006, 
    -1.254802e-006, 4.431849e-007, 1.040349e-006, 4.75593e-008, 4.69262e-007, 
    -1.422564e-006, -1.721705e-006, -1.771127e-006, -9.031346e-007, 
    2.841155e-007, 8.933247e-007, 3.702938e-007, 3.367662e-007, 
    1.112247e-006, 3.670528e-006, 3.058712e-006, 1.217052e-006, 
    2.389525e-006, 2.276525e-006, -1.391271e-006, -1.823158e-006, 
    -4.749125e-006, -1.181661e-006, -1.446035e-006, -2.865991e-006, 
    -2.85854e-006, -5.860255e-006, -1.143329e-005, -7.431085e-006, 
    -1.571079e-006, -1.730521e-006, -1.333654e-006, -2.626082e-006, 
    -3.685676e-006, -3.089508e-006, 1.753991e-006, 4.589432e-006, 
    2.390145e-006, -1.020109e-006, -9.870782e-007, 1.657754e-007, 
    -1.034396e-007, -1.713509e-006, -3.115212e-006, -2.527361e-006, 
    -3.16451e-006, -2.108639e-006, -2.492096e-006, -1.653408e-006, 
    -2.02991e-006, -1.305341e-006, -1.153102e-006, -5.823867e-007, 
    6.581331e-009, -5.985298e-007, 2.48477e-007, 6.927798e-007, 
    3.728271e-006, -7.62444e-007, -7.994971e-006, -5.208204e-006, 
    -4.509092e-006, -4.81382e-006, -2.388781e-006, -5.023802e-006, 
    -4.135072e-006, 7.820618e-007, 1.01688e-006, 7.241961e-007, 
    4.195917e-007, -6.31313e-007, -7.096678e-007, -2.132108e-006, 
    -1.78193e-006, -1.486639e-006, -3.479418e-007,
  -1.566857e-006, -1.216059e-006, 4.316369e-007, 6.046146e-007, 
    -1.281624e-006, -1.73524e-006, -7.146346e-007, 3.80104e-007, 
    -3.433476e-007, -9.0835e-007, -1.732757e-006, -1.598646e-006, 
    1.010794e-007, -2.035251e-006, -3.580377e-006, -4.489222e-006, 
    -1.75784e-006, 1.196315e-006, -1.379723e-006, -4.301473e-007, 
    1.533578e-006, 2.127886e-006, 3.976129e-007, -1.328681e-007, 
    -5.178163e-007, -1.256417e-006, -9.807454e-007, -5.399188e-007, 
    5.589181e-007, 4.188464e-007, 7.014723e-007, 1.070152e-006, 
    1.583373e-006, 1.765291e-006, 1.541028e-006, 2.771243e-006, 9.58393e-007, 
    7.722527e-007, -3.473212e-007, -4.14662e-006, -2.219404e-006, 
    7.943545e-007, 2.411132e-006, -2.864748e-006, -2.258394e-006, 
    -7.945298e-006, -1.064974e-005, -1.215364e-005, -7.011742e-006, 
    -5.59961e-006, -5.451588e-006, -5.230679e-006, -3.880883e-006, 
    1.212084e-006, 5.992006e-006, 6.785493e-006, 6.96443e-006, 1.487384e-006, 
    4.65413e-007, -1.664012e-008, -9.437399e-007, -1.540905e-006, 
    -2.972409e-006, -2.661347e-006, -1.89518e-006, -2.217665e-006, 
    -2.260133e-006, -2.305582e-006, -2.349541e-006, -2.567471e-006, 
    -1.659741e-006, -1.599267e-006, -1.224876e-006, -4.128865e-007, 
    -5.132207e-007, 4.749745e-007, 6.759665e-006, 6.612514e-006, 
    -3.885727e-006, -2.64657e-006, -2.612298e-006, -2.428269e-006, 
    -1.169617e-006, -1.118829e-006, -1.321857e-006, -1.295283e-006, 
    1.304223e-006, 6.428609e-007, -1.845256e-007, -2.558036e-007, 
    -1.581509e-006, -2.459313e-006, -2.732128e-006, -2.539779e-006, 
    -1.707176e-006, -1.46019e-006,
  -1.632794e-006, -1.234437e-006, -6.814796e-007, 1.421198e-006, 
    -1.32223e-006, -7.233275e-007, 2.090136e-006, 1.069407e-006, 
    8.850047e-007, -3.449618e-007, -9.239961e-007, -2.081941e-006, 
    -1.885121e-006, -4.307305e-006, -6.153185e-006, -5.49592e-006, 
    -6.429849e-006, -3.333515e-006, -2.465767e-006, -2.002344e-006, 
    1.828248e-006, 3.110617e-006, 3.515184e-006, 2.978246e-006, 
    3.774589e-006, 1.41114e-006, 4.727399e-007, 1.038362e-006, 3.601144e-008, 
    4.179783e-007, 1.871834e-006, 2.396231e-006, 4.528215e-006, 
    4.051004e-006, 5.406266e-006, 5.640586e-006, 2.603481e-006, 
    3.738578e-006, 3.687417e-006, 4.410371e-006, 1.581634e-005, 
    1.488241e-005, 8.539981e-006, 1.844517e-006, -1.170412e-005, 
    -2.369968e-005, -7.145856e-006, -1.03434e-005, -2.725174e-006, 
    -4.883608e-006, 4.878893e-007, 4.69834e-006, 8.711468e-006, 
    1.515622e-005, 1.82019e-005, 1.191422e-005, 6.048009e-006, 1.033397e-006, 
    -7.792069e-007, -1.450256e-006, -1.397977e-006, -1.335393e-006, 
    -1.395866e-006, -1.383325e-006, -2.145146e-006, -2.287825e-006, 
    -2.634897e-006, -2.641976e-006, -2.647192e-006, -2.807131e-006, 
    -1.852338e-006, -1.749893e-006, -1.653036e-006, -1.614353e-009, 
    1.757094e-007, 8.482362e-006, -1.273176e-006, -9.393934e-007, 
    1.772617e-006, 2.794217e-006, -3.079576e-007, -1.52948e-006, 
    -3.096959e-007, -2.476076e-007, 2.057602e-007, -1.119698e-006, 
    -3.69424e-007, 1.103927e-006, -1.107653e-006, -1.204759e-006, 
    -2.775713e-006, -2.834573e-006, -2.856056e-006, -2.312288e-006, 
    -1.422936e-006, -1.369913e-006,
  -1.064688e-006, -3.563864e-007, -1.351659e-006, -2.077222e-006, 
    -2.433732e-006, -3.033629e-006, 1.986449e-006, 7.091461e-006, 
    1.486018e-006, 7.003546e-007, -2.372017e-006, -3.224487e-006, 
    -3.615022e-006, -3.654633e-006, -9.821852e-006, -8.811181e-006, 
    -8.137151e-006, -9.245177e-006, -3.696852e-006, -7.889168e-006, 
    -7.197385e-006, -9.271025e-007, 4.499158e-006, 8.128336e-006, 
    9.899588e-006, 4.703551e-006, 1.827503e-006, 3.777321e-006, 
    1.812851e-006, 4.15792e-006, 5.244463e-006, 3.146876e-006, 3.042693e-006, 
    3.7464e-006, 9.128824e-006, 1.035531e-005, 1.704879e-005, 2.601147e-005, 
    1.531914e-005, 9.401887e-006, 1.961862e-005, 1.139082e-005, 
    5.577138e-006, 3.537163e-006, -1.720128e-005, -1.942192e-005, 
    -1.407029e-005, -9.414558e-006, 7.613002e-006, 2.249095e-005, 
    2.952702e-005, 2.775043e-005, 2.624144e-005, 2.031202e-005, 
    1.343762e-005, 8.053332e-006, 2.678235e-006, -8.22296e-007, 
    -9.644782e-007, -1.911695e-006, -1.295035e-006, -1.350293e-006, 
    -1.543512e-006, -1.632795e-006, -2.391512e-006, -2.405171e-006, 
    -2.81011e-006, -3.017113e-006, -2.453103e-006, -2.681215e-006, 
    -1.905734e-006, -2.180661e-006, -7.019689e-007, -8.111197e-007, 
    9.508185e-007, 4.296129e-006, -3.167739e-006, 3.089508e-006, 
    2.679852e-006, 1.854934e-005, 3.811841e-006, -1.168624e-006, 
    -2.893285e-008, -6.152936e-007, -8.656332e-007, -6.098301e-007, 
    -5.581724e-007, -4.4629e-007, -1.280009e-006, -1.461804e-006, 
    -2.502898e-006, -2.153963e-006, -2.477194e-006, -1.70519e-006, 
    -1.73611e-006, -1.481424e-006,
  2.236416e-007, -6.371492e-007, 7.948529e-007, 1.803289e-006, 
    -1.409899e-006, 3.976311e-009, 5.866212e-006, 7.357448e-006, 
    1.042461e-005, 7.337208e-006, 6.390119e-007, -1.719097e-006, 
    -4.253537e-006, -5.736201e-006, -8.893014e-006, -7.523966e-006, 
    -5.587313e-006, -9.717296e-006, -1.589469e-005, -1.207391e-005, 
    -9.842468e-006, -1.63056e-006, 2.782668e-006, 4.545102e-006, 
    9.184452e-006, 2.062445e-006, 6.045528e-006, 3.33786e-006, 9.452428e-006, 
    1.657642e-005, 7.341305e-006, 9.9505e-006, 7.731094e-006, 1.838927e-005, 
    2.026906e-005, 9.583891e-007, -8.857125e-006, -8.999683e-006, 
    -1.396114e-006, 1.34971e-005, 2.120336e-005, -9.240954e-006, 
    -1.852342e-006, 6.64244e-006, -8.6613e-006, 1.561282e-005, 2.812868e-005, 
    3.725849e-005, 4.001135e-005, 3.52487e-005, 2.429572e-005, 1.490377e-005, 
    8.113435e-006, 2.179419e-006, -1.173466e-007, -1.193583e-006, 
    -1.105045e-006, -1.471862e-006, -1.094987e-006, -1.665577e-006, 
    -9.698174e-007, -9.905548e-007, -1.417224e-006, -1.597404e-006, 
    -1.697739e-006, -2.00284e-006, -1.753122e-006, -2.431621e-006, 
    -1.76318e-006, -1.048793e-006, -2.192955e-007, 4.11148e-007, 
    6.801138e-007, 1.851841e-006, 4.310159e-007, 1.947952e-006, 
    1.062825e-006, 1.122442e-005, 4.6848e-006, 2.153305e-005, 1.36209e-005, 
    -2.647439e-007, -1.553198e-006, -2.528976e-006, -5.604078e-007, 
    -9.826072e-007, 1.605352e-006, 4.153326e-006, 6.14884e-006, 
    3.121669e-006, 3.715232e-006, 2.13782e-006, 1.417598e-006, 5.139659e-007, 
    -3.861896e-008, -7.809454e-007,
  1.064129e-005, 1.394823e-005, 1.320119e-005, 2.7063e-006, 6.801638e-006, 
    1.131842e-005, 7.969014e-006, 8.67949e-008, 1.57863e-005, 2.031016e-005, 
    3.629177e-006, -4.892536e-008, -1.628573e-006, -4.419686e-006, 
    -2.293411e-006, -5.630172e-007, 1.629196e-006, -6.808215e-006, 
    -2.90667e-005, -1.390974e-005, -5.592032e-006, -3.14576e-006, 
    5.664915e-007, -6.90663e-007, -4.17816e-006, -2.072629e-006, 
    -7.914998e-006, -1.979346e-005, 1.877484e-005, 2.986205e-005, 
    1.058715e-005, 1.178024e-005, 5.804497e-006, 1.555644e-005, 
    1.763031e-005, 2.774468e-006, 3.342211e-006, 1.664092e-006, 
    9.269272e-006, 2.15143e-005, 8.474541e-006, -7.371236e-006, 
    1.098848e-005, 2.609044e-005, 3.55122e-005, 4.534001e-005, 5.830961e-005, 
    6.379646e-005, 5.409345e-005, 3.931485e-005, 2.65417e-005, 1.589892e-005, 
    9.82595e-006, 3.356859e-006, 1.576046e-006, 1.509984e-007, 
    -3.062189e-007, -9.057421e-007, -6.955115e-007, -7.60456e-007, 
    -1.690039e-007, -8.441509e-007, -3.044804e-007, -7.635606e-007, 
    -5.811451e-007, -6.228688e-007, -1.046434e-006, -1.22351e-006, 
    -1.172473e-006, -7.078052e-008, 1.702458e-006, 6.719307e-006, 
    9.779011e-006, 1.211105e-005, 1.618514e-005, 4.843248e-006, 
    -1.552326e-006, 9.266536e-006, 1.070053e-005, 1.597318e-005, 
    3.867472e-006, -1.525133e-006, -8.382773e-006, -7.993853e-006, 
    -2.759447e-006, 3.376335e-007, 6.478156e-006, 1.270324e-005, 
    1.550205e-005, 1.039542e-005, 1.084693e-005, 8.390844e-006, 1.13563e-005, 
    9.674206e-006, 7.28555e-006, 1.074014e-005,
  1.299766e-005, 4.241467e-005, 1.896844e-005, -1.161831e-005, 
    -4.859765e-006, 3.306319e-006, 2.873072e-006, -7.482748e-006, 
    -2.816931e-006, 8.431452e-006, -2.859815e-007, 1.248716e-006, 
    -8.530924e-008, -2.469123e-006, 1.385559e-006, 5.701186e-006, 
    1.020294e-005, 1.531616e-005, 9.335577e-006, 1.043404e-005, 
    1.174709e-005, 5.550195e-006, 4.076712e-006, -2.144028e-006, 
    -5.607428e-006, -5.032744e-006, 3.066038e-006, 5.583461e-006, 
    2.292158e-005, 3.014096e-005, 9.368232e-006, -2.013519e-006, 
    4.839647e-006, 6.222966e-006, 8.556526e-008, 2.733243e-006, 
    7.765244e-006, 7.527065e-006, 1.055449e-005, -2.503904e-006, 
    -1.671302e-005, -1.167021e-005, -9.908283e-006, 3.623602e-006, 
    -1.401582e-006, -1.02807e-005, 5.150709e-006, 1.551423e-005, 
    2.103634e-005, 2.402552e-005, 3.070347e-005, 3.242679e-005, 
    3.737794e-005, 2.467148e-005, 1.975422e-005, 1.500162e-005, 
    1.162117e-005, 9.72785e-006, 7.211043e-006, 5.615999e-006, 5.623822e-006, 
    5.578993e-006, 5.250051e-006, 8.912508e-006, 8.940944e-006, 1.0535e-005, 
    1.124839e-005, 6.243339e-006, 1.731267e-006, 9.916475e-006, 
    6.509446e-006, 1.164911e-005, 1.517907e-005, 2.522704e-005, 
    -1.82775e-006, -6.35584e-006, -6.636983e-006, 9.504711e-006, 
    1.33009e-005, -1.177763e-005, -2.134715e-006, -1.280755e-006, 
    -1.779324e-006, -3.809233e-006, 4.974499e-007, 6.480892e-006, 
    7.376075e-007, -7.262453e-006, -6.392584e-007, 2.540401e-006, 
    8.900221e-006, 1.338472e-005, 6.420167e-006, 7.968411e-007, 
    6.304435e-006, 8.789204e-006,
  7.924558e-006, 9.955838e-006, -4.455447e-006, -6.005415e-006, 
    -1.101689e-006, 1.442968e-007, 4.90708e-006, 1.641114e-006, 
    -1.159745e-005, -1.613647e-005, -2.308736e-005, -2.167499e-006, 
    -3.319606e-006, -4.28607e-006, -2.106031e-006, 4.486863e-006, 
    1.503353e-005, 1.696857e-005, 1.746093e-005, 1.981841e-005, 
    1.667428e-005, 9.032956e-006, 4.807735e-006, 3.361492e-007, 
    4.779416e-006, -7.016337e-006, 3.272071e-007, 1.209677e-005, 
    2.14239e-005, 3.930107e-005, 1.715471e-005, 1.649372e-005, 7.358445e-006, 
    5.088732e-007, 5.099675e-006, 3.037363e-006, 9.484589e-006, 
    9.786963e-006, 5.622707e-006, -3.295645e-007, -5.945563e-006, 
    -4.278998e-006, -9.252253e-006, 3.430905e-007, -4.239511e-006, 
    -2.864289e-005, -1.112745e-005, 3.780675e-006, -4.259738e-006, 
    -2.123764e-005, -1.7053e-005, -1.523868e-005, -5.652546e-007, 
    5.890906e-007, -2.598761e-006, 8.381903e-008, 9.094052e-006, 
    1.001954e-005, 1.175714e-005, -3.741552e-006, -1.029422e-005, 
    1.275638e-005, 1.616577e-005, 2.286521e-005, 1.601651e-005, 
    1.743026e-005, 2.614657e-005, 1.053698e-005, 1.0759e-005, 1.631318e-005, 
    4.821646e-006, 1.08098e-005, -2.21518e-006, -1.975037e-005, 
    -5.258173e-005, -3.940203e-005, -1.78285e-005, -1.409414e-005, 
    -1.57586e-005, -1.075913e-005, -5.976482e-006, 1.687549e-007, 
    2.429759e-006, -5.530317e-006, -9.694486e-007, 9.287396e-006, 
    1.777458e-006, -7.791568e-006, -7.627532e-006, -1.978115e-007, 
    4.379326e-006, 5.036221e-006, 3.801659e-006, -1.032191e-005, 
    -6.666538e-006, 3.024565e-006,
  1.47571e-006, 2.471108e-006, 3.09795e-006, 6.945193e-007, -7.038068e-006, 
    -1.365232e-005, -1.352119e-005, -1.063533e-005, -3.210826e-006, 
    -7.415689e-006, -8.86706e-006, -9.99371e-007, 2.992772e-006, 
    3.445894e-007, 7.078052e-007, -8.37942e-007, 4.759058e-006, 
    6.887443e-006, 8.072333e-006, 1.764086e-005, 2.938298e-005, 
    2.427858e-005, 1.635862e-005, -4.513815e-006, 1.716246e-006, 
    1.216891e-005, 1.647e-005, 1.615151e-005, 2.889708e-005, 2.924961e-005, 
    1.791344e-005, 1.847706e-005, 2.5712e-006, 1.400473e-005, 2.35873e-005, 
    1.287783e-005, 1.426998e-005, 1.942527e-005, 1.527047e-005, 2.39869e-005, 
    8.604176e-006, -3.372879e-006, 3.690511e-007, 4.262234e-006, 
    5.629285e-006, 6.658709e-006, 2.632464e-005, 2.196506e-005, 
    5.964939e-006, -1.198414e-005, -1.320727e-005, -1.196815e-006, 
    2.897283e-006, 4.915397e-006, -2.784283e-006, -1.757344e-006, 
    5.699319e-006, 1.099221e-005, 6.276121e-006, 3.535548e-006, 
    6.322811e-006, 2.184548e-005, 2.250336e-005, 2.111346e-005, 
    1.905722e-005, 2.055553e-005, 1.602372e-005, 1.670668e-005, 
    2.283008e-005, 1.588278e-005, 4.927686e-006, -2.800921e-005, 
    -4.30615e-005, -3.891178e-005, -3.385656e-005, -3.04376e-005, 
    -2.011806e-005, -1.52301e-005, -1.188641e-005, -1.224056e-005, 
    -1.576158e-005, -1.177502e-005, -1.356142e-005, -9.856747e-006, 
    -4.884105e-006, -6.517395e-006, -8.064631e-006, -5.879501e-006, 
    -5.902722e-006, -3.87008e-006, -5.1445e-006, -1.165631e-005, 
    -2.859531e-006, -2.97216e-006, -1.149998e-006, 4.340462e-006,
  -1.4623e-006, -2.363076e-006, -3.153707e-006, -2.263362e-006, 
    -1.576915e-006, -1.454974e-006, -1.340111e-006, -3.705546e-006, 
    -2.652283e-006, -1.967947e-006, -3.447632e-006, -4.575899e-007, 
    8.575616e-007, 4.246955e-006, 1.39003e-006, 2.078091e-006, 2.404426e-006, 
    5.386894e-006, 1.112881e-005, 2.039609e-005, 2.540214e-005, 
    1.452317e-005, 9.628879e-006, -2.782042e-006, 1.202971e-005, 
    2.894861e-005, 2.09144e-005, 1.329395e-005, 1.687581e-005, 2.674956e-005, 
    1.510717e-005, 5.778798e-006, -2.057453e-005, 1.71747e-005, 
    2.684083e-005, 1.857305e-005, 1.709983e-005, 1.993999e-005, 
    1.933127e-005, 1.431107e-005, 1.865003e-006, -1.007269e-005, 
    -1.175503e-005, 7.36217e-006, 6.066264e-006, 6.424758e-006, 
    7.227063e-007, -1.042709e-005, -9.386989e-006, -2.732129e-006, 
    6.269045e-006, 4.128116e-006, 4.577138e-006, 2.48216e-006, 
    -3.888457e-006, 1.523022e-006, 8.934861e-006, 6.974735e-006, 
    2.061699e-006, 4.037965e-006, 8.681292e-006, 1.415424e-005, 1.18571e-005, 
    9.579831e-006, 9.641673e-006, 7.220231e-006, 1.794385e-005, 
    2.696899e-005, 1.855182e-005, 4.367532e-006, -4.24149e-006, 
    -4.652229e-005, -5.210712e-005, -2.176823e-005, -1.843895e-005, 
    -2.584842e-005, -1.423707e-005, -1.189498e-005, -1.826907e-005, 
    -1.278743e-005, -1.259272e-005, -1.408371e-005, -1.049377e-005, 
    -4.619732e-006, -5.82238e-006, -3.629178e-006, -3.666059e-006, 
    -4.1044e-006, -3.254289e-006, -2.718717e-006, -3.242617e-006, 
    -8.6387e-006, -6.700307e-006, -3.861513e-006, -1.07487e-006, 
    -1.477078e-006,
  -6.901721e-007, -2.458692e-007, -1.671414e-007, -6.407499e-008, 
    -1.04184e-007, -1.978129e-007, -7.115305e-008, -5.786618e-008, 
    -4.979471e-008, -1.814217e-007, -3.546353e-006, -7.102886e-008, 
    3.514191e-008, 2.609814e-006, 4.679213e-006, 9.18371e-006, 2.710894e-006, 
    3.185867e-006, 5.338341e-006, 2.299882e-005, 9.827814e-006, 6.31313e-006, 
    8.491188e-007, -1.70985e-007, 8.43071e-006, 2.531521e-005, 1.820326e-005, 
    2.072217e-005, 8.666513e-006, 6.167094e-006, 5.936992e-006, 9.64589e-006, 
    1.278532e-005, 2.001648e-005, 1.361556e-005, 9.75802e-006, 7.665774e-006, 
    -7.867857e-007, -2.258894e-006, -5.375718e-006, -9.724121e-006, 
    -1.836469e-005, -1.056617e-005, 5.878632e-006, 6.509574e-006, 
    4.892303e-006, -6.430968e-006, -1.197755e-005, -1.091361e-005, 
    -2.781177e-006, -3.01165e-006, -4.614514e-006, -5.558381e-006, 
    -3.661216e-006, -3.178866e-008, -9.103369e-007, 2.823646e-006, 
    1.340857e-006, -1.582504e-006, 9.564064e-007, 7.095432e-007, 
    -1.029671e-006, -2.675504e-006, -4.128243e-006, -6.075451e-006, 
    -1.009107e-005, -6.116556e-006, 2.452297e-005, 6.865463e-006, 
    1.592698e-005, 4.103782e-006, -1.560835e-005, -1.223249e-005, 
    -6.491071e-006, -1.030365e-005, -1.761864e-005, -1.886574e-005, 
    -1.549584e-005, -1.143999e-005, -1.15751e-005, -1.045888e-005, 
    -7.164603e-006, -4.846229e-006, -3.19158e-006, -3.162771e-006, 
    -2.109135e-006, -2.348423e-006, -2.049407e-006, -1.378357e-006, 
    -1.34334e-006, -4.978228e-007, -5.554408e-007, -2.341221e-006, 
    -1.34098e-006, 5.026659e-007, -3.052255e-007,
  -1.301244e-006, -6.693105e-007, -1.029546e-006, -7.264316e-008, 
    -7.313987e-008, 7.450573e-010, -1.452863e-008, -2.856056e-009, 
    4.221996e-009, 6.705522e-009, 1.812975e-008, 1.164774e-007, 
    -1.538545e-007, -8.779273e-008, 1.951183e-006, 6.511311e-006, 
    1.13907e-005, 8.001429e-006, 8.366384e-006, 6.990758e-006, 1.154964e-005, 
    1.109279e-005, 9.037802e-006, 5.747253e-006, 1.513822e-005, 
    4.765516e-006, 9.311989e-007, 6.704155e-006, -1.169119e-006, 
    1.288578e-006, 7.368749e-006, 1.157721e-005, 2.286124e-005, 3.08053e-005, 
    2.466328e-005, 1.227098e-005, -2.39275e-006, -7.780021e-006, 
    -5.763271e-006, -4.874419e-006, -3.707908e-006, -4.028647e-006, 
    -5.266691e-006, -5.816171e-006, -7.508694e-006, -5.283953e-006, 
    -5.108741e-006, -1.192018e-005, -1.374707e-005, -1.538284e-005, 
    -1.042585e-005, -6.924072e-006, -6.120155e-006, -5.198146e-006, 
    -4.19418e-006, -1.520415e-006, 4.508838e-007, 1.505141e-006, 
    -1.033147e-006, -2.458816e-006, -1.006325e-006, -1.334523e-006, 
    -1.590327e-006, -6.768853e-007, -1.154964e-006, -3.648674e-006, 
    -1.573066e-005, -1.499058e-006, -1.271546e-007, 1.797081e-006, 
    -1.820177e-006, 4.235902e-006, -2.304958e-006, 2.084795e-006, 
    1.935288e-006, -7.042789e-006, -1.164625e-005, -1.006114e-005, 
    -9.256728e-006, -8.297338e-006, -7.120769e-006, -5.64754e-006, 
    -5.056461e-006, -3.14936e-006, -1.49707e-006, -1.122678e-006, 
    -1.752625e-006, -2.070144e-006, -1.976267e-006, -2.522394e-006, 
    -1.55891e-006, -6.036212e-007, -1.090517e-006, -2.54636e-006, 
    -1.158814e-006, -1.012782e-006,
  -1.704817e-006, -1.155833e-006, -1.152605e-006, -9.549161e-007, 
    -7.752329e-007, -3.652026e-007, -2.918144e-008, -4.221996e-008, 
    -3.72529e-009, -2.483527e-009, 2.438823e-007, 1.627952e-007, 
    8.468827e-008, -5.153318e-008, -1.663963e-007, 1.149128e-006, 
    1.8167e-006, 4.003693e-006, 1.463033e-005, 9.52656e-006, 1.000601e-005, 
    1.427916e-005, 6.873161e-007, 3.001333e-007, 1.650067e-005, 1.76503e-005, 
    2.108217e-005, 4.292153e-006, 4.502512e-006, 1.468261e-006, 
    6.303067e-006, 1.049849e-005, 1.478319e-005, 1.91136e-005, 9.069718e-006, 
    1.76087e-005, 6.924201e-006, 5.292764e-006, -1.53693e-006, 
    -1.176806e-005, -3.297504e-006, -2.881636e-006, -1.641238e-006, 
    -4.009284e-006, -9.853891e-006, -6.370121e-006, -1.022467e-006, 
    -4.322206e-006, -9.242074e-006, -1.149091e-005, -9.043515e-006, 
    -6.031494e-006, -3.601363e-006, -1.860037e-006, -3.295765e-006, 
    -3.30806e-007, -4.336234e-007, -4.277881e-007, 8.607904e-007, 
    -1.398847e-006, -1.143788e-006, 3.053492e-007, 5.215497e-009, 
    1.204512e-007, 3.694245e-007, -2.34209e-006, -4.269306e-006, 
    -1.450007e-006, -4.146241e-007, 8.302432e-007, 4.79867e-006, 
    1.718539e-005, 7.955859e-006, 8.08189e-006, 1.451001e-006, 
    -9.323194e-007, 7.153794e-007, 5.47928e-006, 2.675752e-006, 
    2.825756e-006, 1.511224e-006, -4.18735e-006, -5.19889e-006, 
    -3.187606e-006, -1.597902e-006, -1.331915e-006, -9.883197e-007, 
    -2.550086e-006, -2.268577e-006, -1.639501e-006, -2.57492e-006, 
    -7.43692e-007, 6.581331e-009, -2.07002e-007, -1.433864e-006, 
    -1.816203e-006,
  -2.628317e-006, -3.866355e-006, -2.093489e-006, -1.479809e-006, 
    -2.209966e-006, -1.101444e-006, -7.208437e-007, -5.65499e-007, 
    -4.010896e-007, -1.580765e-007, -1.937151e-008, 2.086163e-008, 
    4.35859e-008, 4.755954e-008, 1.532336e-007, 1.280258e-007, 2.539406e-007, 
    9.586413e-007, 5.089741e-006, 1.472607e-006, 3.570071e-007, 
    1.285523e-005, 5.858637e-006, 2.187118e-006, 3.740935e-006, 
    1.489557e-005, 1.349735e-005, -7.085626e-006, -4.622212e-006, 
    1.67526e-006, 5.089243e-006, 6.599103e-006, 8.763622e-006, 7.518877e-006, 
    5.915761e-006, 1.046955e-005, 8.930634e-006, 1.310668e-005, 
    6.986906e-006, -4.102043e-006, -3.307687e-006, -7.794551e-007, 
    -6.184018e-008, 3.637124e-007, -9.273499e-007, -2.476076e-006, 
    -1.423806e-006, -2.098568e-008, -7.150084e-007, -7.185216e-006, 
    -6.984795e-006, -6.580975e-006, -4.993379e-006, -1.882141e-006, 
    -1.332908e-006, -1.996631e-006, -1.438955e-006, -1.139815e-006, 
    -2.068782e-007, 2.816323e-007, 5.338343e-007, 2.142042e-007, 
    1.187746e-006, 1.140684e-006, -3.815939e-007, -1.040349e-006, 
    -2.127141e-006, -9.374071e-007, 1.710778e-006, 3.372877e-006, 
    6.143004e-006, 1.214445e-006, -7.41953e-007, 3.959238e-006, 
    2.532452e-006, -5.128109e-006, -1.74965e-006, -8.050374e-007, 
    2.474586e-006, 1.142398e-007, -3.128749e-006, -1.844019e-006, 
    -5.080674e-006, -6.645174e-006, -6.861992e-007, -7.847939e-008, 
    -2.163772e-006, -1.911447e-006, -1.350293e-006, -1.219535e-006, 
    -2.157191e-006, -2.102926e-006, -5.512188e-007, -1.015638e-006, 
    -2.007187e-006, -2.110749e-006,
  -2.664948e-006, -5.99958e-006, -6.270285e-006, -5.616248e-006, 
    -2.96769e-006, -3.258263e-006, -3.110741e-006, -2.489487e-006, 
    -2.983212e-006, -2.366304e-006, -1.524886e-007, -3.551443e-008, 
    -7.400911e-008, -4.435578e-007, -9.665886e-007, -2.060086e-007, 
    -1.23928e-007, 1.77572e-008, -7.325164e-007, -9.038799e-007, 
    -1.461558e-007, -2.158806e-006, -2.705057e-006, 1.949593e-008, 
    3.491823e-007, 4.639227e-006, 8.972736e-006, 8.789822e-006, 
    6.729861e-006, -2.930683e-006, 5.893784e-006, 7.473056e-006, 
    7.765368e-006, 2.203635e-006, 3.249696e-006, 8.451567e-006, 
    1.223658e-005, 8.932999e-006, 1.0873e-005, 9.879222e-006, 9.059037e-006, 
    4.92148e-006, 2.218037e-006, 1.734992e-006, 3.178866e-008, -2.05636e-006, 
    -2.401943e-006, 8.828938e-007, 2.261128e-006, -3.228213e-006, 
    -5.940719e-006, -3.716723e-006, -4.289175e-006, -2.597521e-006, 
    -2.422061e-006, -1.149127e-006, -2.554307e-006, -1.704197e-006, 
    6.44477e-008, 4.599497e-007, 8.903444e-007, -5.463789e-009, 
    7.127721e-007, 1.284728e-006, -8.0218e-008, -8.951872e-007, 
    -1.773237e-007, 2.602985e-006, -8.88358e-007, 1.342098e-006, 
    6.835038e-006, 1.592809e-006, -4.414469e-007, 2.781177e-006, 
    1.682465e-006, -2.934659e-006, -4.800037e-006, -3.869456e-006, 
    -1.99303e-007, -2.123539e-006, -4.203863e-006, -3.475074e-006, 
    -4.097074e-006, -6.443632e-006, -2.727036e-006, -1.156952e-006, 
    -2.345318e-006, -2.535681e-006, -1.908715e-006, -4.224476e-007, 
    -8.378174e-007, -1.706183e-006, -1.718104e-006, -1.847247e-006, 
    -5.057578e-006, -2.72654e-006,
  -4.48885e-006, -2.249082e-006, -1.686312e-007, 9.375253e-008, 
    -2.689667e-007, -1.999612e-006, -2.98818e-006, -2.613415e-006, 
    -3.049399e-006, -3.156438e-006, -1.648068e-006, -8.528431e-007, 
    -8.333475e-007, -2.53568e-007, -2.121304e-006, -1.499429e-006, 
    -1.368423e-006, -1.683831e-007, -8.431573e-008, -1.801426e-006, 
    -2.151728e-006, -8.561958e-007, -2.492218e-007, 2.432616e-007, 
    3.331652e-007, 1.399343e-006, 2.578025e-006, 3.268196e-006, 
    2.854442e-006, 6.494174e-006, 8.748226e-006, 6.093331e-006, 
    7.733577e-006, 8.355577e-006, 2.704932e-006, -1.437216e-006, 
    4.693495e-006, 1.052916e-005, 1.415933e-005, 1.669849e-005, 1.50077e-005, 
    1.725517e-005, 1.173131e-005, 5.101538e-006, 7.10773e-006, 6.084891e-006, 
    4.277999e-006, 5.522867e-006, 3.440429e-006, 9.17913e-007, 
    -2.701208e-006, -2.800798e-006, -2.028546e-006, 3.72529e-008, 
    9.477135e-007, 2.806013e-006, 9.801242e-007, -7.713843e-007, 
    -8.506049e-008, 1.631057e-006, 1.558909e-006, 1.731143e-006, 
    1.080086e-006, 1.145278e-006, 1.28746e-006, -2.406537e-007, 
    -1.993279e-006, -1.195445e-006, 5.411603e-007, -1.656141e-006, 
    -1.68875e-008, 1.546616e-006, -1.481796e-006, 1.267717e-006, 
    2.65489e-006, 1.098961e-006, 2.160596e-008, 6.797418e-007, 3.274654e-006, 
    -5.720794e-007, -4.95054e-006, -5.064903e-006, -3.355242e-006, 
    -1.575925e-006, -3.411871e-006, -6.337217e-006, -5.313133e-006, 
    -3.613035e-006, -3.233179e-006, -1.105915e-006, -1.22649e-006, 
    -2.437209e-006, -1.530101e-006, -1.128142e-006, -2.422059e-006, 
    -3.754472e-006,
  -7.110337e-006, -3.955029e-007, -3.388768e-007, -1.057486e-006, 
    -1.998867e-006, -3.282105e-006, -5.045781e-006, -1.969561e-006, 
    -8.672478e-007, -1.144409e-006, -1.931439e-006, -7.269407e-006, 
    -6.393591e-006, -3.094226e-006, -4.716217e-007, -1.390402e-006, 
    -2.270316e-006, -1.836568e-006, -6.334235e-007, -1.045441e-006, 
    -2.293537e-006, -2.507493e-006, -9.30329e-007, -4.156184e-007, 
    1.555929e-007, 3.851951e-007, 6.38639e-007, 1.795838e-006, 1.972914e-006, 
    1.913806e-006, 3.268073e-006, 4.15941e-006, 2.611678e-006, 1.314284e-006, 
    6.542832e-007, -1.779074e-006, -4.779919e-006, -4.185364e-006, 
    -8.805328e-007, 6.66752e-006, 1.56307e-005, 1.97197e-005, 1.909299e-005, 
    1.765129e-005, 1.512244e-005, 1.259931e-005, 9.364634e-006, 
    4.692003e-006, 4.56224e-006, 3.878275e-006, 4.571179e-006, 7.775925e-007, 
    3.700479e-007, -1.703702e-007, -4.464127e-007, 1.502522e-007, 
    3.088639e-006, 2.46639e-006, 2.304712e-006, 3.788124e-006, 2.86388e-006, 
    2.29304e-006, 1.773735e-006, 2.602737e-007, 6.109476e-007, 
    -3.467003e-007, -2.534316e-006, -2.263362e-006, -9.235009e-007, 
    3.483396e-006, 4.500274e-006, 4.736336e-006, 3.535424e-006, 
    2.129873e-006, 1.01862e-006, 1.570825e-007, -2.143161e-006, 
    -1.874443e-006, -3.517544e-006, -4.571553e-006, -6.223469e-006, 
    -5.471456e-006, -7.372846e-006, -6.354599e-006, -4.881869e-006, 
    -5.476673e-006, -9.112557e-006, -7.593631e-006, -3.338233e-006, 
    -1.57977e-006, -6.246082e-007, -1.808003e-007, -2.109012e-006, 
    -4.487112e-006, -5.877267e-006, -5.343681e-006,
  -1.190856e-007, -2.625093e-007, -4.496425e-006, -3.75323e-006, 
    -2.914421e-007, -1.89431e-006, -3.851825e-006, -1.327445e-006, 
    -9.479618e-007, -1.285225e-007, 1.211588e-006, 2.279876e-007, 
    -2.375617e-006, -3.321096e-006, -3.051013e-006, 3.214927e-007, 
    -2.445031e-007, -1.988436e-006, -2.191216e-006, -1.022468e-006, 
    -1.408035e-006, -2.6308e-006, -3.077959e-006, -2.102678e-006, 
    -1.02818e-006, -8.032966e-007, -1.003221e-006, -4.361073e-007, 
    -2.900761e-007, 4.843059e-009, 1.775846e-006, 1.747534e-006, 
    5.081292e-007, 5.883485e-007, -1.288703e-006, -2.662589e-006, 
    -4.014746e-006, -2.157565e-006, -4.381935e-006, -8.417916e-006, 
    -5.389629e-006, -2.512956e-006, -2.296001e-007, 3.797315e-006, 
    4.951034e-006, 7.685769e-006, 8.088478e-006, 9.108957e-006, 
    9.125099e-006, 3.939247e-006, 1.315897e-006, 1.221895e-006, 
    2.415476e-006, 7.124494e-006, 4.000962e-006, 2.297635e-006, 
    5.268059e-006, 5.594018e-006, 3.273908e-006, 4.230189e-006, 
    2.596278e-006, 4.088133e-006, 2.217541e-006, 1.361966e-006, 
    -1.918525e-007, 7.013477e-007, 2.060087e-007, -9.194018e-007, 
    5.08875e-007, -4.959602e-007, -6.793689e-007, -1.077602e-006, 
    -1.248221e-006, -8.588031e-007, -8.715942e-007, -1.743807e-006, 
    -1.88686e-006, -4.703797e-007, -4.056856e-007, -1.400338e-006, 
    -2.457946e-006, -3.523381e-006, -3.726407e-006, -4.030393e-006, 
    -2.337496e-006, -2.657496e-006, -3.167734e-007, -7.034578e-007, 
    -2.544366e-007, -3.290734e-008, -1.483913e-007, 7.917497e-007, 
    1.517437e-007, -7.500239e-007, -1.508743e-006, -6.904211e-007,
  3.69971e-006, 4.021947e-006, 2.553686e-006, 2.785649e-006, 3.099069e-006, 
    1.910452e-006, 4.78949e-007, -1.462425e-006, -1.857677e-006, 
    -7.496528e-007, 6.971259e-007, 7.064391e-007, -7.140143e-007, 
    6.162873e-007, 1.066799e-006, 4.233179e-007, 1.182408e-006, 
    9.736668e-007, -9.83473e-008, -4.624335e-007, -1.392018e-007, 
    -4.644198e-008, -6.861983e-007, -1.171231e-006, -2.367049e-006, 
    -2.707789e-006, -1.851718e-006, 5.52709e-007, 1.050408e-006, 
    -1.177937e-006, 3.501737e-008, -5.108614e-007, -1.721706e-006, 
    -2.307941e-006, -2.278015e-006, -2.365186e-006, -4.092353e-006, 
    -3.843383e-006, -2.890081e-006, -1.223758e-006, -2.037112e-006, 
    -4.289068e-007, 3.495315e-006, 2.80415e-006, 2.004206e-006, 
    2.655514e-006, 3.331279e-006, 3.971287e-006, 2.180415e-006, 
    4.599497e-007, 1.617522e-006, 2.684319e-006, 1.566357e-006, 
    3.891189e-006, 4.073478e-006, 3.075602e-006, 3.268695e-006, 
    5.404152e-006, 8.205079e-006, 5.0772e-006, 2.776087e-006, 4.624948e-006, 
    6.580478e-006, 6.658709e-006, 5.030384e-006, 6.575137e-007, 
    2.032775e-007, -9.16416e-008, -8.299949e-007, -2.520283e-006, 
    -2.273793e-006, 4.94967e-007, -8.856259e-007, -2.363697e-006, 
    -2.431247e-006, -6.587579e-007, 3.741559e-006, 7.195522e-006, 
    5.295875e-006, 3.200272e-006, 3.320849e-006, 3.271176e-006, 
    5.729489e-007, -5.489856e-007, -7.3314e-007, -2.267338e-006, 
    -3.065292e-006, -6.870687e-007, 1.201406e-006, 4.082547e-006, 
    4.584963e-006, 3.255533e-006, 4.212558e-006, 3.343075e-006, 
    2.585102e-006, 2.136454e-006,
  5.205475e-006, 5.916754e-006, 4.999587e-006, 4.543115e-006, 4.806492e-006, 
    5.388882e-006, 2.580135e-006, 2.261258e-007, -4.195917e-007, 
    -6.187711e-007, 1.244494e-006, 1.742816e-006, -3.299374e-007, 
    1.587596e-006, 2.344822e-006, 1.112621e-006, 1.047429e-006, 
    1.152728e-006, 9.063633e-007, 1.659e-007, -3.891691e-007, -8.320058e-009, 
    -9.69444e-007, -1.758586e-006, -7.112831e-007, 7.947283e-007, 
    7.222097e-007, -2.473598e-007, -1.328687e-006, -9.007754e-007, 
    -3.352761e-008, 2.889088e-006, 1.15695e-006, 1.568596e-006, 
    2.012899e-006, 1.00322e-006, 1.187997e-006, 2.103423e-006, 1.088158e-006, 
    1.336261e-006, 3.098199e-006, 6.286056e-006, 7.685769e-006, 
    7.775052e-006, 6.655602e-006, 2.874931e-006, 2.376488e-006, 
    5.954505e-006, 5.475806e-006, 2.445031e-006, 3.578014e-006, 
    4.065907e-006, 1.388416e-006, 2.977129e-006, 1.865872e-006, 
    2.474586e-006, 4.259371e-006, 7.100403e-006, 1.084444e-005, 
    1.010063e-005, 5.935999e-006, 7.221352e-006, 1.169095e-005, 
    1.096651e-005, 5.881984e-006, -2.602737e-007, -1.942118e-006, 
    -7.969629e-007, -5.991515e-007, -4.764643e-007, -2.02399e-008, 
    1.001856e-006, 3.270432e-006, 5.013248e-006, 4.785012e-006, 
    5.343803e-006, 8.09108e-006, 8.640935e-006, 8.565061e-006, 7.410224e-006, 
    3.491466e-006, 4.496673e-006, 3.486373e-006, 1.152359e-006, 
    -6.961345e-007, -3.568857e-007, 2.678109e-006, 2.013272e-006, 
    1.829369e-006, 5.451366e-007, 4.254405e-006, 5.142017e-006, 5.78873e-006, 
    5.557635e-006, 4.606198e-006, 4.174188e-006,
  3.492212e-006, 5.272774e-006, 6.459159e-006, 4.380199e-006, 1.322354e-006, 
    1.175329e-006, 1.282866e-006, 1.952796e-006, 7.224589e-007, 
    4.146001e-006, 5.072108e-006, 4.698337e-006, 5.366528e-006, 
    3.477309e-006, 1.931439e-006, 1.61392e-006, 9.275973e-007, 1.364823e-006, 
    1.400336e-006, 8.761881e-007, 9.403875e-007, 5.810216e-007, 
    2.004199e-007, 3.986133e-008, 1.50241e-006, 2.398963e-006, 1.844515e-006, 
    1.544133e-006, 2.553438e-006, 4.684677e-006, 3.715728e-006, 
    2.425786e-006, 4.007792e-006, 4.359212e-006, 3.248952e-006, 
    1.633167e-006, 4.899503e-006, 3.481284e-006, 3.070632e-006, 
    3.685802e-006, 2.553936e-006, 3.035491e-006, 4.87951e-006, 8.334715e-006, 
    9.722884e-006, 7.254133e-006, 4.937623e-006, 5.368018e-006, 
    5.303697e-006, 4.835178e-006, 4.893416e-006, 4.288304e-006, 
    3.342704e-006, 3.020592e-006, 1.638509e-006, 2.908208e-006, 
    9.204945e-006, 1.016917e-005, 9.238596e-006, 1.22952e-005, 1.594139e-005, 
    1.648565e-005, 1.085375e-005, 5.197151e-006, 1.717608e-006, 
    -2.017869e-007, -8.297466e-007, -4.718713e-007, 1.820426e-007, 
    1.952922e-006, 3.360834e-006, 3.001218e-006, 3.298248e-006, 
    3.228957e-006, 5.737194e-006, 8.189181e-006, 9.082009e-006, 
    8.969382e-006, 7.454804e-006, 6.08315e-006, 5.308539e-006, 5.871803e-006, 
    6.483249e-006, 5.800895e-006, 3.84984e-006, 5.410733e-006, 3.566591e-006, 
    1.860164e-006, 3.191704e-006, 2.848607e-006, 3.853071e-006, 
    2.083929e-006, 1.643351e-006, 3.511333e-006, 5.16052e-006, 2.45149e-006,
  2.582867e-006, 3.647185e-006, 5.471084e-006, 2.802288e-006, 2.116958e-006, 
    9.741634e-007, 8.491188e-007, 2.664452e-006, 3.790979e-006, 
    4.128367e-006, 3.974512e-006, 5.709628e-006, 6.112579e-006, 
    6.089234e-006, 3.327677e-006, 1.857181e-006, 9.956457e-007, 
    4.811827e-007, 1.629443e-006, 1.586477e-006, 7.125254e-007, 
    8.912139e-007, 1.164402e-006, 1.412381e-006, 2.081197e-006, 
    2.408151e-006, 2.061079e-006, 2.093862e-006, 2.532577e-006, 
    3.459802e-006, 2.234926e-006, 1.045937e-006, 7.78834e-007, 1.578283e-007, 
    1.829614e-006, 2.227725e-006, 2.669667e-006, 4.739562e-006, 
    4.866099e-006, 1.865377e-006, 2.350409e-006, 1.591818e-006, 
    1.073131e-006, 1.055994e-006, 2.095849e-006, 1.158316e-006, 
    1.566361e-006, 8.231655e-007, -9.785072e-008, 4.831691e-007, 
    1.057484e-006, 2.895795e-007, 6.935243e-007, 3.076218e-006, 
    3.247835e-006, 4.43657e-006, 6.975359e-006, 8.717921e-006, 9.134041e-006, 
    1.042597e-005, 1.320168e-005, 1.242608e-005, 8.561212e-006, 
    5.972262e-006, 3.85642e-006, 1.878912e-006, 2.161414e-006, 2.000232e-006, 
    1.47422e-006, 4.073358e-006, 3.825874e-006, 3.592547e-006, 3.371511e-006, 
    4.716217e-006, 2.962475e-006, 1.629565e-006, 3.09733e-006, 4.546469e-006, 
    2.895791e-006, 9.765226e-007, 2.991408e-006, 5.177035e-006, 
    4.464266e-006, 3.474455e-006, 4.444395e-006, 7.310759e-006, 
    5.708138e-006, 1.887107e-006, -4.188478e-007, 2.510227e-006, 
    4.908317e-006, 3.190464e-006, 1.390032e-006, 6.886803e-007, 
    2.601988e-006, 3.633399e-006,
  1.034141e-006, 5.878501e-007, 2.384682e-006, 3.226723e-006, 2.274041e-006, 
    2.258023e-006, 1.154964e-006, 9.182841e-007, 1.538918e-006, 
    2.916655e-006, 3.625577e-006, 4.166364e-006, 4.585212e-006, 
    5.214537e-006, 5.078067e-006, 4.632648e-006, 5.159527e-006, 
    4.652018e-006, 3.319481e-006, 2.150362e-006, 2.963345e-006, 
    4.392738e-006, 5.478909e-006, 4.685297e-006, 3.834937e-006, 
    4.117936e-006, 4.834683e-006, 5.190075e-006, 4.332388e-006, 
    2.548595e-006, 1.356006e-006, 5.650018e-007, 6.798655e-007, 
    1.749148e-006, 2.436464e-006, 2.684072e-006, 3.427888e-006, 
    3.478924e-006, 1.90325e-006, 1.482293e-006, 1.168126e-006, 2.342463e-006, 
    2.66681e-006, 2.621609e-006, 3.649418e-006, 3.605957e-006, 3.60012e-006, 
    2.455463e-006, 3.760051e-007, 2.508368e-007, 5.006787e-007, 
    1.888729e-007, 4.646681e-007, 2.160918e-006, 4.362564e-006, 
    3.422796e-006, 1.999488e-006, -1.647944e-006, -3.418572e-007, 
    2.059589e-006, 2.84339e-006, 2.281988e-006, 2.677491e-006, 3.468867e-006, 
    3.414725e-006, 3.309672e-006, 3.045798e-006, 2.983212e-006, 3.64917e-006, 
    3.69437e-006, 3.768379e-006, 4.789854e-006, 4.837166e-006, 3.137191e-006, 
    1.029422e-006, 6.21254e-007, 1.159558e-006, 2.264605e-006, -1.78441e-007, 
    -1.383076e-006, 2.75001e-006, 4.815558e-006, 5.117183e-006, 
    3.581867e-006, -1.246735e-007, -1.615161e-006, -2.640732e-006, 
    -1.17594e-007, 2.396355e-006, 3.153087e-006, 5.104517e-006, 
    4.112846e-006, 1.600509e-006, 1.170238e-006, 1.643473e-006, 2.004206e-006,
  -1.321981e-006, -1.542023e-006, -8.569405e-007, -9.436153e-007, 
    -1.515571e-006, -5.338334e-007, 1.334647e-006, 3.494695e-006, 
    6.287546e-006, 5.899743e-006, 2.730141e-006, 1.693888e-006, 
    2.657001e-006, 3.820905e-006, 4.771104e-006, 5.45842e-006, 5.258248e-006, 
    4.268314e-006, 4.098192e-006, 4.549075e-006, 4.742543e-006, 
    4.824003e-006, 5.107497e-006, 4.622712e-006, 4.328167e-006, 
    4.834432e-006, 5.789101e-006, 5.71919e-006, 5.076826e-006, 3.368657e-006, 
    2.21158e-006, 2.79434e-006, 3.904974e-006, 3.827611e-006, 3.113101e-006, 
    2.153093e-006, 1.792238e-006, 1.211837e-006, 1.767401e-006, 
    1.432746e-006, 1.819183e-006, 2.03078e-006, 2.357985e-006, 2.967069e-006, 
    3.012642e-006, 4.270176e-006, 4.805376e-006, 4.27241e-006, 3.736094e-006, 
    2.586718e-006, 9.540472e-007, 5.894644e-007, 1.864508e-006, 3.20139e-006, 
    1.799564e-006, 1.095235e-006, 1.215314e-006, 1.611686e-006, 
    2.394119e-006, 1.757592e-006, 9.040041e-007, 1.292055e-006, 
    1.561765e-006, 1.949941e-006, 2.954776e-006, 3.731995e-006, 4.63687e-006, 
    3.870204e-006, 3.74727e-006, 3.863498e-006, 3.635759e-006, 4.100427e-006, 
    3.741805e-006, 2.803777e-006, 2.610932e-006, 2.095103e-006, 2.10156e-006, 
    3.185248e-006, 3.887093e-006, 2.261871e-006, 8.759398e-007, 
    3.226096e-007, -5.885977e-008, -1.394501e-007, 1.266351e-006, 
    4.122558e-008, -2.486013e-007, 7.797044e-007, 1.47149e-006, 
    2.177432e-006, 2.371271e-006, 2.637134e-006, 2.818184e-006, 
    1.154964e-006, 5.718321e-007, -1.933422e-007,
  -1.679486e-006, -2.702574e-006, -2.371147e-006, -1.543263e-006, 
    -1.632174e-006, -1.695504e-006, -5.669881e-007, 7.205945e-007, 
    1.112869e-006, 1.959379e-006, 2.115468e-006, 8.650122e-007, 4.65785e-007, 
    7.718791e-007, 1.250456e-006, 2.214809e-006, 2.40927e-006, 2.827372e-006, 
    2.649675e-006, 3.140171e-006, 3.944462e-006, 4.648169e-006, 
    4.753719e-006, 4.461656e-006, 3.180156e-006, 2.571195e-006, 3.26832e-006, 
    2.570202e-006, 2.012153e-006, 2.18538e-006, 1.736978e-006, 2.074863e-006, 
    3.217533e-006, 3.871198e-006, 3.775582e-006, 2.822156e-006, 
    1.983097e-006, 1.972914e-006, 1.807635e-006, 1.308943e-006, 
    8.296224e-007, 8.211778e-007, 1.689543e-006, 2.07449e-006, 1.826634e-006, 
    2.432118e-006, 3.515308e-006, 4.033869e-006, 3.562868e-006, 
    2.386918e-006, 1.479685e-006, 1.0781e-006, 1.114607e-006, 1.651173e-006, 
    2.405916e-006, 2.94124e-006, 2.289812e-006, 1.838059e-006, 1.920015e-006, 
    2.005199e-006, 2.227475e-006, 2.309059e-006, 2.234677e-006, 
    2.636761e-006, 3.138185e-006, 3.759811e-006, 3.948808e-006, 
    3.283347e-006, 2.368291e-006, 2.328555e-006, 2.505009e-006, 
    2.791608e-006, 3.272792e-006, 3.506119e-006, 3.724669e-006, 
    3.871198e-006, 4.530201e-006, 5.507221e-006, 3.61912e-006, 2.387414e-006, 
    1.578157e-006, 4.282842e-007, -6.712971e-007, -7.811932e-007, 
    -2.293536e-007, 3.539026e-007, 7.255626e-007, -4.729882e-007, 
    -2.422308e-006, -3.806254e-006, -3.139177e-006, -6.109476e-007, 
    1.596411e-006, 1.768394e-006, 4.04194e-007, -9.577725e-007,
  5.311031e-007, -3.563855e-008, -2.110937e-008, 4.701324e-007, 
    9.706864e-007, 8.530924e-007, 4.896274e-007, 1.064191e-007, 
    6.755181e-008, 2.719462e-007, 6.68193e-007, 7.804483e-007, 1.152232e-006, 
    1.627952e-006, 1.879161e-006, 1.821419e-006, 1.976018e-006, 
    2.274662e-006, 2.302726e-006, 2.519166e-006, 2.832587e-006, 2.71375e-006, 
    2.641976e-006, 2.73399e-006, 2.335509e-006, 2.184634e-006, 2.614781e-006, 
    3.053621e-006, 3.72678e-006, 4.065534e-006, 3.51059e-006, 2.33762e-006, 
    1.704444e-006, 1.469503e-006, 1.585484e-006, 2.252062e-006, 
    2.943104e-006, 3.388028e-006, 3.620734e-006, 3.488114e-006, 
    3.120304e-006, 3.031889e-006, 2.811352e-006, 2.404054e-006, 
    2.130617e-006, 2.216424e-006, 2.301857e-006, 2.318e-006, 2.553066e-006, 
    2.511342e-006, 2.462666e-006, 2.534191e-006, 2.893681e-006, 
    2.997369e-006, 2.286707e-006, 1.507625e-006, 1.650676e-006, 
    2.090633e-006, 2.160295e-006, 2.064184e-006, 2.008926e-006, 
    1.927961e-006, 1.753245e-006, 1.618142e-006, 1.404931e-006, 
    1.593555e-006, 1.951059e-006, 2.526865e-006, 2.687797e-006, 
    2.860154e-006, 3.188352e-006, 3.818919e-006, 4.156679e-006, 
    3.685057e-006, 2.949188e-006, 2.360344e-006, 1.87022e-006, 1.166636e-006, 
    6.377704e-007, 4.616877e-007, 5.080055e-007, 5.058941e-007, 
    1.370909e-007, -1.73226e-007, 5.28994e-008, -1.660237e-007, 
    -6.561477e-007, -1.129632e-006, -1.264736e-006, -1.654649e-006, 
    -2.076849e-006, -2.289935e-006, -1.14565e-006, 5.441398e-007, 
    1.290193e-006, 1.089151e-006,
  -8.061534e-007, -9.888163e-007, -7.373592e-007, -4.122658e-007, 
    -2.179295e-007, 4.96766e-009, 4.467865e-007, 8.124853e-007, 
    9.181595e-007, 8.653851e-007, 8.294983e-007, 8.481247e-007, 7.28046e-007, 
    5.551919e-007, 9.387732e-007, 1.243874e-006, 1.288701e-006, 
    1.302858e-006, 1.386925e-006, 1.567478e-006, 1.810366e-006, 
    2.053628e-006, 2.220149e-006, 2.170726e-006, 2.337868e-006, 
    2.998114e-006, 3.742923e-006, 4.0556e-006, 3.650412e-006, 2.626206e-006, 
    1.818439e-006, 1.41561e-006, 1.273552e-006, 1.440073e-006, 2.044191e-006, 
    2.736723e-006, 3.18264e-006, 3.393739e-006, 3.530209e-006, 3.475696e-006, 
    3.067901e-006, 2.580384e-006, 2.422184e-006, 2.567967e-006, 
    2.529223e-006, 2.378473e-006, 2.375494e-006, 2.762179e-006, 
    3.400196e-006, 3.656249e-006, 3.284961e-006, 2.772734e-006, 
    2.507121e-006, 2.308935e-006, 2.084921e-006, 2.236168e-006, 
    2.735481e-006, 2.943104e-006, 2.566353e-006, 2.144153e-006, 
    2.047792e-006, 2.088771e-006, 2.155949e-006, 2.205621e-006, 
    2.155204e-006, 2.059216e-006, 2.087652e-006, 1.925851e-006, 
    1.859541e-006, 1.961117e-006, 2.112984e-006, 2.348174e-006, 
    2.327685e-006, 2.250696e-006, 2.388036e-006, 2.73337e-006, 3.203377e-006, 
    3.513073e-006, 3.303339e-006, 2.984579e-006, 2.78689e-006, 2.228345e-006, 
    1.376246e-006, 7.071844e-007, 3.532814e-007, 4.408259e-007, 
    8.334714e-007, 1.060218e-006, 9.849668e-007, 1.040225e-006, 
    1.132737e-006, 8.78671e-007, 2.458692e-007, -9.077303e-008, 
    -9.623636e-008, -3.042323e-007,
  -5.487354e-007, -3.454579e-007, -1.585731e-007, -6.08452e-009, 
    5.43896e-008, 9.896848e-008, 2.235174e-007, 3.335372e-007, 3.520399e-007, 
    3.556415e-007, 2.970301e-007, 1.064191e-007, -1.100198e-007, 
    -2.471106e-007, -1.744675e-007, 5.12855e-008, 2.878414e-007, 
    4.25428e-007, 5.148349e-007, 5.889679e-007, 7.251901e-007, 9.108335e-007, 
    1.107654e-006, 1.346444e-006, 1.62435e-006, 1.923368e-006, 2.212947e-006, 
    2.412002e-006, 2.512087e-006, 2.430876e-006, 2.326692e-006, 
    2.269695e-006, 2.139311e-006, 1.947707e-006, 1.795093e-006, 
    1.733874e-006, 1.704693e-006, 1.54761e-006, 1.31006e-006, 1.138325e-006, 
    1.080334e-006, 1.113738e-006, 1.180296e-006, 1.193334e-006, 
    1.113614e-006, 9.847181e-007, 9.181599e-007, 9.864566e-007, 
    1.237542e-006, 1.523271e-006, 1.697863e-006, 1.707176e-006, 
    1.580641e-006, 1.435478e-006, 1.35377e-006, 1.467392e-006, 1.738842e-006, 
    2.003709e-006, 2.076104e-006, 1.912812e-006, 1.670544e-006, 
    1.554688e-006, 1.55146e-006, 1.561517e-006, 1.525879e-006, 1.462425e-006, 
    1.369417e-006, 1.207615e-006, 9.50818e-007, 6.829696e-007, 6.016344e-007, 
    8.357069e-007, 1.282742e-006, 1.669427e-006, 1.842777e-006, 
    1.805276e-006, 1.713385e-006, 1.716862e-006, 1.800557e-006, 
    1.852711e-006, 1.816079e-006, 1.745671e-006, 1.657754e-006, 
    1.454478e-006, 1.056492e-006, 5.94805e-007, 1.947087e-007, 
    -1.359731e-007, -5.003062e-007, -8.904685e-007, -1.25356e-006, 
    -1.45634e-006, -1.434733e-006, -1.206373e-006, -9.755295e-007, 
    -7.847939e-007,
  3.820905e-007, 4.456688e-007, 4.746016e-007, 4.659096e-007, 4.37597e-007, 
    4.069252e-007, 3.92025e-007, 3.967434e-007, 4.055601e-007, 4.033245e-007, 
    3.930181e-007, 3.843261e-007, 3.854439e-007, 4.044432e-007, 
    4.476551e-007, 5.145866e-007, 6.022556e-007, 6.955115e-007, 
    7.833041e-007, 8.421639e-007, 8.684892e-007, 8.750703e-007, 
    8.786719e-007, 8.997822e-007, 9.392697e-007, 9.855876e-007, 
    1.034513e-006, 1.078347e-006, 1.113117e-006, 1.146023e-006, 
    1.182407e-006, 1.225496e-006, 1.281624e-006, 1.359359e-006, 
    1.459568e-006, 1.565739e-006, 1.659244e-006, 1.722078e-006, 
    1.754488e-006, 1.761938e-006, 1.74207e-006, 1.694138e-006, 1.610816e-006, 
    1.494711e-006, 1.360972e-006, 1.212085e-006, 1.057237e-006, 
    9.037553e-007, 7.61946e-007, 6.402533e-007, 5.50101e-007, 5.072602e-007, 
    5.155803e-007, 5.559373e-007, 6.13431e-007, 6.744012e-007, 7.227063e-007, 
    7.564822e-007, 7.725007e-007, 7.711346e-007, 7.651752e-007, 
    7.722529e-007, 8.061534e-007, 8.697316e-007, 9.590144e-007, 
    1.070773e-006, 1.195446e-006, 1.319374e-006, 1.43672e-006, 1.528114e-006, 
    1.588588e-006, 1.61392e-006, 1.609946e-006, 1.571824e-006, 1.497939e-006, 
    1.375377e-006, 1.186381e-006, 9.362898e-007, 6.526711e-007, 
    3.635887e-007, 9.958967e-008, -1.210719e-007, -2.898278e-007, 
    -4.055601e-007, -4.79693e-007, -5.17939e-007, -5.255142e-007, 
    -5.102402e-007, -4.769618e-007, -4.235662e-007, -3.471969e-007, 
    -2.45248e-007, -1.177195e-007, 2.781599e-008, 1.696253e-007, 2.900761e-007,
  4.667525e-007, 4.59426e-007, 4.483743e-007, 4.370743e-007, 4.271403e-007, 
    4.226702e-007, 4.229183e-007, 4.246568e-007, 4.302448e-007, 
    4.414206e-007, 4.54956e-007, 4.697328e-007, 4.84013e-007, 4.951888e-007, 
    5.054954e-007, 5.13691e-007, 5.155538e-007, 5.059921e-007, 4.847584e-007, 
    4.565702e-007, 4.250295e-007, 3.943578e-007, 3.72627e-007, 3.540006e-007, 
    3.418313e-007, 3.309037e-007, 3.204729e-007, 3.110354e-007, 
    3.007287e-007, 2.890562e-007, 2.725408e-007, 2.545353e-007, 
    2.324317e-007, 2.123153e-007, 1.898393e-007, 1.684809e-007, 1.46005e-007, 
    1.338358e-007, 1.322214e-007, 1.412865e-007, 1.596646e-007, 
    1.847482e-007, 2.16289e-007, 2.515551e-007, 2.878146e-007, 3.191067e-007, 
    3.407135e-007, 3.475434e-007, 3.398445e-007, 3.193554e-007, 
    2.878146e-007, 2.504373e-007, 2.092111e-007, 1.730757e-007, 
    1.468745e-007, 1.334633e-007, 1.354499e-007, 1.50972e-007, 1.802778e-007, 
    2.229942e-007, 2.806121e-007, 3.537518e-007, 4.409237e-007, 
    5.362913e-007, 6.284301e-007, 7.098897e-007, 7.744613e-007, 
    8.082375e-007, 8.166817e-007, 7.98676e-007, 7.575736e-007, 6.966034e-007, 
    6.283062e-007, 5.595125e-007, 4.924573e-007, 4.318592e-007, 
    3.870314e-007, 3.587193e-007, 3.453083e-007, 3.471707e-007, 3.5785e-007, 
    3.769733e-007, 3.994489e-007, 4.195656e-007, 4.36205e-007, 4.52224e-007, 
    4.630272e-007, 4.717197e-007, 4.784251e-007, 4.820261e-007, 
    4.878625e-007, 4.914637e-007, 4.900976e-007, 4.856272e-007, 4.78301e-007, 
    4.722162e-007,
  1.006808e-007, 1.101182e-007, 1.271305e-007, 1.292414e-007, 1.414106e-007, 
    1.672394e-007, 2.000218e-007, 2.172824e-007, 2.182758e-007, 2.00767e-007, 
    1.735724e-007, 1.431491e-007, 1.155819e-007, 1.062687e-007, 
    1.165753e-007, 1.483645e-007, 1.900877e-007, 2.441045e-007, 
    2.965069e-007, 3.152574e-007, 2.972519e-007, 2.684429e-007, 
    2.674495e-007, 2.926574e-007, 3.166233e-007, 3.022188e-007, 
    2.617375e-007, 2.210076e-007, 1.934406e-007, 1.849965e-007, 
    1.904602e-007, 1.986559e-007, 2.17034e-007, 2.64966e-007, 3.378576e-007, 
    4.128601e-007, 4.787978e-007, 5.165474e-007, 5.442388e-007, 
    5.680805e-007, 5.864587e-007, 5.74786e-007, 5.242462e-007, 4.519754e-007, 
    3.88149e-007, 3.357466e-007, 3.090488e-007, 3.249431e-007, 3.751102e-007, 
    4.167093e-007, 4.237877e-007, 3.818154e-007, 2.526726e-007, 
    4.740923e-008, -2.059105e-007, -4.315398e-007, -5.884976e-007, 
    -6.918126e-007, -7.375093e-007, -6.705782e-007, -4.97228e-007, 
    -2.466404e-007, 7.672952e-009, 1.725784e-007, 3.100417e-007, 
    4.838889e-007, 6.612127e-007, 7.56208e-007, 6.988384e-007, 6.062028e-007, 
    5.850927e-007, 6.720161e-007, 7.631618e-007, 8.081138e-007, 
    8.024012e-007, 7.465219e-007, 6.295477e-007, 4.78673e-007, 3.204723e-007, 
    1.764279e-007, 9.310543e-008, 4.865069e-008, -4.609592e-008, 
    -1.795852e-007, -2.573192e-007, -2.173351e-007, -6.857135e-008, 
    1.306071e-007, 3.218393e-007, 4.671253e-007, 5.20645e-007, 4.820265e-007, 
    3.836788e-007, 2.69933e-007, 1.853691e-007, 1.250191e-007,
  1.664944e-007, 1.825131e-007, 2.421177e-007, 3.019707e-007, 3.603334e-007, 
    3.799533e-007, 3.455565e-007, 3.085519e-007, 3.059442e-007, 
    3.311522e-007, 3.569808e-007, 3.951029e-007, 4.422899e-007, 
    4.710989e-007, 4.646417e-007, 4.286305e-007, 3.718819e-007, 2.82475e-007, 
    2.231188e-007, 2.052374e-007, 1.635141e-007, 1.132227e-007, 
    1.077589e-007, 1.594161e-007, 2.62855e-007, 3.443147e-007, 4.148469e-007, 
    4.728372e-007, 4.871175e-007, 4.389371e-007, 3.729995e-007, 
    3.397203e-007, 3.31028e-007, 3.269301e-007, 3.484126e-007, 4.215524e-007, 
    5.299585e-007, 6.230907e-007, 5.965169e-007, 4.985419e-007, 
    5.082274e-007, 6.065751e-007, 7.112557e-007, 7.804218e-007, 
    8.086101e-007, 7.450319e-007, 6.18496e-007, 5.292131e-007, 6.666764e-007, 
    8.913112e-007, 9.095652e-007, 8.041393e-007, 7.629124e-007, 
    6.649375e-007, 5.232528e-007, 3.589671e-007, 2.437318e-007, 
    2.588813e-007, 3.107866e-007, 4.071476e-007, 6.129076e-007, 
    8.648617e-007, 7.840231e-007, 3.359946e-007, -5.652646e-008, 
    -1.230851e-007, 2.510583e-007, 8.052566e-007, 1.296746e-006, 
    1.631154e-006, 1.703921e-006, 1.620723e-006, 1.448242e-006, 1.11756e-006, 
    6.571145e-007, 4.290032e-007, 4.02305e-007, 4.014355e-007, 4.407993e-007, 
    5.562833e-007, 8.058778e-007, 9.820842e-007, 7.617955e-007, 
    3.871551e-007, 1.11856e-007, 2.801148e-007, 7.517365e-007, 1.101541e-006, 
    1.346666e-006, 1.454327e-006, 1.354116e-006, 1.036722e-006, 
    7.045503e-007, 4.116184e-007, 2.220011e-007, 1.679844e-007,
  9.360281e-008, 2.272164e-007, 2.643451e-007, 2.76266e-007, 3.42452e-007, 
    4.855033e-007, 6.351355e-007, 6.466839e-007, 5.958959e-007, 4.81902e-007, 
    3.72006e-007, 3.51517e-007, 3.838028e-007, 3.877764e-007, 4.434073e-007, 
    5.2139e-007, 5.036328e-007, 4.625306e-007, 3.797049e-007, 3.289168e-007, 
    3.453082e-007, 3.737446e-007, 3.603334e-007, 3.702676e-007, 
    4.568185e-007, 5.325661e-007, 5.500749e-007, 6.263191e-007, 
    7.165954e-007, 7.287647e-007, 6.50906e-007, 5.955234e-007, 5.739167e-007, 
    5.791321e-007, 6.408478e-007, 6.917603e-007, 7.286405e-007, 
    7.410582e-007, 7.00701e-007, 7.431692e-007, 9.362633e-007, 1.356973e-006, 
    1.853678e-006, 2.344424e-006, 2.598736e-006, 2.475553e-006, 
    2.479651e-006, 2.340325e-006, 1.958484e-006, 1.927315e-006, 
    2.047766e-006, 1.632892e-006, 1.214667e-006, 8.695802e-007, 
    5.664656e-007, 5.24743e-007, 7.047993e-007, 6.598457e-007, 6.142727e-007, 
    4.218e-007, 3.81815e-007, 1.194922e-006, 1.874415e-006, 2.103147e-006, 
    2.279727e-006, 2.696959e-006, 3.897871e-006, 5.52843e-006, 6.378789e-006, 
    6.067851e-006, 4.987516e-006, 4.038312e-006, 3.124624e-006, 
    2.135683e-006, 1.671387e-006, 1.84126e-006, 2.152819e-006, 2.173184e-006, 
    2.207953e-006, 1.995736e-006, 1.237639e-006, 4.661297e-007, 
    9.496671e-008, 5.581442e-007, 1.574156e-006, 2.125003e-006, 
    1.946064e-006, 1.379697e-006, 1.098437e-006, 1.046035e-006, 
    8.786451e-007, 6.88407e-007, 2.475804e-007, -1.002363e-007, 
    -7.627045e-008, 5.386642e-008,
  -2.523439e-008, 8.55548e-007, 1.215909e-006, 9.755031e-007, 8.689599e-007, 
    1.289794e-006, 1.493318e-006, 1.345921e-006, 1.010397e-006, 
    7.203209e-007, 7.23177e-007, 9.928879e-007, 1.363057e-006, 1.242482e-006, 
    1.008782e-006, 7.78311e-007, 4.995348e-007, 3.720062e-007, 4.994112e-007, 
    7.928395e-007, 1.138919e-006, 1.224228e-006, 1.051747e-006, 
    9.553867e-007, 9.912735e-007, 1.057087e-006, 1.085399e-006, 
    9.911494e-007, 9.78856e-007, 1.189459e-006, 1.443276e-006, 1.730744e-006, 
    1.597378e-006, 1.192191e-006, 8.3953e-007, 9.430935e-007, 1.180642e-006, 
    1.39435e-006, 1.630658e-006, 1.964443e-006, 2.224717e-006, 2.343181e-006, 
    2.380434e-006, 2.488964e-006, 2.590913e-006, 3.190809e-006, 
    3.611643e-006, 3.986032e-006, 3.614497e-006, 1.77495e-006, 5.669626e-007, 
    -9.710675e-009, 1.349526e-007, 8.549268e-007, 1.353868e-006, 
    2.31462e-006, 3.126361e-006, 2.927803e-006, 2.642198e-006, 2.2611e-006, 
    1.710132e-006, 2.713601e-006, 3.875146e-006, 4.845088e-006, 
    5.093689e-006, 4.082021e-006, 3.799521e-006, 4.89041e-006, 4.994222e-006, 
    4.613374e-006, 5.409717e-006, 5.83887e-006, 5.552021e-006, 4.164599e-006, 
    2.624315e-006, 2.312509e-006, 3.189815e-006, 3.077809e-006, 
    1.869324e-006, 8.930501e-007, 1.311046e-007, -7.167637e-008, 
    -1.132503e-008, 1.91827e-007, 1.018219e-006, 1.888447e-006, 
    1.647048e-006, 7.382023e-007, 4.355843e-007, 4.121148e-007, 3.09049e-007, 
    4.612884e-007, 3.1327e-007, -8.235656e-008, -7.387525e-007, -6.756682e-007,
  2.440411e-006, 2.958598e-006, 2.972877e-006, 2.5893e-006, 2.081543e-006, 
    1.963821e-006, 2.113702e-006, 1.893289e-006, 2.067634e-006, 
    2.845971e-006, 2.814555e-006, 3.091094e-006, 3.885078e-006, 
    4.064886e-006, 4.200114e-006, 3.935992e-006, 3.065391e-006, 
    1.980462e-006, 1.699699e-006, 2.215528e-006, 2.734834e-006, 
    2.990761e-006, 3.115931e-006, 2.913772e-006, 2.934134e-006, 
    2.571294e-006, 2.539753e-006, 2.789099e-006, 2.717944e-006, 
    3.515901e-006, 4.406618e-006, 4.529056e-006, 4.195269e-006, 
    2.797915e-006, 2.400922e-006, 3.203971e-006, 4.140757e-006, 4.61747e-006, 
    4.81603e-006, 4.433442e-006, 3.435065e-006, 1.715098e-006, 2.266317e-006, 
    3.842862e-006, 4.788091e-006, 4.938844e-006, 4.44698e-006, 4.3608e-006, 
    3.803994e-006, 3.154302e-006, 2.320457e-006, 2.148596e-006, 
    2.131212e-006, 1.372369e-006, 8.156858e-007, 2.142263e-006, 
    2.917123e-006, 3.046266e-006, 2.772581e-006, 2.209074e-006, 
    3.184353e-006, 3.033724e-006, 2.438174e-006, 2.600721e-006, 
    3.659698e-006, 3.472191e-006, 2.203357e-006, 3.029256e-006, 
    4.354341e-006, 4.981433e-006, 5.652481e-006, 5.710223e-006, 
    6.084865e-006, 6.023273e-006, 5.193154e-006, 4.432075e-006, 
    3.617231e-006, 2.387884e-006, 1.369389e-006, 1.214168e-006, 
    2.010387e-006, 2.551548e-006, 3.050117e-006, 3.36776e-006, 2.717821e-006, 
    2.13146e-006, 8.185434e-007, 3.099176e-007, 8.195366e-007, 1.581731e-006, 
    2.203483e-006, 2.541491e-006, 2.620219e-006, 2.606806e-006, 
    1.742291e-006, 1.357593e-006,
  3.370369e-006, 2.860004e-006, 2.644063e-006, 2.792824e-006, 3.385519e-006, 
    4.268164e-006, 3.253766e-006, 3.562097e-006, 5.842223e-006, 
    6.274606e-006, 5.887051e-006, 4.719172e-006, 5.087357e-006, 
    6.086726e-006, 7.161099e-006, 7.449813e-006, 6.180479e-006, 
    5.911142e-006, 6.135279e-006, 6.559218e-006, 6.439634e-006, 
    5.482731e-006, 4.811558e-006, 5.231522e-006, 5.320929e-006, 4.23749e-006, 
    2.964186e-006, 3.2976e-006, 4.262822e-006, 5.3069e-006, 5.326148e-006, 
    5.461625e-006, 6.197492e-006, 6.615097e-006, 6.383134e-006, 
    7.484829e-006, 9.237825e-006, 7.539093e-006, 5.747104e-006, 
    5.004902e-006, 6.236112e-006, 5.984528e-006, 5.299325e-006, 
    3.316227e-006, 4.118159e-006, 6.209413e-006, 6.508057e-006, 
    7.549648e-006, 6.19029e-006, 3.553654e-006, 3.45357e-006, 3.968527e-006, 
    3.591156e-006, 3.513049e-006, 3.413457e-006, 2.725397e-006, 
    2.360568e-006, 3.948659e-006, 5.631869e-006, 5.853648e-006, 
    6.339425e-006, 5.617216e-006, 5.451813e-006, 5.02154e-006, 4.425867e-006, 
    4.263941e-006, 4.313861e-006, 4.615114e-006, 4.755557e-006, 
    4.495779e-006, 3.651005e-006, 3.44624e-006, 3.649145e-006, 2.982939e-006, 
    2.282584e-006, 2.600103e-006, 3.755687e-006, 4.782751e-006, 
    4.757419e-006, 4.008632e-006, 4.551036e-006, 4.383895e-006, 
    3.818272e-006, 3.980196e-006, 3.714958e-006, 3.446984e-006, 
    3.350003e-006, 2.826599e-006, 2.396079e-006, 1.460783e-006, 1.79072e-006, 
    2.85491e-006, 3.538627e-006, 2.8641e-006, 2.273767e-006, 2.795804e-006,
  3.840997e-006, 3.089855e-006, 3.56843e-006, 3.047635e-006, 2.478908e-006, 
    3.125244e-006, 2.799159e-006, 2.542858e-006, 2.973997e-006, 
    4.370486e-006, 4.360179e-006, 4.403144e-006, 5.681166e-006, 5.89537e-006, 
    6.132797e-006, 7.053564e-006, 6.959437e-006, 5.869293e-006, 
    6.408717e-006, 7.405107e-006, 7.033944e-006, 6.740142e-006, 
    5.725622e-006, 5.189429e-006, 4.846577e-006, 4.590775e-006, 
    5.534017e-006, 5.733818e-006, 4.329631e-006, 3.866329e-006, 
    3.927424e-006, 4.471689e-006, 2.929666e-006, 4.550044e-006, 
    6.320799e-006, 5.975835e-006, 5.400156e-006, 5.921074e-006, 
    5.309259e-006, 4.184221e-006, 5.412325e-006, 5.392456e-006, 
    5.190297e-006, 6.610006e-006, 8.025243e-006, 8.061752e-006, 
    6.850411e-006, 7.602299e-006, 6.134658e-006, 5.396801e-006, 
    4.427109e-006, 3.798654e-006, 4.516267e-006, 7.167184e-006, 7.69183e-006, 
    4.633615e-006, 4.138026e-006, 4.898111e-006, 3.108358e-006, 
    2.110228e-006, 3.934505e-006, 4.225449e-006, 3.485979e-006, 
    5.132555e-006, 5.607533e-006, 5.103127e-006, 5.022164e-006, 
    5.012229e-006, 4.473055e-006, 4.398549e-006, 4.140016e-006, 
    4.741772e-006, 5.535134e-006, 4.206697e-006, 3.620833e-006, 
    3.962195e-006, 5.570027e-006, 7.028604e-006, 5.1184e-006, 3.716948e-006, 
    2.890925e-006, 2.083778e-006, 1.476057e-006, 2.030629e-006, 
    2.266566e-006, 1.646553e-006, 2.847712e-006, 3.777292e-006, 
    2.232538e-006, 1.73124e-006, 1.914028e-006, 2.15617e-006, 3.091096e-006, 
    1.998842e-006, 1.53256e-006, 3.613257e-006,
  4.992238e-006, 4.430092e-006, 5.33248e-006, 4.764372e-006, 4.494414e-006, 
    5.209173e-006, 5.097412e-006, 6.685628e-006, 8.848036e-006, 
    7.024009e-006, 4.666645e-006, 5.73034e-006, 5.305285e-006, 5.183965e-006, 
    5.725373e-006, 8.069575e-006, 9.219695e-006, 7.861951e-006, 
    8.246525e-006, 8.83686e-006, 8.160596e-006, 7.523819e-006, 7.622664e-006, 
    7.285898e-006, 5.834276e-006, 6.98328e-006, 6.92293e-006, 6.367985e-006, 
    5.059539e-006, 5.092073e-006, 6.969371e-006, 5.984903e-006, 
    4.062653e-006, 3.131207e-006, 4.127845e-006, 5.891276e-006, 
    7.191278e-006, 8.484078e-006, 9.507663e-006, 9.244781e-006, 
    7.764475e-006, 7.152781e-006, 6.604294e-006, 7.726101e-006, 
    7.105597e-006, 7.054186e-006, 7.311475e-006, 5.598467e-006, 6.22717e-006, 
    7.282048e-006, 6.495142e-006, 5.949016e-006, 5.557611e-006, 
    4.607042e-006, 2.978097e-006, 1.452838e-006, 2.235645e-006, 
    3.218005e-006, 2.064407e-006, 2.337098e-006, 3.7465e-006, 4.823976e-006, 
    3.563711e-006, 3.231044e-006, 3.148218e-006, 3.219991e-006, 
    2.792949e-006, 4.871536e-006, 6.059532e-006, 5.543703e-006, 5.3521e-006, 
    4.707375e-006, 4.807958e-006, 5.899095e-006, 5.656952e-006, 
    5.578846e-006, 5.357313e-006, 4.396437e-006, 2.546334e-006, 
    7.350991e-007, 5.331894e-007, 5.437414e-007, 5.781403e-007, 
    1.018634e-010, 3.787136e-007, 5.797538e-007, 2.056708e-006, 
    2.796301e-006, 3.313744e-006, 2.919856e-006, 2.082039e-006, 2.5708e-006, 
    2.924702e-006, 2.652259e-006, 1.983943e-006, 3.370991e-006,
  4.826214e-006, 3.330013e-006, 2.714221e-006, 2.307666e-006, 4.153424e-006, 
    6.155271e-006, 8.206047e-006, 7.582803e-006, 5.909278e-006, 
    4.141877e-006, 5.332728e-006, 6.051709e-006, 6.925909e-006, 
    8.931482e-006, 1.007502e-005, 7.617078e-006, 6.663648e-006, 
    5.673715e-006, 5.363772e-006, 6.434544e-006, 7.473032e-006, 
    8.604031e-006, 8.807558e-006, 7.040033e-006, 6.566173e-006, 
    7.022643e-006, 7.928509e-006, 7.171529e-006, 6.104729e-006, 
    6.353952e-006, 7.375424e-006, 6.724989e-006, 5.0948e-006, 4.653601e-006, 
    5.887541e-006, 6.84879e-006, 7.693809e-006, 8.487303e-006, 6.920322e-006, 
    4.820005e-006, 4.443877e-006, 5.179496e-006, 5.049111e-006, 
    5.140129e-006, 5.385005e-006, 6.165581e-006, 6.036435e-006, 
    6.957576e-006, 4.329508e-006, 2.138291e-006, -5.714846e-007, 
    3.707664e-007, 2.229563e-006, 3.172556e-006, 3.036834e-006, 
    1.792585e-006, 1.438433e-006, 1.473079e-006, 2.112585e-006, 
    2.981324e-006, 4.722649e-006, 5.240465e-006, 2.635246e-006, 
    2.581601e-006, 3.509942e-006, 4.507081e-006, 4.909161e-006, 
    5.194644e-006, 4.020432e-006, 3.203475e-006, 4.700794e-006, 
    4.257981e-006, 4.684651e-006, 4.066254e-006, 1.01375e-006, 
    -1.504668e-008, 8.517054e-007, 7.981798e-007, 1.63575e-006, 
    1.389011e-006, -4.999565e-007, -8.101506e-007, 5.254878e-007, 
    2.200009e-006, 2.209195e-006, 4.511076e-007, 6.28308e-007, 2.198145e-006, 
    2.96096e-006, 3.580475e-006, 5.756418e-006, 5.795036e-006, 5.465472e-006, 
    6.136894e-006, 6.458387e-006, 5.870039e-006,
  3.344916e-006, 4.378309e-006, 7.284534e-006, 7.644019e-006, 7.18469e-006, 
    6.839733e-006, 4.441639e-006, 1.336237e-006, 2.542236e-006, 
    4.990623e-006, 6.489308e-006, 6.163842e-006, 5.716807e-006, 
    4.692973e-006, 3.779654e-006, 4.996207e-006, 7.655071e-006, 
    1.073812e-005, 1.042756e-005, 9.498217e-006, 7.918818e-006, 
    6.943414e-006, 7.63818e-006, 8.828159e-006, 8.49189e-006, 7.662395e-006, 
    7.548773e-006, 6.803341e-006, 6.444225e-006, 5.794907e-006, 
    4.569039e-006, 2.270783e-006, 1.042677e-006, 2.519009e-006, 3.2149e-006, 
    3.243829e-006, 2.418306e-006, 2.129975e-006, 1.63774e-006, 8.910647e-007, 
    1.130602e-006, 3.318341e-006, 6.683395e-006, 5.078913e-006, 
    1.882236e-006, 1.892549e-006, 1.909682e-006, 1.620352e-006, 
    -1.455372e-006, -2.050301e-006, -2.430652e-006, -2.383465e-006, 
    4.005669e-007, -1.022991e-006, -2.875327e-006, -2.254819e-006, 
    9.781124e-007, 2.213666e-006, 2.916504e-006, 4.499505e-006, 
    5.328009e-006, 2.818157e-006, 2.927682e-006, 3.319828e-006, 
    9.079522e-007, 1.379325e-006, 3.61065e-006, 5.119768e-006, 5.169812e-006, 
    2.411729e-006, 2.013123e-006, 2.082536e-006, -2.207882e-006, 
    -1.957666e-006, -4.119156e-007, -9.766736e-007, 1.325679e-006, 
    1.805274e-007, -1.372298e-006, -7.598619e-007, -5.591928e-007, 
    -2.002247e-006, -3.267323e-007, -6.710725e-007, -2.079109e-006, 
    2.587603e-007, 1.974502e-006, 3.187333e-006, 3.61922e-006, 5.070719e-006, 
    6.339926e-006, 6.962917e-006, 5.621316e-006, 5.24059e-006, 5.26791e-006, 
    3.78338e-006,
  3.741905e-006, 4.230911e-006, 4.722773e-006, 3.965171e-006, 3.373472e-006, 
    1.213799e-006, 7.361086e-008, 1.280978e-006, 2.16027e-006, 2.40378e-006, 
    4.677699e-006, 5.361535e-006, 5.622307e-006, 6.641047e-006, 
    6.694074e-006, 8.072548e-006, 8.590116e-006, 8.36399e-006, 7.386847e-006, 
    6.950737e-006, 8.256702e-006, 1.007452e-005, 9.694912e-006, 
    5.952363e-006, 3.873527e-006, 3.40426e-006, 1.221742e-006, 4.456379e-007, 
    1.50449e-006, 3.660389e-007, -1.917313e-006, -1.973436e-006, 
    -9.864816e-007, -4.994617e-007, -7.167691e-007, -1.222044e-006, 
    -1.437242e-006, -2.965357e-006, -3.180305e-006, -2.134369e-006, 
    -1.548504e-006, -7.125491e-007, 1.197532e-006, 1.401182e-006, 
    2.318473e-006, 8.189163e-007, 3.207224e-007, 1.30929e-006, 
    -6.945429e-007, -3.308331e-006, -7.229573e-008, -2.638524e-006, 
    -1.846154e-006, -4.545109e-007, -2.050798e-006, -1.610344e-006, 
    -2.147262e-007, 5.811198e-007, 1.179898e-006, 9.638316e-007, 
    1.804505e-006, 7.841481e-007, 1.853679e-006, 2.520506e-006, 
    1.815681e-006, 2.567693e-006, 2.349392e-006, 2.926439e-006, 3.76314e-006, 
    -1.939879e-007, -2.383094e-006, -5.371647e-006, -4.099955e-006, 
    -1.850625e-006, -3.318512e-006, -4.439949e-006, -6.832335e-006, 
    -5.876052e-006, -3.477335e-006, -2.84143e-006, -1.847523e-006, 
    -2.947228e-006, -2.684099e-006, -9.627638e-007, 8.302177e-007, 
    1.920362e-006, 2.321454e-006, 3.230176e-006, 3.751096e-006, 3.12562e-006, 
    4.056688e-006, 3.971752e-006, 2.458168e-006, 2.78699e-006, 3.590907e-006, 
    2.446992e-006,
  6.106711e-006, 6.05009e-006, 3.480141e-006, 8.113439e-007, -1.009794e-007, 
    -1.477947e-007, 3.265577e-007, 3.598605e-006, 3.889549e-006, 
    4.09643e-006, 7.009106e-006, 1.093519e-005, 1.046332e-005, 6.357797e-006, 
    5.494152e-006, 5.3105e-006, 5.342783e-006, 3.525958e-006, 2.287918e-006, 
    2.798159e-006, 2.123514e-006, 9.058385e-007, -2.028075e-006, 
    -3.625108e-006, -4.08692e-006, -5.541271e-006, -4.892943e-006, 
    -4.089274e-006, -6.394483e-006, -6.447759e-006, -4.29901e-006, 
    -3.23606e-006, -1.450777e-006, -6.483497e-007, -2.469893e-006, 
    -4.461555e-006, -3.931449e-006, -4.054133e-006, -3.800318e-006, 
    -4.593556e-006, -2.886753e-006, -8.882562e-007, -5.952024e-007, 
    1.063794e-006, -2.020606e-007, -1.476605e-006, -4.696594e-007, 
    2.879406e-007, -1.647844e-006, -4.288082e-006, -5.047796e-006, 
    -4.801923e-006, -4.689298e-006, -3.631189e-006, -4.271194e-006, 
    -1.221917e-006, -2.536575e-006, -1.961762e-006, -1.426564e-006, 
    1.103655e-006, 2.093338e-006, 4.333506e-007, 1.990149e-006, 
    6.865448e-007, -1.04323e-006, 4.662579e-007, -7.387498e-007, 
    2.684543e-006, -5.713591e-007, -3.548361e-006, -3.060228e-006, 
    -2.201547e-006, -3.489877e-006, -4.158443e-006, -4.849237e-006, 
    -7.119801e-006, -1.117093e-005, -8.158409e-006, -3.194338e-006, 
    -8.019579e-007, -3.219174e-006, -2.851239e-006, -2.903391e-006, 
    -3.321866e-006, -3.299265e-006, -1.425567e-006, 3.004174e-006, 
    5.450693e-006, 6.161721e-006, 7.54865e-006, 6.748083e-006, 4.224694e-006, 
    4.479007e-006, 4.587546e-006, 4.175152e-006, 6.040649e-006,
  -9.818868e-007, -4.954891e-007, -1.201553e-006, -2.351551e-006, 
    -1.71875e-006, -5.847724e-007, 1.175053e-006, 5.824841e-007, 
    1.708393e-006, 1.610419e-006, 1.595025e-006, 6.434529e-007, 
    -4.927719e-006, -4.087044e-006, -2.721725e-006, -3.428908e-006, 
    -5.438575e-006, -8.003561e-006, -6.914906e-006, -6.44875e-006, 
    -9.501253e-006, -9.91116e-006, -1.000665e-005, -1.012983e-005, 
    -1.029921e-005, -8.663934e-006, -8.040444e-006, -9.100663e-006, 
    -7.006181e-006, -5.213198e-006, -3.460449e-006, -3.495218e-006, 
    -3.937908e-006, -4.116472e-006, -3.923006e-006, -3.521171e-006, 
    -2.85658e-006, -1.767181e-006, -1.660885e-006, 2.009256e-008, 
    -7.817143e-007, 6.076953e-007, -6.683149e-008, 9.835767e-007, 
    -4.208578e-007, -8.236875e-007, -2.985349e-006, -5.905727e-006, 
    -4.027312e-006, -6.035989e-006, -1.086893e-005, -1.029585e-005, 
    -5.657745e-006, -3.723948e-006, -2.029934e-006, -2.309953e-006, 
    -2.133873e-006, -3.09723e-007, -9.626383e-007, -2.373235e-007, 
    -5.355003e-006, -3.855825e-006, -2.251963e-006, -2.620025e-006, 
    -9.548203e-007, -1.684981e-006, -1.874105e-007, -1.386332e-006, 
    -9.180658e-007, -3.511941e-007, -3.146888e-007, -2.611951e-006, 
    -2.41451e-006, -1.21745e-006, -2.941888e-006, -6.86499e-006, 
    -8.24223e-006, -1.017317e-005, -3.278032e-006, -1.525159e-006, 
    -4.257537e-006, -3.996269e-006, -2.353167e-006, 8.30958e-007, 
    3.983172e-006, 7.818235e-006, 1.252352e-005, 1.063927e-005, 
    9.045347e-006, 9.193365e-006, 4.22656e-006, 9.130381e-007, 2.580971e-006, 
    4.02068e-006, 5.699167e-006, 2.184359e-006,
  -1.14133e-006, -1.299159e-007, -6.479786e-007, -1.041616e-006, 
    -1.012187e-006, -1.210965e-007, 4.16584e-007, 1.876033e-007, 
    -1.302265e-006, -3.823663e-006, -5.76429e-006, -2.172987e-006, 
    -8.665284e-007, -3.334904e-006, -4.164154e-006, -6.529963e-006, 
    -7.268438e-006, -8.356348e-006, -8.979094e-006, -8.59092e-006, 
    -8.071365e-006, -6.314395e-006, -6.091622e-006, -6.088268e-006, 
    -4.204388e-006, -4.295036e-006, -4.216805e-006, -3.489008e-006, 
    -2.037387e-006, -1.404585e-006, -3.125544e-006, -3.915926e-006, 
    -3.295541e-006, -1.396512e-006, -8.261713e-007, -3.839805e-007, 
    1.857029e-006, 2.415699e-006, 2.139158e-006, 3.692109e-006, 5.1898e-006, 
    3.92432e-006, 1.954882e-006, -3.67585e-007, -2.780562e-007, 
    -3.765797e-006, -3.517443e-006, -4.969437e-006, -5.415975e-006, 
    -1.057674e-005, -6.866354e-006, -4.026937e-006, -3.122041e-007, 
    -1.981382e-006, -2.353414e-006, -2.638397e-006, -9.245159e-007, 
    1.566877e-007, -2.113506e-006, -6.017362e-006, -7.796807e-006, 
    -4.231457e-006, -5.534443e-006, -1.555956e-006, 1.248955e-007, 
    8.937932e-007, -3.647365e-007, -8.12397e-008, 2.410015e-007, 
    -2.862507e-007, 9.479409e-007, 3.192921e-006, 2.886578e-006, 
    -1.15884e-006, -2.036644e-006, -2.039126e-006, -2.572589e-006, 
    -1.357895e-006, -2.883553e-008, 2.385186e-007, -1.977036e-006, 
    3.963063e-006, 7.022642e-006, 1.060388e-005, 1.249708e-005, 
    1.184329e-005, 8.834988e-006, 6.800856e-006, 5.125847e-006, 
    8.171392e-006, 6.044873e-006, 3.10388e-006, 2.401543e-006, 1.452609e-007, 
    -3.638765e-006, -4.44467e-006,
  -8.672732e-007, -1.287238e-006, -1.459595e-006, -1.496228e-006, 
    -9.389237e-007, -4.168865e-007, -1.194478e-006, -3.97069e-006, 
    -1.422963e-006, 2.229439e-006, 2.404153e-006, 2.306952e-007, 
    -2.844037e-006, -5.293665e-006, -5.978125e-006, -6.29229e-006, 
    -5.248713e-006, -4.611439e-006, -4.569469e-006, -1.750789e-006, 
    1.125259e-006, -1.16604e-006, -1.528512e-006, -8.754687e-007, 
    -1.044597e-006, -1.127051e-006, -9.176897e-007, -1.349451e-006, 
    -1.61047e-006, -1.823928e-006, -2.723338e-006, -3.990046e-007, 
    6.771074e-007, 8.110937e-007, 4.503604e-007, 9.913974e-007, 
    1.430858e-006, 1.135814e-006, 2.427497e-006, 1.178159e-006, 
    -7.614763e-007, -4.107778e-006, -5.508489e-006, -4.409652e-006, 
    -2.989449e-006, -2.812865e-006, -3.063828e-006, -4.371777e-006, 
    -5.486261e-006, -4.9261e-006, 1.951401e-006, 6.359045e-006, 
    7.620551e-006, 3.302448e-006, 9.692994e-007, -6.689661e-007, 
    -4.615868e-007, -2.788282e-006, -8.821138e-006, -9.134808e-006, 
    -6.875049e-006, -4.082201e-006, -2.039753e-006, 1.909801e-006, 
    5.065245e-006, 5.843958e-006, 3.273635e-006, 2.321696e-006, 
    1.491459e-006, 4.908792e-006, 4.272759e-006, 2.229188e-006, 
    1.258886e-007, -1.348707e-006, -4.081944e-007, 4.393178e-008, 
    2.144266e-007, 1.83232e-006, 1.775447e-006, 1.38094e-006, 3.535399e-006, 
    3.612884e-006, 1.118926e-005, 1.17627e-005, 1.077785e-005, 9.518455e-006, 
    4.423007e-006, 4.107973e-006, 6.704377e-006, 6.808295e-007, 
    -4.916168e-006, -3.977766e-006, -4.502659e-006, -4.117839e-006, 
    -4.084683e-006, -2.598542e-006,
  -9.584201e-007, -2.542151e-007, -3.706923e-007, -5.486377e-007, 
    1.407896e-007, 1.703434e-007, -1.630463e-006, -3.668691e-006, 
    4.158141e-006, 4.940453e-006, 1.338358e-007, -1.798721e-006, 
    -4.182657e-006, -8.711121e-006, -8.95786e-006, -3.947221e-006, 
    -3.152119e-006, -1.663741e-006, -8.682673e-007, 2.633256e-006, 
    2.685907e-006, 2.1065e-006, 1.310033e-006, 1.254029e-006, 6.199862e-007, 
    -5.354559e-008, -4.470603e-007, -8.307643e-007, -5.690026e-007, 
    -1.090295e-006, -5.014504e-007, -3.346813e-007, -8.8143e-007, 
    3.142641e-007, 5.187821e-007, 1.245213e-006, -7.87677e-007, 
    -5.752113e-007, -9.989012e-007, -1.544036e-006, -2.838821e-006, 
    -4.067299e-006, -4.800312e-006, -4.505268e-006, -2.622134e-006, 
    -3.278159e-006, -7.367407e-006, -5.834203e-006, -3.429774e-006, 
    1.003442e-006, 6.618946e-006, 1.242468e-005, 9.83871e-006, 2.992496e-006, 
    4.810317e-007, -1.188269e-006, -2.468776e-006, -3.881036e-006, 
    -2.007215e-006, 1.612527e-006, 2.937606e-006, 6.830411e-006, 
    6.057537e-006, 8.013812e-006, 5.348618e-006, 3.474179e-006, 
    6.774542e-006, 4.627407e-006, 3.114566e-006, 8.015313e-007, 
    5.022666e-007, -9.714586e-007, -1.297918e-006, -2.791749e-007, 
    -4.172593e-007, -1.101712e-007, 1.079315e-006, 2.196156e-006, 
    1.880003e-006, 4.322319e-007, 1.365661e-006, 6.583177e-006, 
    1.141066e-005, 4.196758e-006, 1.124263e-006, 1.167351e-006, 
    2.894267e-007, 3.086789e-007, -4.512221e-006, -4.9677e-006, 
    -4.841289e-006, -2.889238e-006, -1.674048e-006, -2.719363e-006, 
    -2.269596e-006, -2.134246e-006,
  4.492495e-008, -5.940856e-007, -9.694711e-007, -2.328569e-007, 
    8.863572e-008, 3.728765e-007, -1.311948e-006, 1.327046e-006, 
    1.79507e-006, -1.91557e-006, 1.733973e-006, -4.517797e-007, 
    -3.65491e-006, -1.145703e-005, -9.835414e-006, -1.456244e-006, 
    2.690631e-007, -1.173739e-007, 1.470842e-006, 3.170443e-006, 
    2.001447e-006, 1.776812e-006, 1.989047e-007, 2.568931e-007, 
    4.706008e-007, 2.940214e-008, -5.739685e-007, -9.230293e-007, 
    -8.223219e-007, -8.101529e-007, -6.134572e-007, -6.364301e-007, 
    -4.47061e-007, 1.25726e-006, 7.423e-007, 5.082279e-007, 8.331967e-007, 
    1.265454e-006, 1.933158e-007, -9.121018e-007, 7.95199e-007, 
    -1.720364e-006, -5.631795e-006, -7.639483e-008, -5.870079e-007, 
    -8.924084e-006, -8.667908e-006, -1.528861e-007, 5.578844e-006, 
    1.044916e-005, 9.8212e-006, 1.224971e-005, 8.6789e-006, 1.224224e-006, 
    -3.590711e-006, -1.048113e-005, -9.566946e-006, -3.827885e-006, 
    1.133452e-006, 4.39271e-006, 5.058795e-006, 8.537711e-006, 5.738162e-006, 
    3.390613e-006, 6.093087e-007, 2.695966e-006, 1.147114e-006, 
    -5.686306e-007, -2.76319e-007, -6.27364e-007, -1.171505e-006, 
    -1.080485e-006, -2.329812e-007, -4.547474e-008, -2.44157e-007, 
    3.722544e-007, 4.735823e-007, 1.007789e-006, 1.440667e-006, 
    2.996716e-006, 6.683138e-006, 9.113766e-006, 7.877097e-006, 
    -2.474189e-008, -3.660254e-006, -5.735234e-006, -4.949568e-006, 
    -6.10168e-006, -6.131731e-006, -5.566232e-006, -5.231202e-006, 
    -3.714761e-006, -2.838325e-006, -2.59258e-006, -3.510713e-007, 
    -9.908294e-007,
  -7.190079e-007, -2.740833e-007, -1.775988e-007, 1.907084e-007, 
    1.734481e-007, -1.456739e-006, -7.195058e-007, 2.654615e-007, 
    -6.189221e-007, -2.521675e-006, -5.430493e-007, 9.552641e-007, 
    -2.880915e-006, -2.043014e-005, -5.076356e-006, 2.926572e-007, 
    -2.750781e-006, -2.197327e-006, 7.478866e-007, 2.719559e-006, 
    1.789105e-006, -1.120316e-008, -6.507107e-007, 1.224107e-007, 
    -6.658593e-008, -3.554187e-007, -1.741723e-006, -2.243894e-006, 
    -1.38807e-006, -9.54073e-007, -9.142002e-008, 1.851206e-007, 
    1.34705e-007, 2.055588e-006, 2.081293e-006, 2.030133e-006, 1.46364e-006, 
    7.210658e-007, -6.125881e-007, 1.129978e-006, 2.009643e-006, 
    -3.515333e-006, -3.327456e-006, -4.227982e-006, -5.168989e-006, 
    -5.237162e-006, 3.240979e-006, 8.220813e-006, 1.199963e-005, 
    4.559104e-006, 2.906814e-006, -2.957164e-006, -7.50152e-006, 
    -7.232673e-006, -9.699066e-006, -9.798159e-006, -6.148242e-006, 
    5.254915e-007, 6.226055e-006, 7.422494e-006, 6.557109e-006, 
    1.225098e-006, -2.108663e-006, -1.605129e-006, -1.083342e-006, 
    -1.228752e-006, -1.72521e-006, -1.550245e-006, -1.007843e-006, 
    -1.879561e-006, -1.735266e-006, -1.415513e-006, -8.938478e-007, 
    -5.839036e-007, 2.890692e-008, 5.06489e-007, 6.523965e-007, 
    5.632374e-007, 5.703019e-006, -2.198212e-007, 4.050355e-006, 
    5.382888e-006, 3.608044e-006, -2.658517e-006, -8.450847e-006, 
    -9.387137e-006, -5.615158e-006, -3.335032e-006, -2.434999e-006, 
    -3.59158e-006, -2.350934e-006, -9.791574e-007, -1.52193e-006, 
    -3.069908e-007, -6.802647e-007, -6.230193e-007,
  -3.668433e-007, -3.127022e-007, -5.230413e-008, 1.448118e-006, 
    -9.514652e-007, -1.815484e-006, 3.313246e-006, 1.710006e-006, 
    1.568072e-006, -1.661009e-006, -7.42104e-007, -5.019319e-008, 
    6.103037e-007, -3.235192e-006, -2.78816e-006, -2.472751e-006, 
    -2.516337e-006, -3.03204e-006, -4.076983e-007, 5.808697e-007, 
    2.357585e-006, -1.669196e-007, -1.093897e-006, -1.5079e-006, 
    -7.229819e-007, -1.945124e-006, -1.852861e-006, -2.649329e-006, 
    -1.540061e-006, -4.948689e-007, -8.136169e-008, 2.816058e-007, 
    2.523e-007, 7.467704e-007, 2.175543e-006, 5.506959e-007, -3.783916e-007, 
    -5.214425e-007, 3.697824e-008, 4.87762e-008, 4.635231e-007, 
    -1.023736e-006, -7.658479e-006, -7.946814e-006, -1.391174e-006, 
    4.56184e-006, 7.174458e-008, 5.865812e-006, -8.870229e-007, 
    -7.992643e-006, -9.414707e-006, -9.900985e-006, -8.114584e-006, 
    -7.967679e-006, -3.954548e-006, 2.115317e-006, 3.213536e-006, 
    2.942335e-006, 6.310989e-006, 4.032725e-006, 2.084773e-006, 
    4.347148e-007, -1.594948e-006, -1.983247e-006, -1.430911e-006, 
    -2.327464e-006, -1.631828e-006, -2.129031e-006, -2.305362e-006, 
    -2.624121e-006, -1.896943e-006, -1.838953e-006, -1.24713e-006, 
    -8.584575e-007, -2.472616e-007, 4.641449e-007, 3.117806e-007, 
    2.731853e-006, -1.041371e-006, -3.193101e-006, 3.025278e-006, 
    3.435925e-006, 1.713608e-006, -3.029556e-006, -5.435722e-006, 
    -5.942609e-006, -1.137482e-006, -1.26675e-006, -3.348059e-007, 
    -8.041934e-007, -4.060839e-007, -6.646196e-007, -1.184793e-006, 
    -1.10768e-006, -1.532859e-006, -5.912289e-007,
  -1.148906e-006, -7.757558e-007, -8.046886e-007, 1.060191e-006, 
    -3.046693e-006, -5.79633e-006, 7.877497e-007, 4.933504e-006, 
    1.226836e-006, 9.099379e-007, 1.130982e-007, -2.639146e-006, 
    -1.993057e-006, -2.275682e-006, -1.65977e-006, -2.075263e-006, 
    1.362934e-006, -2.659759e-006, -2.565881e-006, -6.372829e-008, 
    3.463128e-006, 5.886932e-007, -1.697269e-006, -2.789773e-006, 
    -5.37957e-008, -6.62757e-007, -1.093274e-006, -9.271262e-007, 
    -9.221603e-007, -3.919267e-007, 5.19155e-007, 1.600607e-006, 
    2.102278e-006, 3.08265e-006, 2.427621e-006, 1.102287e-006, 1.483644e-007, 
    -2.622866e-007, 1.691255e-006, 3.327651e-006, 7.453411e-006, 
    6.878847e-006, -6.036498e-007, -3.380483e-006, -8.701318e-007, 
    -3.089786e-006, -3.508758e-006, -7.437571e-006, -7.678602e-006, 
    -6.021466e-006, -1.427805e-006, -6.928167e-007, 7.164635e-007, 
    5.221831e-006, 1.081138e-005, 1.056874e-005, 8.354556e-006, 
    6.145587e-006, 4.641191e-006, 3.238616e-006, -5.945831e-007, 
    -1.97828e-006, -1.897563e-006, -2.08768e-006, -1.292206e-006, 
    -1.513861e-006, -2.292447e-006, -2.428545e-006, -2.921648e-006, 
    -3.171737e-006, -2.513106e-006, -2.322994e-006, -2.02286e-006, 
    -9.888431e-007, 1.004436e-006, -1.418221e-008, 4.476773e-006, 
    -3.266607e-006, -5.691407e-006, 6.633592e-006, 6.222446e-006, 
    3.922209e-006, -7.390918e-008, -4.436848e-006, -4.39947e-006, 
    -3.834095e-006, -7.673125e-007, -6.343198e-007, -1.191375e-006, 
    -1.171258e-006, -1.567257e-006, -1.438983e-006, -1.337407e-006, 
    -1.084955e-006, -1.520564e-006, -4.654394e-007,
  -1.768918e-006, -3.108398e-007, -1.61643e-006, 1.427752e-007, 
    -5.097216e-006, -6.507858e-006, 4.51415e-006, 4.554884e-006, 
    3.336966e-006, -4.497861e-008, -5.764377e-008, -2.048191e-006, 
    -3.957402e-006, -7.219516e-006, -1.13367e-005, -3.068799e-006, 
    4.427351e-006, 3.544334e-006, 2.468598e-006, -2.22055e-007, 
    2.784753e-006, -1.89508e-006, 3.567437e-006, 7.492277e-006, 
    2.967787e-006, 1.205104e-006, 1.321831e-006, 1.013625e-006, 
    9.680521e-007, 3.620726e-007, 3.020687e-006, 4.039306e-006, 
    5.139509e-006, 4.39768e-006, 6.117521e-006, 2.11631e-006, 3.17715e-006, 
    3.925064e-006, 3.323926e-006, 5.048361e-006, 8.668845e-006, 
    7.962153e-006, 1.607968e-005, 8.359646e-006, -1.883161e-005, 
    -2.397277e-005, -1.851858e-005, -1.710781e-005, -1.238663e-005, 
    2.882349e-006, 1.258327e-005, 1.955315e-005, 1.835608e-005, 
    1.763723e-005, 1.912561e-005, 1.419903e-005, 8.571989e-006, 
    6.164586e-006, 2.778293e-006, 1.309164e-006, -1.347835e-006, 
    -1.240795e-006, -1.396636e-006, -7.363924e-007, -1.962386e-006, 
    -1.743463e-006, -2.493116e-006, -3.123931e-006, -3.694025e-006, 
    -3.394385e-006, -2.574822e-006, -2.63716e-006, -1.878815e-006, 
    4.553281e-007, 2.886204e-006, 9.225652e-006, -1.969737e-005, 
    -5.69947e-006, 6.278207e-006, 1.797416e-006, 5.796148e-006, 
    2.955616e-006, -2.80219e-006, -1.456615e-006, -7.272042e-007, 
    -1.180943e-006, -1.471143e-006, -3.105915e-007, -1.09191e-006, 
    -1.006724e-006, -1.710929e-006, -1.539938e-006, -1.69727e-006, 
    -1.782701e-006, -1.552354e-006, -7.695476e-007,
  -2.022611e-006, -1.313316e-006, -1.840072e-006, -1.593706e-006, 
    -6.354378e-006, -1.380955e-005, -1.987137e-007, 3.937232e-006, 
    2.771838e-006, 1.397702e-006, -1.594948e-006, -3.550477e-006, 
    -5.871083e-006, -7.739065e-006, -1.465632e-005, -1.584455e-005, 
    -4.913192e-006, 7.196235e-006, 1.271513e-005, 3.398549e-006, 
    9.951327e-007, -6.045557e-006, 6.15005e-006, 1.128326e-005, 1.1058e-005, 
    7.383621e-006, 6.250513e-006, 9.53684e-006, 3.025655e-006, 3.34727e-006, 
    5.607157e-006, 6.09455e-006, 5.741392e-006, 6.021286e-006, 5.382895e-006, 
    9.104953e-006, 1.453655e-005, 2.487871e-005, 1.755701e-005, 
    4.018071e-006, 1.13205e-005, 4.972731e-006, 4.206078e-006, 1.219024e-005, 
    -1.909015e-005, -9.022071e-006, 6.995455e-006, 1.897139e-005, 
    2.611449e-005, 4.037056e-005, 4.76555e-005, 4.164399e-005, 3.562219e-005, 
    2.73364e-005, 1.834691e-005, 1.207165e-005, 7.655818e-006, 4.228178e-006, 
    1.837907e-006, -1.921271e-007, -5.066663e-007, -9.725754e-007, 
    -1.80915e-006, -3.015276e-006, -2.486036e-006, -2.662862e-006, 
    -3.180679e-006, -3.461193e-006, -3.188005e-006, -3.101454e-006, 
    -2.308837e-006, -1.770285e-006, 1.86486e-007, 1.914028e-006, 
    1.778551e-006, 2.676337e-006, 1.309414e-006, 1.042855e-005, 
    -1.286916e-005, -1.051949e-005, 1.536526e-006, 2.695095e-006, 
    4.313615e-007, -5.601851e-007, 3.157541e-007, -5.044305e-007, 
    -1.116993e-006, -7.602284e-008, -2.209363e-007, -1.295309e-006, 
    -1.170638e-006, -2.04546e-006, -1.539938e-006, -1.460463e-006, 
    -1.802196e-006, -1.499952e-006,
  1.42652e-007, 3.304067e-007, 4.040298e-006, 2.621215e-006, 2.697579e-006, 
    6.607392e-006, 2.990644e-006, -8.475181e-006, 2.577437e-005, 
    9.784071e-006, 6.399769e-007, -2.851239e-006, -8.217892e-006, 
    -8.869822e-006, -1.036627e-005, -2.176018e-005, -7.948423e-006, 
    -3.790767e-006, -8.091367e-006, -1.064381e-005, -4.137095e-006, 
    -8.293769e-006, -3.766618e-007, 1.438431e-005, 1.675955e-005, 
    5.271264e-006, 9.720989e-006, 1.035727e-005, 1.21916e-005, 8.904783e-006, 
    4.080532e-006, 6.646631e-006, 9.980518e-006, 1.84142e-005, 2.119974e-005, 
    6.328741e-006, 7.269751e-006, -9.559735e-006, -4.781105e-007, 
    7.338294e-006, -6.389237e-007, -1.130276e-006, 9.697651e-006, 
    3.121029e-006, 2.486107e-006, 1.929845e-005, 4.061916e-005, 
    4.232523e-005, 4.553742e-005, 3.530442e-005, 2.105768e-005, 
    9.985242e-006, 5.126843e-006, 3.306168e-006, 1.945941e-006, 
    8.611364e-007, 8.019151e-008, -1.50528e-007, -1.287974e-007, 
    -7.642079e-007, -7.157794e-007, -8.822992e-007, -1.467791e-006, 
    -8.754696e-007, -1.154991e-006, -1.238437e-006, -1.573713e-006, 
    -1.870867e-006, -9.568057e-007, -5.713619e-007, 6.105483e-007, 
    2.650766e-006, 3.546326e-006, 7.576841e-006, 8.404229e-006, 
    6.145456e-006, 2.59513e-006, 2.219247e-006, -1.471667e-005, 
    -5.033522e-006, -7.801282e-008, -2.674289e-006, -9.479886e-007, 
    -5.66022e-007, -3.366684e-007, 1.306061e-006, 2.427497e-006, 
    4.547063e-006, 3.841616e-006, 1.478417e-006, 8.638685e-007, 
    -9.268788e-007, -7.797303e-007, -4.943727e-007, -1.245267e-006, 
    -5.958245e-007,
  1.327082e-005, 1.803211e-005, 2.65312e-006, -1.470027e-006, 6.81886e-006, 
    -8.089046e-007, -4.609705e-006, -3.182286e-006, 3.139648e-005, 
    2.511563e-005, 9.507288e-006, -1.828027e-006, -5.422187e-006, 
    -2.659268e-006, 6.072441e-006, 8.275209e-006, 1.374294e-005, 
    -8.238509e-006, -2.138704e-005, -1.522243e-005, -4.933929e-006, 
    -3.606401e-007, -5.151487e-006, -8.541003e-006, -5.73822e-006, 
    -8.964569e-006, -7.995986e-006, 2.080778e-007, 2.352591e-005, 
    1.739968e-005, 5.55376e-006, 8.692565e-006, 6.226059e-006, 1.619269e-005, 
    1.867249e-005, 7.510418e-006, 3.181376e-006, 4.609894e-006, 
    1.441609e-005, 1.419384e-005, 4.373724e-006, 2.065013e-005, 
    3.243061e-005, 3.064619e-005, 3.26566e-005, 4.208631e-005, 5.202601e-005, 
    4.271986e-005, 4.33246e-005, 3.676921e-005, 2.271754e-005, 1.130064e-005, 
    8.575095e-006, 5.857868e-006, 3.947042e-006, 2.311641e-006, 
    1.326301e-006, 1.167604e-006, 1.296499e-006, 1.006795e-006, 
    4.903461e-007, -5.074107e-007, -2.449021e-007, -3.646078e-007, 
    -1.989565e-007, 4.819021e-007, 4.647654e-007, 9.95246e-007, 
    2.457795e-006, 4.298464e-006, 6.778261e-006, 6.480241e-006, 
    8.994315e-006, 1.49323e-005, 1.096163e-005, -1.96667e-005, 
    -2.028522e-005, 1.459539e-006, -5.582748e-006, -5.85855e-006, 
    -9.176911e-007, -7.767496e-007, -3.263257e-006, -1.831504e-006, 
    -1.459347e-006, -1.443204e-006, 6.429946e-008, 4.273999e-006, 
    3.420411e-006, 3.419666e-006, 3.044155e-006, 4.830435e-006, 
    7.030715e-006, 7.792412e-006, 8.152898e-006, 9.859577e-006,
  -5.34732e-007, 1.635373e-006, 1.573659e-006, -1.37204e-005, -5.691327e-007, 
    6.941053e-006, 5.338683e-006, -7.086273e-006, -1.312445e-006, 
    4.405447e-007, 5.334965e-006, 8.334435e-006, 4.037443e-006, 
    2.935129e-006, 7.049959e-006, 1.54038e-005, 2.187561e-005, 2.280769e-005, 
    2.725382e-005, 2.89641e-005, 9.711308e-006, -5.668182e-006, 
    -1.731804e-005, -2.169165e-005, -2.293429e-005, -1.460304e-005, 
    -4.551588e-006, 1.266199e-006, 1.07524e-005, 6.912014e-006, 
    3.843226e-006, -1.541681e-006, 6.309747e-006, 1.289828e-005, 
    1.313546e-005, 5.724753e-006, 4.290523e-006, 9.095143e-006, 
    1.177711e-005, 1.406095e-005, 1.362064e-005, 1.604468e-005, 
    1.851625e-005, 1.233278e-005, 4.617454e-006, 5.532522e-006, 
    2.957057e-005, 3.210924e-005, 4.690845e-005, 5.290232e-005, 
    5.403059e-005, 4.971546e-005, 4.984063e-005, 4.170869e-005, 3.56243e-005, 
    2.66394e-005, 2.094815e-005, 1.965373e-005, 1.676216e-005, 1.349247e-005, 
    1.192735e-005, 1.141401e-005, 1.01684e-005, 2.455185e-006, 4.325029e-006, 
    6.306142e-006, 3.240475e-006, 5.91101e-006, 4.661269e-007, 
    -2.040128e-006, 3.069486e-006, -2.496847e-006, 9.826777e-006, 
    1.351196e-005, -1.172375e-005, 3.53888e-007, -4.644353e-006, 
    5.900583e-007, 2.880624e-007, -7.603465e-006, -8.100285e-007, 
    -6.046409e-007, -2.168518e-006, 3.255591e-007, 1.486231e-006, 
    -9.003124e-007, -1.328714e-006, 9.786017e-007, -4.299764e-006, 
    -3.183915e-006, -9.765259e-006, -3.243636e-006, -3.920526e-006, 
    -8.116062e-006, 1.443899e-006, 2.713845e-006,
  -3.859714e-007, -5.624242e-007, -3.643581e-007, -3.095369e-006, 
    -3.136967e-006, 1.671015e-006, 3.166962e-006, 9.211726e-008, 
    -3.803794e-006, -1.717561e-005, 5.620816e-006, 8.159106e-006, 
    1.106048e-005, 1.200484e-005, 3.337085e-006, 8.847284e-006, 
    2.683758e-005, 3.26345e-005, 3.370143e-005, 3.190708e-005, 2.729753e-005, 
    1.505759e-005, -1.152186e-005, -1.634374e-005, -1.180796e-005, 
    -1.347254e-005, -1.21944e-005, -1.161578e-006, 7.209645e-006, 
    -9.586562e-006, -1.106489e-005, -5.249094e-007, 1.821527e-005, 
    2.587484e-005, 7.105831e-006, 4.736925e-006, 4.589907e-006, 
    1.146371e-006, -2.734596e-007, 7.40424e-006, 6.201837e-006, 
    -5.460053e-006, 4.025904e-006, 5.389971e-006, 8.193994e-006, 
    8.463976e-006, 1.272607e-005, 1.774143e-005, 1.746551e-005, 
    1.841482e-005, 1.127207e-005, -3.005407e-007, -2.933448e-006, 
    -9.827971e-006, -5.384078e-006, -2.629095e-006, 4.59524e-006, 
    9.467061e-006, 1.015064e-005, 4.480375e-006, 7.504445e-006, 
    6.569266e-006, -2.903151e-006, -1.055117e-005, -4.351918e-006, 
    -7.877163e-006, -9.448857e-006, 3.453191e-006, 1.905828e-006, 
    8.632589e-006, 2.108127e-005, 2.606322e-005, 2.110511e-005, 
    2.927918e-006, -4.297079e-005, -2.180167e-005, 1.014196e-007, 
    -9.878495e-007, -5.832093e-006, -6.473711e-006, -9.114072e-006, 
    -6.316004e-006, -7.008166e-006, -1.497607e-005, -1.653648e-005, 
    -8.862e-006, -1.299483e-005, -9.643561e-006, -7.933901e-006, 
    -4.522655e-006, -1.043928e-005, -1.553238e-005, -1.106427e-005, 
    -7.101917e-007, -7.362723e-007, 7.124618e-008,
  -1.251477e-006, -1.397259e-006, -9.731971e-007, -1.81921e-006, 
    -2.04608e-006, -1.245267e-006, -2.291329e-006, -2.418361e-006, 
    -4.884501e-006, -5.400455e-006, 2.893034e-006, 2.439045e-006, 
    8.470787e-006, 1.174606e-005, 1.350502e-005, 2.119004e-005, 
    2.312894e-005, 2.715758e-005, 2.988536e-005, 2.838295e-005, 
    2.256518e-005, 2.109478e-006, -2.495563e-005, -1.600201e-005, 
    -6.341219e-006, -1.646853e-005, -1.947174e-005, -6.764094e-007, 
    -2.345965e-006, -8.532188e-006, -8.457049e-006, -6.896284e-006, 
    3.075205e-006, 2.905289e-005, 7.120383e-006, 9.623327e-007, 4.54644e-006, 
    -1.923894e-006, -4.942616e-006, -2.595072e-006, -2.280649e-006, 
    2.101784e-006, 8.430179e-006, 2.053937e-005, 2.045256e-005, 
    -5.466391e-006, 8.369832e-006, 2.311267e-005, 1.413223e-005, 
    5.322676e-006, -8.938609e-006, 3.227033e-007, -3.179441e-006, 
    6.49377e-006, 1.179027e-005, 8.165181e-006, 2.984671e-006, 7.625513e-006, 
    1.529663e-005, 7.034312e-006, 5.060774e-006, 4.194648e-006, 
    -3.100962e-006, -2.250479e-006, 4.704889e-006, 5.558104e-006, 
    4.161244e-006, 1.483531e-005, 1.662619e-005, 2.364898e-005, 
    3.363586e-005, 2.62285e-005, 5.884318e-006, -1.344683e-005, 
    -3.365654e-005, -2.418037e-005, -8.487856e-006, -4.621867e-006, 
    -7.840768e-006, -1.314062e-005, -1.077282e-005, -9.030251e-006, 
    -2.048925e-005, -1.589695e-005, -8.329029e-006, -6.949927e-006, 
    -4.321861e-006, -2.865521e-006, -3.658386e-006, -5.132109e-006, 
    -8.015857e-006, -7.690895e-006, -2.401472e-006, -5.005822e-007, 
    -1.47251e-006, -4.712765e-007,
  -3.699474e-007, -4.374995e-007, -3.31453e-007, -1.142686e-007, 
    -4.684074e-008, 2.555286e-007, 2.24112e-007, -2.90599e-007, 
    -2.951934e-007, -2.107795e-006, 2.456045e-008, 1.659342e-006, 
    5.651486e-006, 8.833009e-006, 1.069863e-005, 1.383831e-005, 
    1.450154e-005, 2.157362e-005, 3.022425e-005, 2.743761e-005, 
    1.334768e-005, -6.033504e-006, -2.519889e-005, -2.056413e-005, 
    -1.258902e-005, -4.433125e-006, 3.293504e-006, -3.764557e-006, 
    -5.873568e-006, 3.803747e-006, 1.245163e-005, 2.354469e-005, 
    -1.40193e-005, -1.599299e-006, 1.773442e-006, -6.136543e-008, 
    -2.527515e-006, -4.740832e-006, -5.545116e-006, 4.419126e-007, 
    -5.219285e-006, 1.200956e-005, 1.119198e-005, 4.706751e-006, 
    -1.692431e-006, -1.336542e-006, 6.863935e-006, -4.403628e-007, 
    -7.931922e-006, -2.387693e-006, -3.997891e-006, -9.478681e-007, 
    1.264085e-006, 3.505218e-006, 6.641047e-006, 4.322923e-006, 
    -2.260313e-007, -2.11077e-006, 5.273372e-006, -5.221864e-007, 
    -1.358883e-006, -2.6158e-006, 1.262633e-007, -4.845631e-006, 
    1.750232e-006, 6.107955e-006, 1.345857e-005, 1.153347e-005, 1.05192e-005, 
    4.174535e-006, -4.043332e-006, -1.257101e-005, -1.845598e-005, 
    -2.227011e-006, -8.629046e-006, -2.532353e-006, -7.524246e-006, 
    -7.732982e-006, -5.16924e-006, -6.575039e-006, -6.483395e-006, 
    -8.499399e-006, -1.013729e-005, -7.092855e-006, -6.881259e-006, 
    -4.755485e-006, -2.344476e-006, -2.53198e-006, -2.175844e-006, 
    -2.772388e-006, -5.729522e-006, -4.310187e-006, -1.980267e-006, 
    -1.631952e-006, -8.241848e-007, 3.312857e-008,
  -1.319014e-007, -4.274413e-007, -1.982117e-007, -1.121574e-007, 
    5.933003e-008, -5.689904e-008, 1.301105e-007, 1.071379e-007, 
    9.286921e-009, -3.670915e-007, -2.829509e-006, 2.314248e-006, 
    1.985553e-006, 2.700436e-006, 5.6721e-006, 1.114741e-005, 1.382403e-005, 
    1.856483e-005, 2.494873e-005, 2.275578e-005, 5.067859e-006, 
    -2.214709e-006, -9.664676e-006, -2.014167e-006, -6.600007e-006, 
    -5.993061e-007, 6.521215e-006, 2.102404e-006, 7.020036e-006, 
    8.02636e-006, 1.048182e-005, 1.470593e-005, 8.082119e-006, 3.205962e-006, 
    -3.629451e-006, -1.181255e-005, -1.496712e-005, 6.007322e-007, 
    -5.707552e-007, 4.527072e-006, -3.313304e-006, 7.174014e-006, 
    6.165945e-006, -2.440465e-006, 2.541241e-006, -5.002843e-006, 
    -5.024205e-006, -9.377705e-006, -4.114241e-006, -6.408991e-007, 
    -5.58039e-006, -8.365416e-006, 6.094342e-008, -8.898751e-007, 
    -1.413391e-007, 1.820898e-006, 3.561399e-008, -3.553083e-006, 
    -2.692293e-006, 4.559515e-007, -1.181192e-006, -2.289342e-006, 
    -5.422808e-006, -5.898156e-006, -3.628459e-006, -6.490969e-006, 
    -7.564362e-006, 6.65932e-007, -4.321113e-006, -4.763553e-006, 
    -1.553099e-006, -6.560264e-006, -3.720721e-006, 1.229703e-005, 
    9.689822e-006, 1.396037e-005, 1.502878e-006, -3.677265e-006, 
    -2.431774e-006, -1.755383e-006, -2.075263e-006, -3.31839e-006, 
    -5.557413e-006, -4.644842e-006, -3.773498e-006, -3.67577e-006, 
    -4.031908e-006, -2.809391e-006, -1.591595e-006, -2.082712e-006, 
    -1.522056e-006, -5.225602e-007, -1.136613e-006, -8.181003e-007, 
    -4.125286e-008, 2.331888e-008,
  -3.120815e-007, -2.789262e-007, -1.059002e-006, -2.275173e-007, 
    -2.268965e-007, -1.343851e-007, -1.590962e-007, -4.746167e-008, 
    1.673752e-008, -1.640586e-009, 2.667161e-008, 1.206223e-006, 
    1.251919e-006, 8.581565e-007, 2.878009e-006, 5.007881e-006, 
    6.650114e-006, 1.075712e-005, 1.06779e-005, 1.026402e-005, 1.156116e-005, 
    8.391688e-006, 2.788231e-006, -1.555334e-006, -2.862544e-006, 
    -2.31492e-006, 1.983814e-006, 3.997091e-006, 3.787727e-006, 
    3.213161e-006, -1.459844e-006, 1.212183e-006, 4.146965e-006, 
    3.799767e-006, 7.038034e-007, -4.094127e-006, -4.517937e-006, 
    -1.331384e-005, -9.841009e-006, 8.044233e-006, 1.517903e-006, 
    6.590129e-006, 6.642291e-006, 5.028989e-006, -3.616296e-007, 
    -5.077854e-007, -6.510716e-006, -4.963598e-006, -9.987762e-007, 
    -4.620875e-006, -8.852683e-006, -1.049937e-006, 1.5641e-006, 
    4.157482e-008, 2.001823e-006, 1.845359e-006, -2.745313e-006, 
    1.524859e-008, 9.722735e-007, 3.726262e-006, -4.152735e-007, 
    -2.509631e-006, -7.165227e-007, 5.307024e-007, 8.842339e-007, 
    -7.853061e-006, -1.088247e-005, -5.773233e-006, -9.637602e-006, 
    -3.253448e-006, -3.835214e-006, 2.085264e-006, 6.011218e-006, 
    9.684481e-006, 1.120081e-005, 6.265167e-006, 3.582209e-006, 
    3.825218e-006, 5.897105e-006, 6.668117e-006, 7.231876e-006, 3.61698e-006, 
    6.163864e-007, -2.035275e-006, -2.634552e-006, -4.627706e-006, 
    -3.379238e-006, -1.552232e-006, -2.362853e-006, -2.782445e-006, 
    -7.955005e-007, -5.27155e-007, -1.034415e-006, -1.001757e-006, 
    -1.076263e-006, -2.827758e-007,
  -2.753252e-007, -1.857939e-007, -8.061659e-008, -8.475297e-007, 
    -8.937233e-007, -5.369647e-007, -3.221397e-007, -2.367064e-007, 
    -3.342974e-008, 6.678057e-008, -1.109158e-007, 1.292413e-007, 
    3.533796e-007, 6.183719e-007, 2.278113e-006, 1.680204e-006, 
    2.894285e-007, 1.106385e-006, 3.671744e-006, 7.590128e-006, 
    6.350227e-006, 8.423972e-006, 1.703549e-006, 1.679833e-006, 
    7.260278e-007, -1.219812e-005, 2.139408e-006, 2.175293e-007, 
    1.645309e-006, 6.643906e-006, 2.785992e-006, 5.089723e-007, 
    -9.532032e-007, -9.812684e-007, -9.771684e-007, 6.386072e-007, 
    5.927403e-006, -3.158832e-006, -3.916677e-006, -3.194218e-006, 
    -2.207882e-006, 8.406834e-006, 1.635934e-005, 1.234025e-005, 
    7.114035e-006, 2.756195e-006, -1.220906e-007, 1.113467e-006, 
    -2.510933e-008, -3.95293e-006, -2.018014e-006, -1.072536e-006, 
    -4.557514e-007, 2.100805e-007, -1.042099e-007, -9.129708e-007, 
    -2.371546e-006, -8.985662e-007, -1.77637e-006, -2.040741e-006, 
    -1.16207e-006, -1.581783e-006, 2.218762e-007, -3.966452e-007, 
    1.114332e-006, 1.529588e-007, -3.10964e-007, -2.031676e-006, 
    -4.861529e-006, -3.342232e-006, -8.583347e-007, 4.630627e-006, 
    2.229899e-007, -2.195837e-006, -1.470507e-007, -4.623987e-006, 
    -3.75673e-006, -1.651861e-007, 4.256981e-006, 3.037323e-006, 
    7.11664e-006, 6.644521e-006, 3.672114e-006, 1.196788e-006, 
    -1.142671e-007, -4.828997e-006, -3.959887e-006, -3.734506e-006, 
    -3.387433e-006, -2.3446e-006, -1.688328e-006, -5.649049e-007, 
    -1.026717e-006, -4.310423e-007, -5.514935e-007, -9.82137e-007,
  -1.323125e-006, -1.1309e-006, -9.216629e-007, -1.347576e-007, 
    -1.191498e-006, -1.397259e-006, -1.188021e-006, -1.595071e-006, 
    -7.208703e-007, 2.294632e-008, 7.373438e-008, -6.225222e-007, 
    -1.070532e-008, 1.740689e-007, 1.476554e-006, 1.761291e-006, 
    4.67001e-007, -1.270588e-007, 2.835416e-006, 3.50187e-006, 2.204228e-006, 
    3.850805e-006, 3.352487e-006, 2.08713e-006, 3.699436e-006, 3.779282e-006, 
    2.532675e-006, 1.10874e-006, 1.600602e-006, 4.950387e-006, 7.854627e-006, 
    6.961052e-006, 2.636611e-006, -8.446732e-007, -4.354517e-006, 
    -7.069648e-007, 7.613839e-006, 9.568004e-006, 2.840006e-006, 
    3.160629e-006, 3.55874e-006, 1.218838e-005, 1.63006e-005, 1.136906e-005, 
    1.262486e-005, 1.234596e-005, 6.537488e-006, 4.295609e-006, 
    7.753315e-007, 1.816054e-006, 2.993867e-006, 3.403647e-006, 
    1.753717e-006, 1.853803e-006, 1.752973e-006, -2.196581e-006, 
    -1.25632e-006, -1.049557e-007, 8.426332e-007, -1.082844e-006, 
    -1.84392e-006, -2.519191e-006, -1.246881e-006, -3.236296e-007, 
    2.837168e-007, 3.120288e-007, 3.317728e-007, 8.46484e-007, 
    -2.295799e-006, -1.021624e-006, 2.652132e-007, -1.502809e-006, 
    -9.868545e-007, -4.224879e-006, -4.218915e-006, -9.838805e-007, 
    -2.836096e-006, -5.455717e-006, -4.605979e-006, -2.743363e-007, 
    1.119788e-006, 3.646906e-006, -2.465204e-007, -2.892968e-006, 
    -2.826651e-006, -3.670553e-006, -5.254671e-006, -5.367301e-006, 
    -3.929463e-006, -2.801569e-006, -2.193104e-006, -1.396887e-006, 
    -2.362233e-006, -1.969835e-006, -1.760723e-006, -3.639015e-006,
  -1.802074e-006, -3.571337e-006, -4.202526e-006, -1.761095e-006, 
    -1.486913e-006, -4.455473e-006, -4.553822e-006, -2.951574e-006, 
    -7.414837e-007, 5.673346e-007, -2.175716e-008, -1.546258e-007, 
    -6.025221e-008, -8.136203e-008, 3.013492e-007, 1.483509e-006, 
    1.863737e-006, 1.375723e-006, 1.443151e-006, 2.191809e-006, 
    1.548949e-006, 1.546589e-006, 6.776036e-007, -1.109156e-007, 
    6.557493e-007, 2.411974e-006, 2.751225e-006, 7.610119e-006, 
    8.537092e-006, 6.534257e-006, 6.22779e-006, 5.043275e-006, 3.80126e-006, 
    1.812205e-006, 2.390152e-007, 1.936009e-006, 3.49839e-006, 5.852151e-006, 
    9.540163e-007, -1.507411e-006, -1.069562e-006, -7.052295e-007, 
    9.995416e-006, 1.15634e-005, 1.266422e-005, 1.277461e-005, 7.872997e-006, 
    7.026614e-006, 7.352453e-006, 4.898859e-006, 2.033115e-006, 7.2494e-008, 
    -1.579423e-006, -2.97674e-007, -5.026923e-007, -1.931838e-006, 
    -3.509496e-006, -1.487879e-007, -1.052047e-006, -1.577314e-006, 
    -1.824302e-006, -1.793877e-006, -1.184545e-006, -1.682854e-007, 
    -1.825654e-007, 1.326089e-008, 1.447629e-007, -2.15472e-007, 
    1.315125e-006, -1.939662e-006, -5.125003e-007, 2.503492e-006, 
    4.343383e-008, 3.635432e-008, -8.931056e-008, 2.326815e-007, 
    -2.41811e-006, -2.349199e-006, -4.530975e-006, -4.1618e-006, 
    -5.047921e-006, -5.643971e-006, -2.469031e-006, -3.822923e-006, 
    -3.273442e-006, -4.728663e-006, -5.983586e-006, -3.117346e-006, 
    -3.982112e-006, -3.048181e-006, -4.100577e-006, -3.979754e-006, 
    -3.850486e-006, -2.035276e-006, -4.285474e-006, -3.046071e-006,
  -7.697963e-007, -1.644494e-006, 1.038587e-006, 2.116065e-006, 
    -1.569842e-007, -5.815577e-006, -4.293298e-006, -2.277048e-006, 
    -2.724952e-006, -3.442317e-006, -2.4366e-007, 1.239626e-006, 
    1.935138e-006, 2.536274e-006, 1.075093e-006, 1.020455e-006, 
    1.047774e-006, 7.760759e-007, 4.681185e-007, 5.495776e-007, 
    3.330151e-007, 1.586202e-006, 1.546466e-006, 2.388258e-006, 
    2.631519e-006, 2.332129e-006, 3.418051e-006, 8.106454e-006, 
    1.164995e-005, 1.058526e-005, 7.134153e-006, 5.622805e-006, 
    6.626151e-006, 7.348606e-006, 5.837379e-006, -9.221567e-007, 
    -1.084334e-006, 1.678345e-006, 2.613262e-006, -2.407935e-006, 
    -7.364062e-006, -8.514311e-006, -5.257658e-006, 5.250025e-006, 
    1.256054e-005, 1.302136e-005, 1.182839e-005, 7.930743e-006, 
    3.222842e-006, 3.739788e-006, 1.242355e-006, 7.857561e-007, 
    2.164241e-006, 8.246279e-007, -3.2229e-006, -3.845271e-006, 
    -1.959907e-006, 1.08068e-006, 2.933519e-006, 2.811827e-006, 
    2.418185e-006, 3.738696e-007, 1.688895e-006, 3.899854e-006, 
    4.568048e-006, 2.195784e-006, 1.658224e-006, 2.338587e-006, 
    1.528088e-006, 1.042682e-006, 3.658212e-006, 2.623945e-006, 
    3.241597e-006, 3.20596e-006, 1.087759e-006, -1.792387e-006, 
    -4.673653e-006, 8.400275e-007, 3.459274e-006, -2.531986e-006, 
    -3.106921e-006, -5.068658e-006, -9.375719e-006, -1.04106e-005, 
    -9.775809e-006, -8.059691e-006, -7.741299e-006, -4.054506e-006, 
    -1.395641e-006, -9.414052e-007, -3.472214e-007, -4.517933e-006, 
    -3.94573e-006, -2.66485e-006, -4.921383e-006, -3.521791e-006,
  8.566658e-007, 2.469222e-006, 1.51679e-006, -1.097746e-006, -3.597634e-007, 
    -2.844285e-006, -7.749622e-006, -2.397746e-006, -9.166952e-007, 
    -3.206136e-006, -3.602754e-006, -3.947469e-006, -1.677773e-006, 
    -1.265626e-007, -9.71334e-007, -1.399121e-006, -6.153191e-007, 
    -2.11498e-007, 7.219348e-007, 1.335863e-006, 8.84731e-007, 1.143017e-006, 
    1.737821e-006, 1.191446e-006, 9.573733e-007, 1.390376e-006, 
    1.983318e-006, 3.226696e-006, 6.289132e-006, 7.066599e-006, 
    7.327249e-006, 7.573488e-006, 7.447821e-006, 7.546669e-006, 
    7.606772e-006, 4.582331e-006, 1.939236e-006, 3.68019e-006, 2.837904e-006, 
    2.226952e-006, 3.021927e-006, -1.234344e-006, 7.194467e-007, 
    1.706896e-006, 3.950146e-006, 5.262933e-006, 5.06264e-006, 6.760005e-006, 
    1.178096e-005, 1.052889e-005, 1.043426e-005, 8.763214e-006, 
    5.774295e-006, 6.392194e-006, 7.399267e-006, 4.700043e-006, 
    1.932029e-006, 2.147353e-006, 4.550908e-006, 6.989361e-006, 
    8.642895e-006, 6.914979e-006, 7.343267e-006, 9.136125e-006, 
    9.612215e-006, 7.675191e-006, 5.496887e-006, 2.89055e-006, 1.53206e-006, 
    7.528542e-007, 4.317958e-006, 3.669385e-006, 5.499496e-006, 
    6.143351e-006, 4.556377e-006, 1.869574e-006, -6.86472e-007, 
    -1.782826e-006, -1.181686e-006, -4.653139e-007, 2.804496e-006, 
    5.123118e-006, 4.212776e-006, 8.195348e-007, -2.208253e-006, 
    -1.765566e-006, -3.619272e-006, -3.743073e-006, 8.683382e-007, 
    2.063165e-006, -1.769731e-007, 6.612136e-007, -1.905119e-007, 
    -4.830708e-007, -3.566121e-006, -2.182423e-006,
  -1.276681e-006, 1.240373e-006, -5.455331e-007, -2.808398e-006, 
    -5.560869e-007, -4.826388e-006, -5.74467e-006, -1.786676e-006, 
    -1.167905e-006, -2.737121e-006, -1.229123e-006, 2.758925e-007, 
    4.483736e-007, 4.011881e-007, 1.676117e-007, 4.513545e-007, 6.12039e-007, 
    1.079563e-006, 1.902113e-007, 8.616335e-007, 2.229311e-006, 
    2.647039e-006, 2.631393e-006, 2.624068e-006, 1.714352e-006, 
    1.428994e-006, 1.304446e-006, 1.08751e-006, 1.251174e-006, 1.951529e-006, 
    2.655609e-006, 3.237624e-006, 3.038692e-006, 2.473192e-006, 
    2.303444e-006, 4.567799e-006, 4.239231e-006, 3.086006e-006, 
    4.560472e-006, 1.591419e-006, 3.609774e-006, 7.62154e-006, 7.670591e-006, 
    1.019708e-005, 1.349545e-005, 1.308666e-005, 7.499351e-006, 
    6.564303e-006, 5.152913e-006, 8.243733e-007, 2.827343e-006, 
    4.769459e-006, 3.613877e-006, 2.034845e-006, 4.236001e-006, 2.58979e-006, 
    -6.946721e-007, -3.579786e-006, 2.519228e-007, 4.045884e-006, 
    6.574486e-006, 1.359517e-005, 1.721268e-005, 1.598483e-005, 1.38177e-005, 
    9.940537e-006, 6.539971e-006, 5.024396e-006, 5.126592e-006, 
    2.763019e-006, 2.742904e-006, 3.357331e-006, 1.465503e-006, 
    3.107241e-006, 5.797769e-006, 5.031356e-006, 2.922712e-006, 
    4.448339e-006, 2.191686e-006, -2.297493e-007, 8.652569e-008, 
    1.860135e-006, 4.332978e-006, 1.16754e-005, 7.882685e-006, 4.260583e-006, 
    2.902925e-007, -7.828385e-007, 1.785338e-007, 2.356592e-006, 
    4.712707e-006, 4.879854e-006, 3.685775e-006, 3.128103e-006, 
    1.208335e-006, 9.825835e-007,
  -3.171717e-007, -1.11277e-006, 8.684619e-007, 1.460066e-007, 
    -8.198385e-007, -2.813118e-006, -2.320883e-006, -2.510003e-006, 
    -2.265997e-006, -1.74098e-006, -1.051304e-006, -7.707895e-007, 
    -5.030633e-007, 5.6299e-007, 1.412604e-006, 4.837639e-007, 7.934614e-007, 
    1.140036e-006, 6.161363e-007, 5.28592e-007, 1.884721e-006, 2.2123e-006, 
    2.994485e-006, 3.96865e-006, 1.586202e-006, 1.129233e-006, 8.478482e-007, 
    1.756835e-007, 1.221991e-006, 1.582104e-006, 1.311772e-006, 
    1.472581e-006, 1.737821e-006, 1.514305e-006, 1.339959e-006, 
    1.726272e-006, 3.185343e-006, 3.1697e-006, 1.419437e-006, 1.137681e-006, 
    2.471577e-006, 3.730227e-006, 7.864677e-006, 7.570754e-006, 
    8.615447e-006, 1.120775e-005, 1.282254e-005, 1.175202e-005, 
    9.606625e-006, 1.024899e-005, 8.098377e-006, 5.298694e-006, 
    7.143215e-006, 4.926915e-006, 3.600588e-006, 5.458263e-006, 
    4.438156e-006, 2.636607e-006, 2.069119e-006, 2.202854e-006, 
    3.751091e-006, 8.738505e-006, 1.417445e-005, 1.94825e-005, 1.566183e-005, 
    8.460855e-006, 5.265177e-006, 4.5226e-006, 4.291134e-006, 3.25836e-006, 
    3.030002e-006, 5.023652e-006, 5.667631e-006, 5.655093e-006, 
    8.301657e-006, 6.667249e-006, 4.97522e-006, 6.317314e-006, 4.876125e-006, 
    1.50648e-006, -1.526529e-006, 1.147364e-006, 2.943445e-006, 
    4.137029e-006, 5.678678e-006, 9.008469e-006, 5.428337e-006, 
    1.437365e-008, -2.315923e-006, -2.676315e-007, 5.250396e-006, 
    7.231873e-006, 9.474996e-006, 6.333707e-006, 2.955123e-006, 4.724643e-007,
  2.474064e-006, 1.372124e-006, 1.310409e-006, 2.549441e-006, 9.007508e-007, 
    -1.307102e-006, -9.564319e-007, -1.251352e-006, -2.163426e-006, 
    -1.095634e-006, -1.391424e-006, -1.664239e-006, -5.162283e-007, 
    -1.787175e-007, 6.721393e-007, 1.870319e-006, 3.142255e-006, 
    2.542856e-006, 1.534296e-006, 2.414457e-006, 2.787981e-006, 
    2.592278e-006, 2.317851e-006, 1.015862e-006, 1.041444e-006, 
    1.287184e-006, 1.614514e-006, 6.79217e-007, 1.871067e-007, 1.1717e-006, 
    1.397951e-006, 1.399068e-006, 1.647793e-006, 1.88733e-006, 8.870884e-007, 
    -2.405568e-007, -2.291081e-006, -1.350197e-006, -1.488153e-006, 
    -1.399367e-006, 1.010521e-007, -4.13158e-007, -8.531169e-007, 
    4.729591e-007, 4.029866e-006, 5.045378e-006, 7.333576e-006, 
    9.289477e-006, 9.235213e-006, 1.233515e-005, 1.329118e-005, 
    1.225568e-005, 1.183459e-005, 1.047685e-005, 5.631864e-006, 
    3.664412e-006, 4.149075e-006, 7.569761e-006, 6.289374e-006, 4.87153e-006, 
    5.36364e-006, 8.192997e-006, 9.81264e-006, 8.266637e-006, 6.375802e-006, 
    5.432317e-006, 4.750714e-006, 4.404135e-006, 3.261588e-006, 
    4.428973e-006, 4.926422e-006, 3.202855e-006, 3.243586e-006, 
    6.881455e-006, 8.827796e-006, 7.42597e-006, 8.370822e-006, 6.922306e-006, 
    6.348488e-006, 4.53688e-006, 3.595625e-006, 4.461999e-006, 4.160254e-006, 
    2.871177e-006, 3.635603e-006, 7.701634e-006, 8.376657e-006, 
    3.143992e-006, 6.522641e-007, 1.849574e-006, 6.312803e-007, 
    5.035818e-006, 8.920179e-006, 8.77315e-006, 8.343377e-006, 5.244558e-006,
  1.635373e-006, -1.767185e-006, -3.237557e-006, 2.258494e-007, -1.1345e-006, 
    -1.271714e-006, -7.445888e-007, -2.672095e-008, -2.149736e-007, 
    1.93193e-007, 8.827428e-007, 1.972912e-007, -5.121292e-007, 
    1.628921e-006, 1.767499e-006, 9.692958e-007, 8.464849e-007, 
    2.443267e-006, 2.588553e-006, 2.292889e-006, 2.709252e-006, 
    2.785124e-006, 2.323064e-006, 1.666792e-006, 1.802146e-006, 
    1.374359e-006, 1.597751e-006, 1.932529e-006, 2.944816e-006, 
    3.022054e-006, 3.141015e-006, 3.916371e-006, 2.065894e-006, 
    2.048261e-006, 1.918374e-006, 1.573163e-006, -4.39115e-007, 
    -1.121213e-006, -3.124553e-006, -5.35451e-006, -1.706207e-006, 
    2.057952e-006, 6.712726e-007, -6.107257e-007, 2.496665e-006, 
    5.163223e-006, 7.280058e-006, 7.572613e-006, 8.920924e-006, 
    1.166572e-005, 1.076978e-005, 9.759238e-006, 1.007303e-005, 
    7.850773e-006, 5.998434e-006, 6.653212e-006, 4.86321e-006, 4.933121e-006, 
    2.172434e-006, -2.382345e-006, -4.847381e-006, -3.579116e-007, 
    6.136637e-006, 8.002138e-006, 2.858269e-006, 2.257127e-006, 
    2.315613e-006, 1.867213e-006, 2.150337e-006, 2.821138e-006, 
    3.997955e-006, 6.299193e-006, 6.626024e-006, 5.263933e-006, 
    5.468701e-006, 3.284315e-006, 2.526094e-006, 5.033464e-006, 
    4.229918e-006, 1.807362e-006, 2.605939e-006, 1.792087e-006, 2.6987e-006, 
    3.520745e-006, 2.610159e-006, 4.083638e-006, 3.51913e-006, 5.282182e-006, 
    4.352722e-006, 5.404745e-006, 5.011603e-006, 2.712106e-006, 
    1.803877e-006, 2.131084e-006, 3.274752e-006, 3.001318e-006,
  1.003933e-006, 3.852168e-006, 4.171052e-006, 1.974498e-006, -3.62852e-008, 
    -5.472684e-007, -1.542321e-008, 1.60781e-006, 7.374565e-007, 
    -1.753615e-007, -4.921367e-007, -5.134953e-007, -1.721479e-006, 
    -2.142067e-006, -1.603366e-007, 7.54344e-007, 2.298239e-007, 
    1.101045e-006, 2.622952e-006, 3.151942e-006, 2.038824e-006, 
    1.821267e-006, 2.196282e-006, 3.604939e-006, 4.900967e-006, 
    3.791823e-006, 3.007654e-006, 4.083887e-006, 5.320807e-006, 
    4.428724e-006, 2.007531e-006, 1.425145e-006, 1.524859e-006, 
    1.306681e-006, 1.887081e-006, 1.925574e-006, 1.596385e-006, 
    7.008248e-007, -3.716868e-007, 1.514682e-007, 1.809221e-006, 
    3.580473e-006, 5.286035e-006, 4.493917e-006, 4.389982e-006, 5.81478e-006, 
    6.926655e-006, 5.828315e-006, 3.246068e-006, 2.571045e-006, 
    4.674344e-006, 5.739405e-006, 4.837761e-006, 4.395195e-006, 6.91312e-006, 
    9.320276e-006, 7.948624e-006, 4.831796e-006, 3.234887e-006, 
    5.007714e-007, 9.574906e-007, 6.26067e-007, 2.057577e-006, 3.461888e-006, 
    2.558256e-006, 2.065894e-006, 1.516538e-006, 3.288413e-006, 
    3.449344e-006, 5.065376e-006, 4.253512e-006, 4.258352e-006, 
    4.293993e-006, 5.669245e-006, 6.463975e-006, 6.484588e-006, 6.66092e-006, 
    6.771683e-006, 5.027503e-006, 1.974255e-006, 3.458063e-007, 
    8.744246e-007, 2.831319e-006, 9.948762e-007, 1.200497e-007, 
    6.301671e-007, 1.733206e-007, 3.345776e-006, 5.098402e-006, 
    5.505452e-006, 1.942586e-006, -4.485519e-007, -2.787165e-006, 
    -4.942867e-006, -3.263132e-006, -1.78978e-006,
  -2.969457e-006, -9.8499e-007, 4.067788e-007, 2.168837e-006, 1.533554e-006, 
    1.154318e-006, 1.497418e-006, 2.090483e-006, 2.197276e-006, 
    3.158773e-006, 3.478652e-006, 1.243228e-006, 5.579022e-007, 
    -7.502604e-008, 3.327659e-007, 2.000579e-006, 2.390494e-006, 
    1.824252e-006, 2.309531e-006, 2.946555e-006, 2.945808e-006, 
    3.506339e-006, 2.634996e-006, 2.921721e-006, 4.639327e-006, 
    4.872903e-006, 4.536633e-006, 4.237119e-006, 3.530927e-006, 1.99325e-006, 
    1.366286e-006, 1.02418e-006, 1.600233e-006, 2.78587e-006, 3.767978e-006, 
    3.304182e-006, 2.834049e-006, 2.297483e-006, 2.046026e-006, 
    3.636725e-006, 3.332866e-006, 3.524843e-006, 5.053949e-006, 
    4.991241e-006, 4.72898e-006, 4.224948e-006, 3.143869e-006, 3.730727e-006, 
    4.281824e-006, 4.554888e-006, 3.247433e-006, 1.881245e-006, 1.6617e-006, 
    3.333486e-006, 4.650378e-006, 5.156149e-006, 4.071469e-006, 
    3.699684e-006, 2.740919e-006, 1.947681e-006, 2.270786e-006, 
    1.508467e-006, 2.008649e-006, 2.805366e-006, 3.180627e-006, 3.0341e-006, 
    2.501012e-006, 2.850691e-006, 3.317591e-006, 3.555887e-006, 
    4.881345e-006, 4.991368e-006, 5.668004e-006, 6.74188e-006, 4.383026e-006, 
    3.902835e-006, 4.894881e-006, 5.064383e-006, 3.728866e-006, 
    3.070483e-006, 2.628787e-006, 1.786499e-006, 2.019455e-006, 
    1.509461e-006, -2.603507e-006, -2.44816e-006, -9.032883e-007, 
    -1.099485e-006, -1.290842e-006, 8.168026e-007, 3.326157e-006, 
    1.794197e-006, 7.496292e-007, -5.798047e-007, -2.320012e-006, 
    -2.530738e-006,
  1.298984e-006, 2.031005e-006, 3.927302e-006, 5.038308e-006, 4.95548e-006, 
    4.768346e-006, 3.606552e-006, 2.777551e-006, 1.630659e-006, 
    2.173807e-006, 2.357834e-006, 2.635617e-006, 3.25799e-006, 3.146726e-006, 
    3.273388e-006, 2.90955e-006, 1.732358e-006, 1.111723e-006, 1.43781e-006, 
    2.328278e-006, 2.185476e-006, 2.265446e-006, 2.396577e-006, 
    3.473684e-006, 3.127108e-006, 3.695091e-006, 4.032974e-006, 
    3.105748e-006, 2.295247e-006, 1.767128e-006, 1.660956e-006, 
    2.411851e-006, 3.33361e-006, 3.360061e-006, 2.935999e-006, 1.872801e-006, 
    1.064041e-006, 1.431479e-006, 2.668772e-006, 3.453813e-006, 
    3.230421e-006, 2.763394e-006, 2.372487e-006, 2.431344e-006, 
    2.863976e-006, 2.192555e-006, 2.023552e-006, 2.319339e-006, 
    3.635608e-006, 4.928159e-006, 3.763136e-006, 3.367387e-006, 
    2.666907e-006, 1.131343e-006, 1.982448e-006, 3.540488e-006, 
    2.420543e-006, 6.07567e-007, 7.025628e-007, 2.448606e-006, 3.48759e-006, 
    2.513302e-006, 1.664061e-006, 2.007035e-006, 2.750603e-006, 
    3.666403e-006, 4.716811e-006, 3.879739e-006, 2.385772e-006, 
    2.702173e-006, 3.79207e-006, 4.182853e-006, 4.406867e-006, 3.251159e-006, 
    2.558751e-006, 2.47071e-006, 2.394961e-006, 2.575514e-006, 3.03683e-006, 
    3.354473e-006, 3.518883e-006, 3.198506e-006, 3.422148e-006, 
    3.947415e-006, 1.620227e-006, -3.77895e-007, 4.501126e-007, 
    2.568688e-006, 4.022542e-006, 5.967888e-006, 5.19228e-006, 3.662935e-007, 
    -3.028188e-006, -1.424451e-006, 1.676126e-007, 1.197408e-006,
  1.969662e-006, 1.59415e-006, -1.204753e-007, -4.936264e-007, 1.62867e-006, 
    3.784498e-006, 4.284431e-006, 4.443378e-006, 3.646415e-006, 
    2.014736e-006, 1.054355e-006, 1.606693e-006, 3.030746e-006, 
    4.216758e-006, 4.084755e-006, 3.476664e-006, 3.266928e-006, 
    2.401668e-006, 1.460908e-006, 1.564222e-006, 2.254271e-006, 
    2.421784e-006, 2.537144e-006, 2.871799e-006, 2.658464e-006, 
    2.512557e-006, 2.243219e-006, 2.316234e-006, 2.378944e-006, 
    1.863984e-006, 1.138547e-006, 1.145004e-006, 1.436445e-006, 1.7336e-006, 
    2.289165e-006, 2.470088e-006, 2.096195e-006, 1.728384e-006, 
    1.737449e-006, 2.111965e-006, 2.487971e-006, 2.722416e-006, 2.71807e-006, 
    3.198384e-006, 3.185097e-006, 3.323554e-006, 3.797039e-006, 4.10959e-006, 
    3.886321e-006, 2.813561e-006, 1.895899e-006, 1.352626e-006, 
    1.194922e-006, 8.987613e-007, 6.353839e-007, 1.856534e-006, 2.3854e-006, 
    2.379813e-006, 2.098057e-006, 1.869945e-006, 2.348521e-006, 
    2.792203e-006, 2.95686e-006, 3.353852e-006, 3.471943e-006, 2.890054e-006, 
    2.192556e-006, 1.505984e-006, 1.536034e-006, 1.389506e-006, 
    1.188093e-006, 1.193309e-006, 2.023551e-006, 3.378066e-006, 
    4.250406e-006, 4.133556e-006, 3.052974e-006, 2.639465e-006, 
    3.169203e-006, 2.512683e-006, 1.83977e-006, 2.030754e-006, 2.793817e-006, 
    3.493178e-006, 3.14747e-006, 2.744519e-006, 3.061417e-006, 3.397438e-006, 
    4.584565e-006, 6.305029e-006, 7.241568e-006, 5.284672e-006, 
    9.681771e-007, -1.081849e-006, 4.312387e-007, 1.623208e-006,
  9.186315e-007, -2.920751e-008, -7.403669e-007, -4.906487e-007, 
    6.45814e-007, 1.498905e-006, 2.052235e-006, 2.692736e-006, 2.873537e-006, 
    2.300216e-006, 1.183498e-006, 6.235859e-007, 5.925422e-007, 
    4.008152e-007, 6.292985e-007, 1.234162e-006, 1.514428e-006, 1.73484e-006, 
    1.429491e-006, 1.326052e-006, 1.533426e-006, 1.456934e-006, 
    1.638356e-006, 2.190941e-006, 2.303692e-006, 1.875656e-006, 
    1.554288e-006, 1.3679e-006, 1.565838e-006, 1.551308e-006, 1.671635e-006, 
    2.063288e-006, 2.287674e-006, 2.378075e-006, 2.659211e-006, 
    2.805739e-006, 2.667033e-006, 2.462391e-006, 2.190693e-006, 
    1.767376e-006, 1.720809e-006, 1.675112e-006, 1.641336e-006, 
    1.831326e-006, 2.070366e-006, 2.209568e-006, 2.132578e-006, 
    2.102776e-006, 1.92123e-006, 1.374482e-006, 7.399403e-007, 7.309995e-007, 
    9.512887e-007, 1.421668e-006, 1.197033e-006, 1.371749e-006, 
    1.918621e-006, 1.876401e-006, 1.764643e-006, 2.123389e-006, 
    2.575391e-006, 2.733095e-006, 2.481763e-006, 2.148224e-006, 1.80823e-006, 
    1.412355e-006, 1.262598e-006, 1.53976e-006, 1.514925e-006, 1.18983e-006, 
    8.643638e-007, 7.382014e-007, 1.036722e-006, 1.260612e-006, 
    1.338098e-006, 1.383919e-006, 2.056458e-006, 2.72763e-006, 3.117048e-006, 
    3.728616e-006, 3.788096e-006, 3.667149e-006, 3.869556e-006, 
    3.439534e-006, 2.213169e-006, 1.413597e-006, 1.944327e-006, 
    3.413085e-006, 4.920087e-006, 6.098272e-006, 6.097901e-006, 
    5.279456e-006, 4.182855e-006, 2.812942e-006, 1.42403e-006, 1.086395e-006,
  3.854905e-006, 3.152067e-006, 2.224344e-006, 1.491828e-006, 1.388016e-006, 
    1.640343e-006, 1.886087e-006, 1.79606e-006, 1.415086e-006, 1.080059e-006, 
    8.478482e-007, 8.304642e-007, 1.148976e-006, 1.462025e-006, 
    1.800779e-006, 2.273766e-006, 2.632636e-006, 2.569926e-006, 
    1.851316e-006, 9.244659e-007, 4.384401e-007, 6.008627e-007, 
    1.093967e-006, 1.753715e-006, 2.229933e-006, 2.417563e-006, 
    2.617985e-006, 3.043413e-006, 3.574018e-006, 3.720297e-006, 
    3.562842e-006, 3.434816e-006, 3.421157e-006, 3.195901e-006, 
    2.764139e-006, 2.557634e-006, 2.538883e-006, 2.447489e-006, 
    2.257996e-006, 1.959104e-006, 1.765761e-006, 1.790721e-006, 
    1.585582e-006, 1.278866e-006, 1.078818e-006, 1.061806e-006, 
    1.138919e-006, 1.265952e-006, 1.291159e-006, 1.232051e-006, 
    1.255024e-006, 1.473698e-006, 1.827477e-006, 2.178399e-006, 
    2.306798e-006, 2.306425e-006, 2.255264e-006, 2.264454e-006, 
    2.209816e-006, 2.119788e-006, 1.996606e-006, 1.824124e-006, 
    1.877023e-006, 1.994618e-006, 2.001696e-006, 2.063908e-006, 
    2.101657e-006, 1.777558e-006, 1.594025e-006, 1.60545e-006, 1.75322e-006, 
    1.874292e-006, 1.766879e-006, 1.371874e-006, 9.301784e-007, 
    7.126214e-007, 7.616713e-007, 1.099307e-006, 1.573163e-006, 1.98667e-006, 
    2.214409e-006, 2.221116e-006, 2.0803e-006, 1.845482e-006, 1.534545e-006, 
    1.237515e-006, 1.093347e-006, 1.171453e-006, 1.499528e-006, 
    1.574157e-006, 1.241364e-006, 9.476862e-007, 1.268187e-006, 
    2.214536e-006, 3.148714e-006, 3.829449e-006,
  2.924574e-006, 2.842121e-006, 2.792699e-006, 2.860374e-006, 2.927678e-006, 
    2.882726e-006, 2.709874e-006, 2.455437e-006, 2.169832e-006, 
    1.921106e-006, 1.768866e-006, 1.712738e-006, 1.692994e-006, 
    1.654996e-006, 1.575896e-006, 1.480032e-006, 1.389134e-006, 
    1.272284e-006, 1.202125e-006, 1.298983e-006, 1.496298e-006, 
    1.687406e-006, 1.893042e-006, 2.083901e-006, 2.271656e-006, 
    2.482631e-006, 2.756192e-006, 2.980082e-006, 3.050366e-006, 
    3.004297e-006, 2.867454e-006, 2.684542e-006, 2.512061e-006, 
    2.353861e-006, 2.195163e-006, 1.966306e-006, 1.658721e-006, 
    1.330771e-006, 1.076831e-006, 1.016357e-006, 1.200759e-006, 
    1.518651e-006, 1.786251e-006, 1.940974e-006, 2.011879e-006, 
    2.062046e-006, 2.09694e-006, 2.097808e-006, 2.111343e-006, 2.229311e-006, 
    2.426503e-006, 2.545216e-006, 2.548569e-006, 2.494303e-006, 
    2.435444e-006, 2.351997e-006, 2.181628e-006, 1.835051e-006, 
    1.469724e-006, 1.222614e-006, 1.169963e-006, 1.292028e-006, 
    1.405152e-006, 1.40714e-006, 1.420551e-006, 1.555655e-006, 1.748004e-006, 
    1.936876e-006, 2.007409e-006, 1.820896e-006, 1.525729e-006, 
    1.276258e-006, 1.147736e-006, 1.039703e-006, 8.620063e-007, 
    6.305413e-007, 4.674971e-007, 3.640589e-007, 3.253153e-007, 
    3.572286e-007, 4.195654e-007, 4.549561e-007, 4.367021e-007, 
    3.440664e-007, 3.243217e-007, 3.847958e-007, 3.738683e-007, 3.09421e-007, 
    2.771358e-007, 3.155064e-007, 4.663807e-007, 7.555855e-007, 
    1.201007e-006, 1.843743e-006, 2.492192e-006, 2.867329e-006,
  1.114083e-006, 1.177164e-006, 1.259618e-006, 1.365169e-006, 1.487359e-006, 
    1.611535e-006, 1.72441e-006, 1.821392e-006, 1.91142e-006, 1.997971e-006, 
    2.082783e-006, 2.172191e-006, 2.269917e-006, 2.368762e-006, 2.4573e-006, 
    2.534041e-006, 2.599109e-006, 2.646669e-006, 2.669765e-006, 
    2.658838e-006, 2.611899e-006, 2.548445e-006, 2.479031e-006, 
    2.407878e-006, 2.33362e-006, 2.259487e-006, 2.191065e-006, 2.141271e-006, 
    2.111841e-006, 2.091724e-006, 2.06813e-006, 2.042053e-006, 2.007284e-006, 
    1.96196e-006, 1.901859e-006, 1.835424e-006, 1.778179e-006, 1.743782e-006, 
    1.740926e-006, 1.768866e-006, 1.821144e-006, 1.877272e-006, 
    1.913034e-006, 1.920485e-006, 1.913158e-006, 1.895774e-006, 
    1.865351e-006, 1.823131e-006, 1.780166e-006, 1.745397e-006, 
    1.717953e-006, 1.695105e-006, 1.662447e-006, 1.618613e-006, 
    1.557766e-006, 1.49158e-006, 1.44402e-006, 1.420055e-006, 1.423034e-006, 
    1.442158e-006, 1.46662e-006, 1.488102e-006, 1.502632e-006, 1.502632e-006, 
    1.481894e-006, 1.437812e-006, 1.382305e-006, 1.31972e-006, 1.244966e-006, 
    1.162141e-006, 1.079687e-006, 9.927639e-007, 9.016185e-007, 
    8.099764e-007, 7.218105e-007, 6.345144e-007, 5.456041e-007, 
    4.560729e-007, 3.697705e-007, 2.896768e-007, 2.258503e-007, 
    1.790354e-007, 1.570565e-007, 1.630169e-007, 2.006423e-007, 
    2.710499e-007, 3.783384e-007, 5.194033e-007, 6.754935e-007, 
    8.236357e-007, 9.506675e-007, 1.032004e-006, 1.062799e-006, 
    1.065654e-006, 1.063047e-006, 1.078196e-006,
  2.326343e-007, 2.424442e-007, 2.666588e-007, 3.009316e-007, 3.353285e-007, 
    3.632681e-007, 3.827638e-007, 3.913319e-007, 3.951814e-007, 
    3.995275e-007, 4.030046e-007, 4.094619e-007, 4.180299e-007, 
    4.297026e-007, 4.41996e-007, 4.566488e-007, 4.726675e-007, 4.847127e-007, 
    4.893071e-007, 4.874445e-007, 4.871961e-007, 4.945225e-007, 
    5.092994e-007, 5.270568e-007, 5.465523e-007, 5.624471e-007, 
    5.640613e-007, 5.504019e-007, 5.295402e-007, 5.110384e-007, 
    4.946471e-007, 4.824777e-007, 4.721711e-007, 4.668316e-007, 
    4.647203e-007, 4.662104e-007, 4.685695e-007, 4.729158e-007, 
    4.763926e-007, 4.689421e-007, 4.501915e-007, 4.202648e-007, 
    3.811492e-007, 3.402954e-007, 3.02173e-007, 2.7175e-007, 2.471631e-007, 
    2.305233e-007, 2.197201e-007, 2.192232e-007, 2.425686e-007, 
    2.866509e-007, 3.468763e-007, 4.206372e-007, 4.971298e-007, 
    5.672891e-007, 6.298742e-007, 6.758196e-007, 7.056221e-007, 
    7.192814e-007, 7.150593e-007, 7.017723e-007, 6.754474e-007, 
    6.493703e-007, 6.313646e-007, 6.282603e-007, 6.335997e-007, 
    6.388152e-007, 6.430373e-007, 6.489979e-007, 6.593043e-007, 
    6.739572e-007, 6.86623e-007, 6.920868e-007, 6.896034e-007, 6.751989e-007, 
    6.604221e-007, 6.496186e-007, 6.463899e-007, 6.50612e-007, 6.568207e-007, 
    6.609187e-007, 6.599253e-007, 6.532196e-007, 6.384428e-007, 
    6.134833e-007, 5.823149e-007, 5.4767e-007, 5.063191e-007, 4.616156e-007, 
    4.131871e-007, 3.674901e-007, 3.240284e-007, 2.857822e-007, 
    2.562281e-007, 2.388432e-007,
  4.305714e-007, 3.71836e-007, 3.03291e-007, 2.657895e-007, 2.448037e-007, 
    2.403334e-007, 2.455487e-007, 2.600774e-007, 2.876445e-007, 
    3.129763e-007, 3.272566e-007, 3.438962e-007, 3.62026e-007, 3.817701e-007, 
    4.033767e-007, 4.231208e-007, 4.520538e-007, 4.839672e-007, 
    5.050771e-007, 4.931563e-007, 4.530472e-007, 4.011416e-007, 
    3.599151e-007, 3.493602e-007, 3.606602e-007, 3.481184e-007, 
    3.082578e-007, 2.567247e-007, 2.207136e-007, 2.039496e-007, 
    1.815979e-007, 1.489395e-007, 1.501813e-007, 1.670693e-007, 
    1.685595e-007, 1.294439e-007, 7.319204e-008, -7.895096e-009, 
    -9.394932e-008, -1.909309e-007, -2.490456e-007, -2.602213e-007, 
    -2.428368e-007, -2.428367e-007, -2.799654e-007, -4.011615e-007, 
    -5.666889e-007, -6.224445e-007, -5.791062e-007, -4.920589e-007, 
    -3.960708e-007, -2.695351e-007, -1.256149e-007, -2.776324e-008, 
    3.606283e-008, 8.896222e-008, 1.340386e-007, 2.043225e-007, 
    3.481186e-007, 5.535062e-007, 7.75161e-007, 9.403152e-007, 9.888672e-007, 
    9.326163e-007, 8.574889e-007, 7.556655e-007, 6.185742e-007, 
    5.069396e-007, 4.139317e-007, 3.353284e-007, 2.502675e-007, 
    1.388814e-007, 3.109631e-008, -5.694483e-008, -1.216408e-007, 
    -1.000342e-007, -3.136438e-008, 4.27417e-009, -1.509738e-008, 
    -2.366551e-008, -7.606786e-008, -1.996234e-007, -3.752086e-007, 
    -5.377556e-007, -6.246789e-007, -6.372209e-007, -6.06301e-007, 
    -5.432194e-007, -4.494661e-007, -3.409359e-007, -2.01486e-007, 
    -1.994022e-008, 1.72533e-007, 3.183161e-007, 4.075989e-007, 4.428648e-007,
  6.791727e-007, 5.816946e-007, 5.199789e-007, 3.765549e-007, 2.142564e-007, 
    1.633441e-007, 2.092893e-007, 3.071402e-007, 4.20389e-007, 5.232068e-007, 
    5.768511e-007, 5.589696e-007, 5.489115e-007, 5.332653e-007, 
    4.638507e-007, 3.655029e-007, 3.036631e-007, 2.690181e-007, 
    2.659137e-007, 2.568486e-007, 2.215828e-007, 1.66945e-007, 1.154119e-007, 
    1.637165e-007, 3.155842e-007, 4.401331e-007, 4.742815e-007, 4.69687e-007, 
    4.294538e-007, 3.52092e-007, 2.505157e-007, 1.814738e-007, 1.853232e-007, 
    2.342487e-007, 2.973301e-007, 3.050293e-007, 1.779969e-007, 
    6.673486e-008, 6.598998e-008, 8.076722e-008, -2.155457e-008, 
    -1.836045e-007, -3.498765e-007, -4.47852e-007, -4.438789e-007, 
    -3.329883e-007, -1.390258e-007, -8.14066e-008, -8.98508e-008, 
    7.058452e-008, 2.974552e-007, 4.059848e-007, 2.382226e-007, 
    -6.116625e-008, -2.614634e-007, -1.772714e-007, -3.024707e-008, 
    -2.330271e-007, -5.827073e-007, -7.486065e-007, -7.243921e-007, 
    -6.451669e-007, -5.325396e-007, -3.271525e-007, -5.197762e-008, 
    2.327588e-007, 6.653895e-007, 1.021899e-006, 1.082745e-006, 
    9.293872e-007, 8.057077e-007, 7.973877e-007, 7.978847e-007, 
    5.756092e-007, 3.597916e-007, 2.292818e-007, -6.901701e-009, 
    -3.974365e-007, -6.357309e-007, -6.492658e-007, -6.536122e-007, 
    -7.802721e-007, -9.824309e-007, -1.049486e-006, -7.63881e-007, 
    -4.066255e-007, -4.417675e-007, -5.190054e-007, -2.731358e-007, 
    1.819703e-007, 6.103783e-007, 8.398565e-007, 9.372113e-007, 
    9.928422e-007, 9.68131e-007, 8.428369e-007,
  4.6472e-007, 3.253942e-007, 2.625611e-007, 1.577563e-007, 1.488154e-007, 
    2.774623e-007, 3.917045e-007, 4.105793e-007, 4.85706e-007, 5.270566e-007, 
    4.790004e-007, 4.06233e-007, 4.156703e-007, 4.25232e-007, 3.391776e-007, 
    2.030803e-007, 1.442207e-007, 1.209998e-007, 1.360251e-007, 
    1.403714e-007, 1.655793e-007, 1.932706e-007, 2.344973e-007, 
    2.885138e-007, 3.738231e-007, 3.876066e-007, 2.955918e-007, 
    3.736986e-007, 4.478319e-007, 4.09834e-007, 2.654169e-007, 1.268363e-007, 
    6.512039e-008, 6.536879e-008, 3.941602e-008, 1.197304e-008, 
    2.128627e-008, -1.013029e-008, -7.569531e-008, -3.072844e-007, 
    -4.639949e-007, -6.709968e-007, -6.397047e-007, -3.165978e-007, 
    6.632945e-009, 7.877952e-008, 1.368953e-007, 2.580909e-007, 
    7.307067e-007, 1.004018e-006, 6.615401e-007, 3.369432e-007, 
    3.887249e-007, 3.878554e-007, 3.134737e-007, -3.15852e-007, 
    -1.243574e-006, -1.144606e-006, -3.825353e-007, -4.299709e-007, 
    -9.82307e-007, -1.431454e-006, -1.246307e-006, -6.110204e-007, 
    4.518042e-007, 2.197226e-006, 4.437744e-006, 6.347824e-006, 
    6.634299e-006, 5.331563e-006, 3.782215e-006, 3.156986e-006, 
    3.175862e-006, 3.275079e-006, 3.287247e-006, 3.030947e-006, 
    2.377782e-006, 1.5571e-006, 5.018496e-007, -1.797553e-007, 
    -8.801094e-007, -1.066871e-006, -4.698309e-007, 2.485299e-007, 
    8.242105e-007, 7.805011e-007, 2.761999e-008, -2.736319e-007, 
    -1.603839e-007, 1.326725e-007, 6.958117e-007, 1.222444e-006, 
    1.742991e-006, 2.13216e-006, 1.861579e-006, 1.062878e-006,
  5.567354e-007, 1.552721e-007, 1.859441e-007, -4.775575e-008, 
    -1.932906e-007, 2.592083e-007, 4.906724e-007, 3.268838e-007, 
    1.919047e-007, 2.176091e-007, 3.014284e-007, 5.305337e-007, 
    1.021155e-006, 1.262801e-006, 9.174671e-007, 6.251558e-007, 
    3.210481e-007, 2.222037e-007, 1.700495e-007, 1.125561e-007, 
    2.152499e-007, 5.839292e-007, 5.949814e-007, 6.522268e-007, 
    7.894409e-007, 7.038836e-007, 9.464002e-007, 1.049963e-006, 
    1.234241e-006, 1.273729e-006, 1.141109e-006, 1.068962e-006, 
    9.055459e-007, 4.473352e-007, 1.279536e-007, 5.766992e-008, 
    1.757617e-007, 1.286992e-007, 1.421099e-007, 5.183392e-008, 
    -1.343064e-007, -1.834806e-007, -1.449857e-007, 1.363983e-007, 
    3.317273e-007, -2.687893e-007, -4.323301e-007, 6.915889e-007, 
    1.56815e-006, 1.47539e-006, 1.395421e-006, 2.001402e-006, 2.308241e-006, 
    1.950986e-006, 1.254357e-006, 8.083152e-007, 9.312498e-007, 5.468e-007, 
    -4.473559e-007, 2.004717e-007, 1.531145e-006, 2.069202e-006, 
    1.635205e-006, 1.055301e-006, 1.391322e-006, 2.439868e-006, 
    3.920175e-006, 4.382484e-006, 4.869255e-006, 4.394031e-006, 
    3.530261e-006, 3.766196e-006, 3.831015e-006, 3.348218e-006, 
    3.181077e-006, 2.772909e-006, 1.716789e-006, 2.068457e-006, 
    2.311844e-006, 1.857357e-006, 8.355105e-007, 6.605469e-007, 
    7.187859e-007, 7.526855e-007, 8.367529e-007, 1.149428e-006, 
    1.165695e-006, 8.058323e-007, 8.037218e-007, 1.254233e-006, 
    2.076032e-006, 4.369817e-006, 5.167774e-006, 4.75377e-006, 3.76632e-006, 
    1.979672e-006,
  1.500599e-006, 1.027611e-006, 1.428079e-006, 1.800981e-006, 2.032074e-006, 
    2.175e-006, 1.222445e-006, 1.942915e-006, 2.588632e-006, 2.052936e-006, 
    1.963032e-006, 2.969605e-006, 3.559442e-006, 3.085585e-006, 
    2.492023e-006, 1.951112e-006, 1.459001e-006, 1.216359e-006, 1.05431e-006, 
    1.30825e-006, 1.580693e-006, 1.964647e-006, 1.457385e-006, 1.366985e-006, 
    2.202693e-006, 3.555221e-006, 3.452776e-006, 2.528531e-006, 
    2.133401e-006, 3.267876e-006, 3.302273e-006, 2.408577e-006, 
    1.637069e-006, 8.779789e-007, 7.72181e-007, 9.188325e-007, 3.072455e-008, 
    -3.213154e-007, -7.919443e-007, -8.565157e-007, -5.163965e-007, 
    -5.731463e-007, -4.471076e-007, 1.116148e-006, 3.314772e-007, 
    -1.164723e-006, -5.376323e-007, 1.897837e-006, 2.743728e-006, 
    3.101231e-006, 3.316304e-006, 2.52108e-006, 2.46371e-006, 1.694686e-006, 
    1.406846e-006, 1.535739e-006, 2.907143e-006, 2.867159e-006, 
    2.330344e-006, 2.0769e-006, 2.119492e-006, 3.045849e-006, 3.371563e-006, 
    2.876844e-006, 2.379394e-006, 2.536974e-006, 2.681764e-006, 
    2.361265e-006, 2.134394e-006, 1.623285e-006, 9.871292e-007, 
    1.504944e-006, 1.777387e-006, 2.176738e-006, 2.706722e-006, 
    3.487918e-006, 3.913221e-006, 3.480093e-006, 3.526038e-006, 
    2.928005e-006, 9.896112e-007, 8.946181e-007, 9.390733e-007, 
    4.943977e-007, 9.182113e-007, 1.091934e-006, 1.162342e-006, 
    1.845809e-006, 2.272106e-006, 1.907276e-006, 3.115512e-006, 4.52007e-006, 
    4.76271e-006, 4.087066e-006, 3.211997e-006, 2.57522e-006,
  4.281652e-006, 3.332572e-006, 3.640528e-006, 3.960158e-006, 3.602408e-006, 
    3.457492e-006, 3.88404e-006, 3.223668e-006, 2.389575e-006, 2.759746e-006, 
    3.077016e-006, 3.8823e-006, 4.835976e-006, 5.607363e-006, 4.743961e-006, 
    3.922534e-006, 3.226029e-006, 4.664737e-006, 6.569851e-006, 
    6.546255e-006, 4.809153e-006, 2.890877e-006, 3.690944e-006, 5.58513e-006, 
    5.659637e-006, 4.6928e-006, 4.88875e-006, 4.012313e-006, 4.092409e-006, 
    5.964739e-006, 4.992313e-006, 3.530385e-006, 3.831388e-006, 
    5.269104e-006, 5.354661e-006, 3.751047e-006, 2.111921e-006, 
    2.149049e-006, 1.472785e-006, 3.175701e-007, 4.165358e-007, 2.2613e-006, 
    3.246392e-006, 2.964391e-006, 2.085222e-006, 2.339038e-006, 
    4.528638e-006, 5.323741e-006, 5.219557e-006, 4.96152e-006, 4.253715e-006, 
    2.13154e-006, 2.226658e-006, 3.38684e-006, 4.185788e-006, 4.050436e-006, 
    3.475872e-006, 1.600809e-006, 1.494887e-006, 1.829296e-006, 
    1.992709e-006, 1.760995e-006, 1.253363e-006, 1.607763e-006, 
    1.508172e-006, 1.553622e-006, 2.359775e-006, 2.303896e-006, 
    2.530516e-006, 3.224291e-006, 3.689703e-006, 3.157482e-006, 
    3.752535e-006, 4.684106e-006, 5.680994e-006, 5.615184e-006, 
    4.318533e-006, 3.139478e-006, 2.311594e-006, 2.057281e-006, 
    1.781982e-006, 2.100371e-006, 2.373558e-006, 2.291726e-006, 
    2.571992e-006, 2.865792e-006, 3.463081e-006, 2.684867e-006, 2.2654e-006, 
    2.463585e-006, 2.399138e-006, 3.53709e-006, 3.654312e-006, 2.705852e-006, 
    3.228263e-006, 4.566265e-006,
  4.56589e-006, 4.638659e-006, 4.355039e-006, 5.316912e-006, 4.245766e-006, 
    2.421118e-006, 2.071064e-006, 2.149915e-006, 1.629367e-006, 
    1.722997e-006, 3.387581e-006, 5.73427e-006, 8.050157e-006, 6.927106e-006, 
    4.750045e-006, 5.417371e-006, 6.227124e-006, 7.148388e-006, 
    7.794726e-006, 7.087667e-006, 5.858196e-006, 6.229734e-006, 
    6.977896e-006, 6.204647e-006, 5.261158e-006, 4.881673e-006, 4.96487e-006, 
    3.90465e-006, 3.358897e-006, 3.629106e-006, 4.81859e-006, 3.622525e-006, 
    4.683237e-006, 4.43526e-006, 4.244775e-006, 3.628982e-006, 3.987107e-006, 
    3.116878e-006, 4.887757e-006, 4.521562e-006, 4.677404e-006, 
    5.642129e-006, 6.84155e-006, 6.178076e-006, 4.170515e-006, 5.019881e-006, 
    4.897816e-006, 4.3199e-006, 4.534104e-006, 4.075397e-006, 4.538204e-006, 
    3.627618e-006, 3.803823e-006, 5.262895e-006, 3.73627e-006, 2.19996e-006, 
    2.452662e-006, 3.173005e-006, 3.468298e-006, 3.588626e-006, 
    4.491882e-006, 6.172735e-006, 7.373768e-006, 6.16839e-006, 4.465061e-006, 
    3.29445e-006, 3.281786e-006, 4.063228e-006, 4.217456e-006, 5.36559e-006, 
    5.35963e-006, 4.808661e-006, 5.5942e-006, 6.345588e-006, 6.397122e-006, 
    6.733765e-006, 5.413895e-006, 4.810646e-006, 2.653576e-006, 
    2.559824e-006, 3.14991e-006, 3.61495e-006, 3.42136e-006, 2.65047e-006, 
    1.515252e-006, 2.023133e-006, 2.740251e-006, 3.469415e-006, 
    3.913967e-006, 3.158851e-006, 3.929241e-006, 3.805934e-006, 
    2.591487e-006, 2.303771e-006, 3.890123e-006, 4.31704e-006,
  6.958398e-006, 6.072649e-006, 3.020517e-006, 2.117877e-006, 2.080875e-006, 
    3.111911e-006, 4.676038e-006, 5.114751e-006, 5.545646e-006, 
    6.435741e-006, 7.65304e-006, 8.126774e-006, 8.224624e-006, 8.492101e-006, 
    8.237417e-006, 6.9245e-006, 7.03216e-006, 7.2897e-006, 6.625605e-006, 
    5.755252e-006, 6.792005e-006, 6.583134e-006, 8.71872e-006, 8.05984e-006, 
    6.264625e-006, 5.419604e-006, 4.960524e-006, 3.861067e-006, 
    4.222173e-006, 5.184414e-006, 4.648842e-006, 3.163943e-006, 
    3.413163e-006, 4.242786e-006, 4.903155e-006, 5.826405e-006, 
    5.942882e-006, 8.201529e-006, 7.537681e-006, 6.92934e-006, 6.627841e-006, 
    7.292185e-006, 5.577309e-006, 5.194723e-006, 5.718994e-006, 
    6.453498e-006, 7.894934e-006, 8.055245e-006, 6.965973e-006, 
    6.467408e-006, 7.117344e-006, 6.555818e-006, 5.726199e-006, 
    5.275935e-006, 5.453256e-006, 5.31803e-006, 6.733144e-006, 7.590206e-006, 
    7.049295e-006, 5.806165e-006, 4.824054e-006, 6.038128e-006, 
    7.621873e-006, 6.718368e-006, 5.81337e-006, 6.698743e-006, 8.06133e-006, 
    5.684597e-006, 6.160068e-006, 5.950955e-006, 6.011929e-006, 
    6.737861e-006, 6.937036e-006, 3.794137e-006, 2.966377e-006, 
    4.612955e-006, 4.992562e-006, 3.613461e-006, 3.171641e-006, 
    2.314453e-006, 1.304403e-006, 1.218717e-006, 1.327498e-006, 
    2.007984e-006, 1.779128e-006, 1.756278e-006, 2.703744e-006, 
    3.118617e-006, 4.297548e-006, 4.860689e-006, 4.432899e-006, 
    2.651712e-006, 3.936815e-006, 3.458486e-006, 3.56031e-006, 5.288475e-006,
  4.609232e-006, 5.148029e-006, 4.074278e-006, 3.974937e-006, 5.397624e-006, 
    6.863775e-006, 6.832855e-006, 5.808526e-006, 5.983862e-006, 
    7.433868e-006, 8.059469e-006, 7.799445e-006, 7.884255e-006, 
    6.402461e-006, 4.684603e-006, 5.506899e-006, 5.886754e-006, 6.57171e-006, 
    6.545013e-006, 7.70991e-006, 5.852482e-006, 5.703843e-006, 6.07426e-006, 
    6.240036e-006, 7.022594e-006, 8.531462e-006, 7.827755e-006, 
    7.917657e-006, 6.946471e-006, 6.218552e-006, 5.431399e-006, 
    3.047835e-006, 1.033819e-006, 2.532626e-006, 2.478611e-006, 
    3.475621e-006, 4.744952e-006, 4.060867e-006, 4.582782e-006, 
    5.853477e-006, 4.517835e-006, 1.949247e-006, 1.827804e-006, 
    3.895091e-006, 5.626727e-006, 4.522304e-006, 3.834988e-006, 
    5.783935e-006, 6.402583e-006, 5.460459e-006, 5.470021e-006, 
    6.205268e-006, 3.906394e-006, 2.4318e-006, 2.194496e-006, 4.534355e-006, 
    5.925376e-006, 3.896954e-006, 5.732281e-006, 4.404714e-006, 
    4.328716e-006, 5.612201e-006, 6.803675e-006, 5.687329e-006, 
    6.577549e-006, 6.121698e-006, 5.866639e-006, 4.840944e-006, 
    5.637658e-006, 5.824169e-006, 4.960526e-006, 5.147036e-006, 
    5.463313e-006, 4.242536e-006, 2.575967e-006, 8.96358e-007, 1.609842e-007, 
    7.441176e-007, -4.233862e-007, -2.75182e-006, -2.237481e-006, 
    -2.53267e-007, 1.629993e-006, 3.781222e-006, 3.01195e-006, 2.934959e-006, 
    3.378145e-006, 3.858213e-006, 4.02349e-006, 2.44583e-006, -7.612707e-007, 
    9.100168e-007, 2.268505e-006, 3.489657e-006, 2.874982e-006, 3.359024e-006,
  5.920527e-006, 5.116612e-006, 5.349191e-006, 5.838199e-006, 5.489386e-006, 
    3.464696e-006, 3.808293e-006, 4.08533e-006, 5.225142e-006, 6.100836e-006, 
    3.898322e-006, 3.355543e-006, -3.033128e-007, -1.86135e-006, 
    -6.245536e-007, 5.030437e-006, 6.475229e-006, 6.539303e-006, 
    7.123797e-006, 3.402733e-006, 2.161218e-006, 5.313803e-006, 
    7.010298e-006, 6.983359e-006, 4.850877e-006, 3.696165e-006, 
    5.110283e-006, 5.612823e-006, 4.830385e-006, 3.068075e-006, 
    1.828546e-006, 1.87126e-006, 3.428308e-006, 4.388936e-006, 4.306115e-006, 
    3.374791e-006, -5.9376e-007, -3.42674e-007, 1.832028e-006, 1.668115e-006, 
    8.040934e-007, 2.519468e-006, 3.065221e-006, 1.447452e-006, 
    1.506432e-006, 4.430663e-006, 5.241536e-006, 6.314296e-006, 
    5.743332e-006, 5.192363e-006, 3.457744e-006, 1.724367e-006, 
    -1.725512e-007, -2.407251e-007, 7.845993e-007, 1.647501e-006, 
    -5.875481e-007, -1.494554e-007, 1.030219e-006, 2.44347e-006, 
    3.290974e-006, 5.592583e-006, 4.747437e-006, 4.930724e-006, 1.56902e-006, 
    2.289618e-006, 1.291985e-006, -1.18372e-006, -9.897594e-007, 
    2.425961e-006, 3.219573e-006, 2.081619e-006, 1.061635e-006, 
    -6.608134e-007, -7.313465e-007, -1.982549e-006, -3.090568e-006, 
    -4.343769e-006, -3.898336e-006, -3.550275e-006, -3.347994e-006, 
    -4.41243e-006, -2.936966e-006, -8.624756e-007, -8.774259e-008, 
    -1.020802e-006, -9.404594e-007, 7.274775e-007, 1.088085e-006, 
    1.10013e-006, 1.574484e-006, 1.36177e-006, 2.50767e-006, 4.512871e-006, 
    4.437241e-006, 5.076998e-006,
  2.583041e-006, 4.336725e-007, -7.035851e-008, 9.55959e-007, 9.683772e-007, 
    6.774317e-007, -3.95079e-007, 6.126902e-008, 1.657309e-006, 
    3.130413e-006, 2.195366e-006, 1.085973e-006, 1.828179e-006, 
    2.877467e-006, 6.942377e-006, 5.469774e-006, 2.921421e-006, 2.60564e-006, 
    3.630721e-006, 3.651701e-006, 6.310194e-006, 8.376737e-006, 5.39278e-006, 
    1.744105e-006, 2.392557e-006, 4.234586e-006, 4.499208e-006, 
    1.963283e-006, -1.368378e-006, -3.498993e-006, -3.04835e-006, 
    -2.491048e-006, -1.708862e-006, -1.939456e-006, -2.236486e-006, 
    -2.117527e-006, -2.038923e-006, -6.322516e-007, -1.6993e-006, 
    -8.70672e-007, -8.525785e-008, -3.835285e-007, -3.24716e-006, 
    -3.067476e-006, -9.42322e-007, 2.399633e-006, 1.583299e-006, 
    -5.788552e-007, 1.08908e-006, 4.465928e-007, -4.4847e-007, 6.565733e-007, 
    -1.907296e-006, -6.404662e-009, -6.515002e-007, -1.681916e-006, 
    -2.178496e-006, -3.73595e-007, -2.080646e-006, 1.503082e-006, 
    5.33264e-007, 7.547987e-007, 2.72175e-006, -1.632865e-006, 
    -4.531141e-006, -4.370953e-006, -2.87277e-006, -2.789324e-006, 
    -2.856128e-006, -1.984659e-006, -3.232382e-006, -4.314703e-006, 
    -4.615085e-006, -5.789545e-006, -6.881055e-006, -9.540414e-006, 
    -1.12163e-005, -8.691171e-006, -5.735157e-006, -2.706869e-006, 
    -1.868182e-006, -1.337701e-006, -1.968267e-006, -6.075425e-007, 
    -1.665921e-007, 7.213912e-007, 8.22969e-007, 1.417149e-006, 
    -4.081157e-007, 3.345485e-008, 1.607394e-006, 4.391299e-006, 
    4.48394e-006, 3.631092e-006, 3.620786e-006, 2.672081e-006,
  -1.384764e-006, -1.899349e-006, -5.028633e-007, -6.420651e-007, 
    -2.425109e-006, -3.11851e-006, -1.89252e-006, -7.221552e-007, 
    -9.382238e-007, -1.091457e-006, 1.559209e-006, 4.093275e-006, 
    4.810146e-006, 5.238431e-006, 4.05317e-006, 4.144811e-006, 4.492624e-006, 
    2.462843e-006, -5.160837e-008, 1.664484e-007, -1.834898e-006, 
    -3.353081e-006, -4.182955e-006, -4.039532e-006, -3.977319e-006, 
    -5.515489e-006, -6.673927e-006, -8.159075e-006, -7.942886e-006, 
    -6.12718e-006, -5.077643e-006, -4.849406e-006, -3.708228e-006, 
    -3.934601e-006, -3.299439e-006, -4.24616e-006, -3.770689e-006, 
    -3.952107e-006, -4.974079e-006, -6.84877e-006, -3.64502e-006, 
    -4.19475e-006, -5.391188e-006, -3.602056e-006, -2.740893e-006, 
    -3.637073e-006, -2.686626e-006, -1.237242e-006, -1.674342e-006, 
    -1.198621e-006, 9.678824e-007, -5.591137e-007, -3.023146e-006, 
    -2.217486e-006, -3.186187e-006, -5.908878e-006, -4.893984e-006, 
    -3.84482e-006, 1.047354e-006, 1.074177e-006, 1.744729e-006, 
    4.389562e-006, 1.848044e-006, -2.457025e-006, -2.138388e-006, 
    -3.93783e-006, -5.861937e-006, -5.553859e-006, -2.646519e-006, 
    -3.488682e-006, -4.937821e-006, -7.014918e-006, -5.95557e-006, 
    -7.25706e-006, -7.893093e-006, -7.882167e-006, -1.090722e-005, 
    -1.266755e-005, -5.385106e-006, -4.355185e-006, -2.138761e-006, 
    -1.809818e-006, -1.291133e-006, -2.253128e-006, -1.018074e-006, 
    3.607624e-006, 5.448288e-006, 1.83066e-006, -1.29424e-006, 2.260433e-006, 
    4.499827e-006, 3.743222e-006, 2.71367e-006, 9.105097e-007, 
    -1.141005e-006, -1.077678e-006,
  -3.37245e-006, -2.456154e-006, -1.699922e-006, -1.719916e-006, 
    -2.513651e-006, -1.776167e-006, -2.598465e-006, -2.608771e-006, 
    -9.444348e-007, 6.039227e-007, 1.13341e-006, -1.430948e-006, 
    -4.669233e-006, -6.833005e-006, -5.893857e-006, -5.78992e-006, 
    -7.545026e-006, -8.659757e-006, -7.933453e-006, -8.517578e-006, 
    -9.156713e-006, -9.396124e-006, -7.613817e-006, -7.016781e-006, 
    -7.366089e-006, -8.111147e-006, -6.062114e-006, -6.606256e-006, 
    -5.244537e-006, -3.934848e-006, -4.999538e-006, -4.682885e-006, 
    -3.017433e-006, -3.042516e-006, -3.444228e-006, -3.155518e-006, 
    -3.952732e-006, -3.099763e-006, -4.132913e-006, -4.820973e-006, 
    -3.0491e-006, -2.515635e-006, -1.561091e-006, -4.475636e-006, 
    -2.13541e-006, -3.363513e-006, -5.420368e-006, -8.064726e-007, 
    -3.971891e-007, -1.788087e-006, -3.971978e-006, -5.538086e-006, 
    -7.662371e-006, -8.772384e-006, -1.102395e-005, -1.025914e-005, 
    -9.518686e-006, -5.170155e-006, -4.467365e-007, -4.262474e-007, 
    -3.694196e-006, -4.019412e-006, -5.834745e-006, -4.369716e-006, 
    -4.349848e-006, -5.425585e-006, -5.442969e-006, -2.878853e-006, 
    -2.719906e-006, -3.309868e-006, -3.949253e-006, -5.569133e-006, 
    -6.320401e-006, -6.476243e-006, -5.687599e-006, -5.876099e-006, 
    -7.855594e-006, -1.076331e-005, -3.377422e-006, -4.737277e-006, 
    -5.707916e-007, 2.609468e-007, 1.50991e-006, 4.003869e-006, 7.1012e-006, 
    8.433984e-006, 1.083121e-005, 1.087877e-005, 8.902753e-006, 
    6.520677e-006, 1.769691e-006, -9.580945e-007, -1.733701e-006, 
    -2.482735e-006, -1.095061e-006, -3.199475e-006,
  9.274008e-007, -3.57204e-007, -3.316218e-007, -8.331708e-007, 
    -8.134271e-007, -1.994841e-006, -2.594364e-006, -2.208581e-007, 
    -1.570315e-007, -1.092452e-006, -4.171028e-006, -4.382378e-006, 
    -4.851021e-006, -6.663127e-006, -5.730313e-006, -6.917935e-006, 
    -5.438747e-006, -3.537109e-006, -3.542449e-006, -6.294322e-006, 
    -7.752029e-006, -6.836602e-006, -5.232492e-006, -3.701026e-006, 
    -4.488799e-006, -4.46769e-006, -3.564059e-006, -2.667999e-006, 
    -2.41977e-006, -2.852774e-006, -2.477886e-006, -2.765603e-006, 
    -1.382278e-006, -9.734904e-007, -1.292499e-006, -2.34477e-006, 
    -1.443623e-006, 5.406855e-008, 5.008533e-007, 1.093921e-006, 
    3.575709e-006, 5.111269e-006, 1.734796e-006, -2.632361e-006, 
    -3.115159e-006, -1.233018e-006, 1.693197e-006, 4.901758e-007, 
    -3.337309e-006, -4.262551e-006, -6.507658e-006, -8.589723e-006, 
    -8.879426e-006, -1.01459e-005, -8.351304e-006, -1.015199e-005, 
    -8.571222e-006, -6.104347e-008, -1.391718e-006, -5.546905e-006, 
    -3.957322e-006, -4.835005e-006, -6.134509e-006, -5.719881e-006, 
    -7.115623e-006, -5.189897e-006, 1.601184e-006, -3.7384e-006, 
    -1.655468e-006, -3.298323e-006, -6.307237e-006, -4.854129e-006, 
    -5.480347e-006, -4.334448e-006, -2.758277e-006, -1.406741e-006, 
    -2.343031e-006, -3.266158e-006, -2.440012e-006, 3.308855e-006, 
    9.127632e-006, 9.444033e-006, 1.284324e-005, 1.835381e-005, 
    1.811043e-005, 1.737357e-005, 1.670016e-005, 1.240863e-005, 
    9.257772e-006, 4.46543e-006, 1.349348e-006, 1.610988e-006, 2.178596e-006, 
    -4.667254e-007, -2.04637e-006, -2.051216e-006,
  4.909211e-007, 3.723326e-007, 3.722087e-007, -3.400669e-007, 
    -9.826798e-007, -9.15252e-007, 6.13235e-007, 6.426551e-006, 
    9.546606e-006, 3.330584e-006, -2.712732e-007, -1.675853e-007, 
    1.207916e-006, 3.879446e-006, 2.326002e-006, -1.562512e-009, 
    -1.01037e-006, -2.673587e-006, -3.681779e-006, -4.19624e-006, 
    -6.829187e-007, -5.448346e-007, -6.421888e-007, -5.240972e-007, 
    -6.245555e-007, -5.904058e-007, -1.678336e-007, -4.21669e-008, 
    -9.975802e-007, -1.313113e-006, -1.450452e-006, -1.393951e-006, 
    8.829461e-007, 5.345082e-007, -2.201718e-006, -1.648264e-006, 
    5.36369e-007, 1.181714e-006, 1.531642e-006, 9.341056e-007, 
    -3.072071e-006, -5.094778e-006, -5.326865e-006, -3.251629e-006, 
    -1.358316e-006, 1.394179e-006, -2.01735e-007, -8.238567e-007, 
    -1.923936e-006, -1.366756e-006, -5.338165e-006, -7.31058e-006, 
    -5.950847e-006, -6.194359e-006, -6.049322e-006, -6.737257e-006, 
    -1.194647e-006, -2.915482e-006, -4.084359e-006, -2.499246e-006, 
    -5.050699e-006, -2.978444e-006, -8.115745e-006, -5.385853e-006, 
    -8.162682e-006, -4.815258e-006, -3.906038e-006, -4.508294e-006, 
    -5.99357e-006, -7.752032e-006, -5.635693e-006, -2.722637e-006, 
    -2.548544e-006, -1.489318e-006, -9.983255e-007, 2.034535e-007, 
    -3.117545e-007, 3.093753e-007, 1.800858e-006, 1.295835e-005, 
    1.455949e-005, 1.349752e-005, 1.907205e-005, 1.635867e-005, 
    1.447951e-005, 1.019977e-005, 6.508628e-006, 6.701048e-007, 
    -1.94852e-006, -8.966272e-007, 4.414274e-006, 3.380381e-006, 
    7.852195e-007, 7.411354e-007, 5.639358e-007, 1.119874e-006,
  -8.359029e-007, -2.110478e-007, 2.091383e-008, 1.719127e-007, 
    -4.890784e-007, 1.676806e-006, 5.51013e-006, 8.167011e-006, 
    5.845533e-006, -3.040408e-006, -1.052216e-006, 1.761865e-006, 
    2.583663e-006, 3.15227e-006, 8.865463e-007, -1.168077e-006, 
    -3.36041e-006, -1.642429e-006, -1.650874e-006, -2.980681e-006, 
    -3.999668e-006, -2.485711e-006, -1.06265e-006, -7.568024e-007, 
    6.718446e-007, 9.791811e-007, 5.402198e-007, 1.864414e-007, 
    -7.82507e-007, -4.89078e-007, -7.877227e-007, -2.208569e-007, 
    -1.442877e-006, -2.072699e-006, 1.432302e-006, 2.399759e-006, 
    1.676557e-006, -2.77234e-007, -8.643401e-007, -1.236285e-007, 
    -5.727581e-006, -6.321268e-006, -1.967274e-006, -4.509038e-006, 
    2.745717e-006, 4.927246e-006, 5.861051e-006, 5.6913e-006, 8.285346e-006, 
    6.074139e-006, 1.135399e-006, -3.757894e-006, -8.73538e-006, 
    -3.780748e-006, -3.541581e-006, -3.694318e-006, -5.977543e-006, 
    -3.864938e-006, -6.074188e-007, -9.097894e-007, -6.207403e-006, 
    -8.930463e-006, -5.936698e-006, -2.475528e-006, -5.460228e-006, 
    -3.118887e-006, -2.361037e-006, -1.344653e-006, -1.515646e-006, 
    -1.372967e-006, -2.293027e-007, -4.698322e-007, -8.904158e-007, 
    2.649199e-007, 1.673184e-007, 4.410022e-007, 4.264742e-007, 
    1.940432e-006, 1.513389e-006, 9.233678e-006, 1.284001e-005, 
    1.184797e-005, 1.351653e-005, 6.067439e-006, 1.180477e-006, 
    -7.169401e-007, 4.479552e-007, 2.79439e-006, 8.797197e-007, 
    1.347491e-006, -5.433449e-007, 1.257176e-007, 1.784093e-006, 
    1.291735e-006, 2.931092e-007, -7.094918e-007,
  -1.340577e-007, -1.874546e-007, -5.376307e-007, -2.46438e-007, 
    7.278491e-007, 5.880178e-006, 6.143433e-006, 1.222317e-006, 
    -3.424235e-006, -5.647016e-007, 1.375305e-006, 2.009847e-006, 
    8.661827e-007, -3.679661e-006, -6.826291e-006, -5.01754e-006, 
    -1.822981e-006, -5.345282e-007, -4.390455e-006, -5.966124e-006, 
    -5.980406e-006, -2.314098e-006, -3.446985e-008, 6.74826e-007, 
    3.01925e-007, 3.058976e-007, 2.192237e-007, -2.623324e-007, 
    -6.615592e-007, -1.194276e-006, -1.01658e-006, -4.674718e-007, 
    -8.161594e-007, 4.475846e-007, 9.740909e-007, 2.219084e-006, 
    -1.294648e-007, 1.859444e-007, -2.322822e-007, -3.942049e-006, 
    -4.660161e-006, -1.111327e-006, 1.216607e-006, -1.020305e-006, 
    9.468997e-006, 8.817939e-006, 8.255667e-006, 6.162176e-006, 
    4.429423e-006, -5.292964e-006, -1.988632e-006, -5.973827e-006, 
    -9.458581e-006, -1.106306e-005, -1.157293e-005, -9.022357e-006, 
    -1.160671e-005, -7.503928e-006, -4.397531e-006, -4.88244e-006, 
    -2.04103e-006, -2.442066e-007, 1.548407e-006, 2.081244e-006, 
    -1.895749e-006, 6.893551e-007, 1.020038e-006, 1.302536e-006, 
    1.678127e-007, 5.957254e-007, 5.459315e-007, -9.195974e-007, 
    3.472501e-007, 6.029286e-007, 1.582202e-008, -1.652263e-007, 
    3.334658e-007, 2.135017e-006, -9.12768e-007, 6.683913e-007, 
    8.654901e-006, 5.000642e-006, 1.179694e-005, 5.352176e-006, 
    1.412936e-006, -9.317015e-006, -7.021374e-006, -4.939062e-006, 
    -2.907291e-006, 6.586833e-007, 2.830502e-007, -3.26072e-008, 
    3.258911e-007, -2.850566e-007, -9.645501e-007, -6.90492e-007,
  -1.019932e-006, -6.973228e-007, 2.137594e-007, 1.234835e-007, 
    4.279636e-007, 7.746676e-007, 4.675541e-006, 1.606095e-007, 
    -3.198234e-006, -1.793551e-006, 3.425084e-006, 5.39067e-006, 
    5.574206e-006, -1.214948e-005, -5.828289e-006, -2.096294e-006, 
    -1.296226e-006, -4.41566e-006, -7.58017e-006, -3.702889e-006, 
    -3.25871e-006, 7.215158e-007, 9.960695e-007, 1.596834e-006, 
    4.921621e-007, -1.30442e-006, -1.160375e-006, -1.652983e-006, 
    -1.158886e-006, -4.969016e-007, -3.624185e-007, -8.128339e-008, 
    -6.340224e-008, -4.281078e-007, 3.948087e-007, 7.422541e-007, 
    -6.427081e-008, -2.294255e-007, -1.672851e-006, -3.697546e-006, 
    -2.996695e-006, 4.519288e-007, 3.464695e-006, 5.341251e-006, 
    3.87336e-006, 3.942523e-006, 3.980349e-007, -2.757661e-006, 
    -3.961919e-006, -1.147893e-005, -1.199774e-005, -8.45562e-006, 
    -1.326037e-005, -1.504602e-005, -1.480673e-005, -1.260186e-005, 
    -6.522678e-006, -3.734549e-006, 9.867654e-007, 7.323975e-006, 
    1.291539e-005, 1.053654e-005, 3.695164e-006, -2.943796e-006, 
    -6.27535e-007, 9.373334e-007, 9.853911e-007, -7.823837e-007, 
    -7.961671e-007, -1.364771e-006, -1.683406e-006, -1.320686e-006, 
    -1.141254e-006, -1.06178e-006, -2.923832e-007, -3.660189e-007, 
    6.092614e-007, 1.275592e-006, -3.538479e-006, -2.168556e-006, 
    9.923981e-006, 4.62115e-006, 6.140577e-006, 4.060246e-006, -1.67434e-006, 
    -4.935089e-006, -6.437745e-006, -3.688856e-006, -2.654217e-006, 
    -1.637088e-006, -6.444234e-007, -1.179499e-006, -9.842943e-007, 
    -1.55414e-006, -1.576118e-006, -1.637958e-006,
  -1.755304e-006, -4.027759e-007, 3.778496e-009, 3.049047e-007, 
    -5.109432e-006, -4.532632e-006, -9.096657e-007, -5.520455e-006, 
    -3.01917e-006, -5.020149e-006, -3.244676e-006, -3.696925e-006, 
    -2.893004e-006, -7.719742e-006, -1.129838e-005, -3.412064e-006, 
    -9.111758e-006, -1.232234e-005, -1.018567e-006, -1.860482e-006, 
    -2.457151e-006, -2.412074e-006, -3.742161e-007, -8.7648e-009, 
    -9.193491e-007, -1.77927e-006, -2.334587e-006, -1.410094e-006, 
    -9.878947e-007, -4.299704e-007, -1.09332e-006, 8.145253e-007, 
    2.113534e-006, 1.480707e-007, 1.070576e-006, 5.507741e-007, 
    3.564382e-007, 4.895555e-007, 1.047355e-006, -5.897864e-007, 
    7.587687e-007, -1.134551e-006, 8.172574e-007, -4.220219e-007, 
    -3.140492e-006, 3.414654e-006, -1.077547e-006, -4.142719e-006, 
    -7.132636e-006, -1.720855e-005, -1.472018e-005, -1.136618e-005, 
    -5.220922e-006, 5.813199e-007, 1.506945e-006, 1.835637e-006, 
    7.013165e-006, 1.255429e-005, 1.252138e-005, 8.327195e-006, 
    5.828642e-006, -2.070738e-007, -2.95013e-006, -1.574504e-006, 
    -8.110683e-007, -1.058676e-006, -1.852784e-006, -2.134416e-006, 
    -1.616351e-006, -2.660054e-006, -2.322418e-006, -2.856625e-006, 
    -1.817641e-006, -1.883207e-006, -6.387118e-007, -6.673954e-007, 
    2.198447e-007, -1.024649e-006, -2.153484e-005, 1.071908e-005, 
    1.714334e-005, -1.818138e-006, 3.012949e-006, 7.356386e-006, 
    -3.473777e-006, -3.495513e-006, -3.3018e-006, -1.991612e-006, 
    -1.643547e-006, -2.129448e-006, -1.86843e-006, -1.655841e-006, 
    -1.953988e-006, -2.153042e-006, -1.836144e-006, -1.845334e-006,
  -2.109083e-006, -1.408728e-006, -1.061904e-006, 1.431026e-007, 
    2.941546e-006, 2.6208e-006, -3.063615e-006, -3.636938e-006, 
    -5.383612e-006, -7.219189e-006, -5.442475e-006, -1.166383e-005, 
    -9.885751e-006, -1.315196e-005, -1.196297e-005, -9.255804e-006, 
    -1.813441e-005, -9.091273e-006, 1.767206e-006, 1.869033e-006, 
    -3.148565e-006, -3.281557e-006, 8.048373e-007, -1.280331e-006, 
    -1.036945e-006, -1.850672e-006, -1.7034e-006, -2.242105e-007, 
    -3.912282e-007, -5.041056e-007, -1.478144e-006, 2.799485e-006, 
    9.54996e-006, 6.724702e-006, 2.530389e-006, 1.077159e-006, 2.496467e-007, 
    -2.408497e-007, 7.244694e-008, -2.325647e-006, 2.561314e-006, 
    3.599176e-006, -1.537006e-006, -2.748708e-006, -3.791414e-006, 
    4.507419e-006, 9.599891e-006, 9.48416e-006, 1.613615e-005, 2.048619e-005, 
    1.023679e-005, 1.616709e-005, 2.648526e-005, 1.917066e-005, 
    1.550485e-005, 2.07498e-005, 2.57649e-005, 1.824008e-005, 1.004604e-005, 
    3.264522e-006, 3.334644e-007, -2.896487e-006, -2.202837e-006, 
    -9.873993e-007, -9.058149e-007, -1.687754e-006, -2.333595e-006, 
    -2.70215e-006, -3.517119e-006, -3.142852e-006, -3.79602e-006, 
    -2.969501e-006, -3.104232e-006, -2.524701e-006, -2.38118e-007, 
    3.481186e-007, 9.500789e-006, 2.538982e-006, -4.438254e-006, 
    1.843367e-005, 6.30624e-006, 4.489273e-006, 7.671297e-006, 8.087289e-006, 
    6.04794e-007, -4.285523e-006, -2.068105e-006, -2.434053e-006, 
    -1.425741e-006, -1.69123e-006, -1.863339e-006, -2.644284e-006, 
    -2.488566e-006, -2.974841e-006, -2.407975e-006, -2.050099e-006,
  -1.947281e-006, -1.189061e-006, -1.239104e-006, -1.534644e-006, 
    -2.214878e-006, 3.908881e-006, -7.899784e-006, 6.223658e-006, 
    -1.143977e-006, -1.964837e-005, -3.644895e-006, -1.234507e-005, 
    -7.028946e-006, -2.805209e-006, -2.558969e-006, 3.891255e-006, 
    1.09467e-005, 8.658259e-006, 3.11702e-006, 2.315821e-006, 7.752009e-006, 
    3.1534e-007, 1.252865e-006, 2.092922e-006, -1.74202e-006, 4.387666e-007, 
    2.684495e-006, 6.314542e-006, 2.281667e-006, 1.081502e-006, 
    2.168168e-006, 4.720612e-006, 5.769405e-006, 3.833997e-006, 
    3.810153e-006, -2.135284e-006, -2.261572e-006, -1.387247e-006, 
    6.636501e-007, -1.157789e-005, -7.704595e-006, -7.700495e-006, 
    -1.094484e-005, 1.311731e-005, 2.092291e-005, 2.457615e-005, 
    4.182308e-006, -5.676426e-006, 2.260534e-005, 3.743574e-005, 
    3.183215e-005, 3.415313e-005, 3.963752e-005, 3.823383e-005, 
    3.850229e-005, 3.034727e-005, 2.808465e-005, 1.810223e-005, 
    9.800919e-006, 2.814384e-006, -9.628111e-007, -1.740901e-006, 
    -1.483731e-006, -1.446229e-006, -1.655096e-006, -2.819621e-006, 
    -3.319679e-006, -4.200462e-006, -3.948507e-006, -4.488177e-006, 
    -3.761993e-006, -3.164458e-006, -3.079025e-006, -1.202595e-006, 
    2.524681e-006, 1.487402e-005, 8.982708e-006, -8.866635e-006, 
    4.50269e-006, 2.309505e-006, 1.001973e-005, 2.640918e-006, 1.183045e-005, 
    6.103814e-006, 6.593036e-007, -7.445083e-007, -2.016572e-006, 
    -1.930891e-006, -1.283311e-006, -1.760148e-006, -2.308138e-006, 
    -2.231025e-006, -2.455039e-006, -2.418902e-006, -2.28591e-006, 
    -2.187066e-006,
  -1.465973e-006, -1.17093e-006, -7.843696e-007, -2.090705e-006, 
    -4.401503e-006, 2.241199e-006, 8.071394e-006, 1.498067e-005, 
    7.957773e-006, 4.100802e-007, -3.39605e-006, -6.263403e-006, 
    -4.040889e-006, -5.416077e-007, 1.524593e-005, 1.854874e-005, 
    1.039707e-005, 1.020836e-005, 1.499336e-005, 1.807939e-005, 1.5765e-005, 
    1.23381e-005, 1.110107e-005, 5.342117e-006, -3.985388e-006, 
    1.413184e-006, 1.642113e-005, 1.649837e-005, 9.439809e-006, 5.61965e-006, 
    4.086449e-006, 4.1237e-006, 5.139336e-006, 2.751676e-006, 2.362358e-007, 
    -3.667628e-007, -4.024754e-006, -1.196954e-005, 1.892011e-006, 
    -3.206427e-006, -2.264635e-005, -3.161162e-005, -2.034895e-005, 
    1.083346e-005, 2.135478e-005, 2.840973e-005, 2.455979e-005, 
    2.926519e-005, 5.260426e-005, 6.671764e-005, 5.764657e-005, 
    4.981937e-005, 4.86239e-005, 5.334224e-005, 4.853153e-005, 3.770695e-005, 
    3.110002e-005, 2.238296e-005, 1.577082e-005, 8.617894e-006, 
    5.710548e-006, 2.415032e-006, 1.29223e-006, -4.895755e-007, 
    -1.915741e-006, -2.557484e-006, -3.214624e-006, -3.380151e-006, 
    -3.388967e-006, -2.843587e-006, -2.108587e-006, -1.607535e-006, 
    -6.624282e-007, 7.499521e-007, 3.336421e-006, 8.672789e-006, 
    3.693458e-007, 8.466643e-006, -8.222392e-006, -3.465451e-006, 
    -4.583788e-006, -1.410811e-005, -8.626845e-006, -3.910633e-006, 
    -5.05097e-007, 2.207134e-007, -9.50145e-007, 6.470109e-007, 
    2.121977e-006, 1.440747e-006, 7.179151e-007, -1.786384e-007, 
    -2.042028e-006, -1.639323e-006, -1.919465e-006, -1.739286e-006,
  5.940772e-006, 7.918778e-006, 5.09687e-006, 3.820584e-006, -7.271214e-006, 
    -6.706032e-007, -1.208801e-005, -2.529903e-005, 1.485898e-005, 
    1.505149e-005, 1.340054e-005, -1.74711e-006, -3.989851e-006, 
    1.104119e-006, 1.026136e-005, 1.060544e-005, -2.693354e-005, 
    -2.003976e-005, -2.738278e-006, 7.580282e-006, 1.976063e-005, 
    1.482884e-005, 1.49478e-006, -4.850757e-006, -3.193752e-006, 
    1.095837e-005, 2.546143e-005, 1.063279e-005, 1.843291e-005, 
    1.740858e-005, 2.553617e-006, 9.398336e-006, 6.805163e-006, 
    5.354166e-006, 6.033537e-006, -1.907665e-006, -7.641633e-006, 
    4.179725e-006, 1.548883e-005, 4.149922e-006, 5.918264e-008, 
    -7.284361e-006, -6.178823e-006, 1.482225e-005, 2.743732e-005, 
    3.316409e-005, 5.878811e-005, 7.170929e-005, 7.235674e-005, 
    6.691657e-005, 4.592706e-005, 3.347055e-005, 2.474939e-005, 
    1.627423e-005, 1.155913e-005, 8.105537e-006, 5.271337e-006, 
    3.994433e-006, 3.352193e-006, 1.765343e-006, 1.522578e-006, 
    1.038538e-006, 6.841387e-007, 8.799652e-007, 1.896692e-007, 
    -2.049628e-007, -1.278495e-007, -7.445351e-008, -7.274593e-009, 
    8.574891e-007, 1.181714e-006, 2.21362e-006, 3.221062e-006, 5.912831e-006, 
    3.426081e-006, -8.957431e-007, 1.029606e-006, -2.048218e-006, 
    -1.790331e-005, -5.110302e-006, -9.411509e-006, -1.090661e-005, 
    -3.296456e-006, -1.6392e-006, -1.196884e-006, -5.818583e-008, 
    -1.308272e-007, 3.851381e-006, 7.227487e-006, 7.662975e-006, 
    5.601896e-006, 4.534103e-006, 3.6789e-006, 2.848409e-006, 1.726104e-006, 
    3.419497e-006,
  -3.255722e-006, 6.18404e-006, 1.791341e-007, -8.82415e-006, 2.212888e-006, 
    -2.697154e-006, -2.491899e-006, 1.096571e-005, 3.568213e-005, 
    2.66093e-005, 1.667346e-005, 5.59581e-006, 6.478575e-006, 1.670277e-005, 
    3.246672e-005, 3.983432e-005, -2.743007e-006, 1.402192e-005, 
    1.797023e-005, 1.072616e-005, 1.755748e-005, 3.989844e-006, 
    -1.132458e-005, 2.153829e-007, 3.119501e-006, 1.114613e-005, 
    7.836947e-005, 8.755364e-006, 1.669558e-005, 3.188147e-005, 
    1.941391e-005, 3.890697e-005, -3.471025e-006, -8.322619e-006, 
    -4.719746e-006, -1.974957e-006, -9.917523e-006, -6.18217e-006, 
    4.085596e-006, 9.472104e-006, 8.906485e-006, 1.958168e-005, 
    1.405644e-005, 2.238035e-005, 4.026535e-005, 3.890251e-005, 
    6.809227e-005, 8.788684e-005, 7.545891e-005, 5.442568e-005, 
    5.168188e-005, 4.179372e-005, 3.306784e-005, 2.444007e-005, 
    1.701929e-005, 1.202392e-005, 7.616904e-006, 5.258547e-006, 3.95569e-006, 
    3.683744e-006, 3.171517e-006, 3.627615e-006, 3.571861e-006, 
    3.641895e-006, 2.536354e-006, 2.314948e-006, 1.060394e-006, 
    1.543812e-006, 2.409569e-006, 1.874493e-006, 5.187272e-006, 
    4.272586e-006, 8.501907e-006, 8.9405e-006, 1.078565e-005, -1.34603e-005, 
    -3.544421e-005, -4.090936e-006, -5.274334e-006, -1.589316e-005, 
    -6.761599e-006, -1.67459e-006, -2.926039e-006, -3.299438e-006, 
    -3.94627e-006, -2.90505e-006, -2.380661e-006, 6.308655e-007, 
    2.750185e-006, 1.839724e-006, 3.72087e-006, 9.251688e-006, 4.691559e-006, 
    4.436379e-006, 4.529506e-006, 2.267989e-007,
  3.659032e-006, 1.352125e-005, -3.167937e-006, -9.028188e-006, 
    -1.925799e-006, 5.096865e-006, 1.576436e-005, 1.215009e-005, 
    1.626181e-005, 1.260134e-005, 3.949223e-005, 1.277891e-005, 
    8.007437e-006, 1.109348e-005, 2.218082e-005, 4.012269e-005, 
    5.236211e-005, 3.25432e-005, 3.406264e-005, 2.590164e-005, 6.413284e-006, 
    1.187878e-005, 3.318928e-006, -1.215644e-005, -9.000622e-006, 
    -1.962926e-006, 1.525943e-006, -9.532709e-006, 1.846798e-006, 
    2.186302e-006, -7.293565e-007, -4.37296e-007, 3.185414e-008, 
    1.632288e-007, -5.844908e-006, -6.922019e-006, -6.545262e-006, 
    -3.002766e-006, 4.709582e-006, 5.989343e-006, 1.737989e-005, 
    1.268563e-005, 4.385074e-007, 2.348192e-005, 1.188694e-005, 
    4.853093e-006, 1.557684e-005, 1.735307e-005, 2.37319e-005, 3.110425e-005, 
    4.677814e-005, 4.996388e-005, 5.779458e-005, 5.763092e-005, 
    5.556524e-005, 5.225136e-005, 4.5464e-005, 3.572671e-005, 3.056806e-005, 
    2.838888e-005, 1.885078e-005, 2.106571e-005, 1.788108e-005, 
    1.350548e-005, 6.994913e-006, 5.052061e-007, 1.371216e-006, 
    -5.063979e-006, 4.314432e-006, 4.723101e-006, 3.345111e-006, 
    4.148424e-006, 4.314817e-006, -7.913193e-006, -2.172731e-005, 
    -3.091612e-005, -2.199741e-005, -6.637298e-006, -9.712279e-006, 
    -1.298085e-005, -2.28442e-006, -1.592136e-006, -5.182697e-006, 
    -6.331946e-006, -1.07988e-005, -1.224285e-005, -1.47465e-005, 
    -1.432988e-005, -1.368232e-005, -1.341758e-005, -5.563179e-006, 
    -3.887912e-006, -6.0487e-006, 1.449684e-006, 1.040153e-006, 5.645728e-006,
  -1.109463e-006, -1.321929e-006, -2.347253e-006, -7.258827e-007, 
    -9.508904e-007, -9.919922e-007, 1.244672e-006, 3.060502e-006, 
    2.612599e-006, 6.809014e-006, 2.157061e-005, 3.659032e-006, 
    5.683728e-006, 2.646377e-006, 9.170239e-006, 2.467936e-005, 
    3.077666e-005, 2.743061e-005, 1.831198e-005, 1.491686e-005, 
    8.730516e-006, 3.340519e-006, 1.012224e-006, -1.543295e-005, 
    -1.059542e-005, -5.394912e-006, -3.640796e-006, -2.526567e-006, 
    -9.274208e-007, -1.561823e-005, -3.528303e-005, -1.898016e-005, 
    -1.104367e-006, 1.44404e-005, -1.374538e-005, -1.891124e-005, 
    -1.053566e-006, 2.211227e-005, 2.712911e-005, 1.417206e-005, 
    1.372999e-005, 9.493218e-006, 1.947166e-005, 2.071452e-005, 
    1.457129e-005, 7.258292e-006, -2.640045e-006, -1.09575e-005, 
    -2.149436e-005, -2.811383e-005, -1.752009e-005, -1.915363e-005, 
    -1.143881e-005, -9.133597e-006, -2.784026e-005, -2.75148e-005, 
    -2.547807e-005, -2.396808e-005, -2.310244e-005, -1.3727e-005, 
    -1.219465e-006, 5.565038e-006, 2.728098e-006, -1.043016e-006, 
    -5.32846e-006, -9.949195e-006, -5.128546e-006, 7.078706e-007, 
    7.307346e-006, 4.889254e-006, 5.316055e-006, 1.086934e-005, 8.34516e-007, 
    -1.166532e-005, -1.645056e-005, -1.687564e-005, -1.585466e-005, 
    -1.191715e-005, -3.058907e-006, -3.431065e-006, -1.112218e-005, 
    -9.111015e-006, -1.07376e-005, -2.03378e-005, -2.348877e-005, 
    -2.128464e-005, -2.290589e-005, -1.300121e-005, -1.206231e-005, 
    -5.076403e-006, -2.776282e-006, -2.355118e-007, 1.660534e-006, 
    6.89728e-007, -9.009718e-007, -1.336705e-006,
  2.372288e-007, 5.870335e-007, 4.010174e-007, 1.227383e-007, 2.333794e-007, 
    5.940831e-008, 2.28785e-007, 9.388253e-007, 4.012659e-007, 2.161466e-006, 
    3.287745e-006, 1.271121e-006, 4.177467e-006, 3.122218e-006, 
    1.267671e-005, 1.565173e-005, 8.871331e-006, 1.867444e-005, 
    1.323987e-005, 1.115519e-005, 1.804581e-006, -5.692684e-006, 
    -8.604122e-006, -9.883013e-006, -1.459191e-005, -1.086413e-005, 
    -4.642654e-006, -1.30169e-006, -5.80519e-006, -1.022562e-005, 
    -7.973555e-006, -1.064881e-005, -5.201808e-006, 1.683489e-005, 
    -4.464819e-006, -2.832763e-006, 1.337535e-005, 2.70171e-005, 
    2.35819e-005, 1.501736e-006, -1.693828e-006, 5.872484e-006, 
    2.936082e-006, 1.158273e-005, 2.766086e-006, 3.792287e-006, 
    4.880436e-006, 3.828281e-006, -5.40186e-006, -8.151495e-006, 
    -1.135675e-005, -1.179595e-005, -6.781993e-007, -7.305978e-006, 
    -2.156664e-005, -1.867047e-005, -7.588977e-006, -1.396009e-005, 
    -8.917552e-006, -4.25112e-006, -5.37392e-006, 1.927525e-006, 
    -6.582646e-006, -4.414913e-006, -5.533358e-006, 7.962859e-006, 
    1.236305e-005, 1.203784e-005, 1.499808e-005, 1.133512e-005, 
    1.545305e-005, 1.101996e-005, -1.592882e-006, -1.324584e-005, 
    -1.64738e-005, -1.35122e-005, -1.203996e-005, -9.39227e-006, 
    -9.799938e-006, -1.079335e-005, -1.347842e-005, -8.995408e-006, 
    -1.486659e-005, -1.330209e-005, -8.64759e-006, -6.404718e-006, 
    -5.197972e-006, -3.160361e-006, -1.562459e-006, -8.57759e-007, 
    9.616742e-007, -2.218521e-007, 1.282021e-007, 1.542276e-009, 
    2.907491e-007, 7.058429e-008,
  1.931462e-007, 3.784173e-007, 7.025177e-007, 8.409742e-007, 2.926116e-007, 
    1.741474e-007, -2.579864e-007, 2.775862e-007, 4.360353e-007, 
    5.402193e-007, 2.499598e-006, 2.180465e-006, 5.519566e-006, 
    4.021379e-006, 6.115985e-006, 4.330081e-006, 2.432418e-006, 
    4.334923e-006, 1.314772e-005, 1.217977e-005, 2.045485e-006, 
    -2.862835e-006, -7.207927e-007, 1.203942e-006, -1.009859e-005, 
    -3.974088e-006, 7.421299e-007, 8.896518e-007, -6.911141e-007, 
    -3.627018e-006, 5.20255e-006, 4.478235e-006, -9.029922e-006, 
    -6.334791e-006, -5.608723e-006, -1.983281e-006, 5.077018e-007, 
    9.573574e-006, 3.276291e-007, -1.056673e-005, -1.393996e-005, 
    -3.188914e-006, 6.275186e-007, 1.788321e-006, 2.742359e-006, 
    -4.85847e-006, -9.290328e-006, -8.855215e-006, -1.052452e-005, 
    -1.424211e-005, -1.052178e-005, -8.524155e-006, 5.617767e-008, 
    -2.578217e-006, -6.123824e-006, -4.292477e-006, -5.835755e-007, 
    3.801219e-006, 8.878291e-006, 4.071044e-007, -9.688956e-007, 
    -1.358436e-006, -1.228695e-005, -8.781206e-006, -2.484092e-006, 
    6.527011e-006, 1.832736e-005, 1.735854e-005, 1.140875e-005, 2.34773e-006, 
    4.639751e-007, -9.782098e-007, -5.398266e-006, -8.918043e-006, 
    -3.531273e-006, -5.690454e-006, -9.809999e-006, -1.254846e-005, 
    -1.486523e-005, -1.335909e-005, -1.032558e-005, -1.355219e-005, 
    -1.271263e-005, -7.873848e-006, -8.898924e-006, -6.183187e-006, 
    -3.73393e-006, -3.348364e-006, -2.518864e-006, -1.931138e-006, 
    -1.070597e-006, 1.900421e-007, 2.793247e-007, 2.724951e-007, 
    4.633541e-007, 1.866891e-007,
  1.919045e-007, 2.525979e-008, 2.666587e-007, 4.149253e-007, 4.94274e-007, 
    2.317651e-007, -1.324439e-007, -1.525607e-007, 2.954677e-007, 
    1.398747e-007, 8.374255e-006, 1.855992e-006, 7.120791e-007, 
    9.579485e-007, 2.274093e-006, 2.421119e-006, 3.271851e-006, 
    9.898613e-007, 6.195458e-006, 6.477338e-006, 2.270493e-006, 
    2.199341e-006, -2.736546e-006, -4.571871e-006, -4.818859e-006, 
    -4.911743e-006, 3.65009e-006, 1.958809e-006, 2.153767e-006, 
    1.986375e-006, 3.86488e-007, 1.601555e-006, 7.272061e-006, 2.379769e-006, 
    4.476366e-006, -9.326817e-006, -1.092633e-005, 4.828158e-006, 
    3.460846e-006, -3.927893e-006, -2.581321e-006, 7.509479e-007, 
    3.095894e-006, 1.005508e-006, 2.472403e-006, -1.05222e-006, 
    -5.813634e-006, -4.116764e-006, -5.744096e-006, -7.187151e-006, 
    -7.660883e-006, -8.153736e-006, -6.48493e-006, -3.956082e-006, 
    -3.785835e-006, 1.957444e-006, 3.941781e-006, 6.991924e-006, 
    5.847265e-006, 1.269013e-006, -2.562201e-006, -5.813139e-006, 
    -4.632222e-006, -1.626782e-006, -5.000531e-006, -1.173665e-006, 
    1.084337e-005, 1.139621e-005, 3.567021e-006, 1.796107e-007, 
    1.904424e-006, -3.175384e-006, -3.285159e-006, 4.236572e-006, 
    4.346228e-006, 4.932466e-006, -2.711702e-006, -5.022259e-006, 
    -6.324746e-006, -8.657276e-006, -8.353167e-006, -9.041476e-006, 
    -1.054923e-005, -1.142777e-005, -7.277428e-006, -3.761998e-006, 
    -3.477136e-006, -2.392206e-006, -2.667753e-006, -2.81043e-006, 
    -1.478515e-006, 3.30831e-008, -2.205138e-008, 1.248495e-007, 
    5.493803e-008, 1.495605e-007,
  -3.444131e-007, -2.484247e-007, -5.797272e-007, -7.805482e-008, 
    1.198823e-007, 1.037394e-007, 3.755335e-008, -4.750737e-008, 
    -3.459309e-008, 4.103308e-007, 4.035013e-007, 8.851812e-007, 
    1.556479e-006, -9.757257e-007, -1.401434e-007, 7.248696e-007, 
    5.568245e-006, -1.419161e-006, 1.508024e-007, 2.120239e-006, 
    3.675299e-006, 4.775874e-006, 8.291772e-007, -6.093901e-006, 
    -2.896982e-006, -2.661916e-006, -4.251124e-006, 1.317811e-006, 
    2.552e-006, 9.328651e-007, 1.452418e-006, 5.937372e-007, 6.124183e-006, 
    4.535596e-006, 3.593959e-008, 3.65519e-006, 1.737029e-006, 2.753288e-006, 
    1.592489e-006, 2.748529e-007, -1.429464e-006, -2.23015e-006, 
    7.718118e-007, -2.154777e-006, 3.445697e-006, 8.368752e-007, 
    -1.768341e-006, -3.221829e-006, -3.785339e-006, -1.113809e-006, 
    -4.466199e-006, -4.797625e-006, -4.252242e-006, -2.513276e-006, 
    -1.679557e-006, 1.52444e-006, 1.158245e-006, 4.455249e-006, 
    6.717219e-007, 1.5309e-006, -1.193408e-006, -5.317429e-006, 
    -5.143209e-006, -6.934733e-007, 2.214583e-007, -4.411563e-006, 
    -9.758496e-007, 4.011196e-006, 3.2983e-006, 3.025238e-006, 2.923616e-007, 
    2.485442e-006, 4.890113e-006, 7.637769e-006, 7.683961e-006, 
    8.217798e-006, 5.077625e-006, 4.166668e-006, -4.117137e-007, 
    -1.598342e-006, 8.265706e-007, 7.811213e-007, -2.051846e-006, 
    -5.099624e-006, -3.303287e-006, -2.644036e-006, -1.92369e-006, 
    -5.046013e-007, -7.463723e-007, -1.096673e-006, -1.830059e-006, 
    -1.084628e-006, -2.630776e-007, -2.661818e-007, -6.441747e-007, 
    -5.583687e-007,
  -4.195399e-007, -1.356727e-007, -7.647499e-007, -8.551502e-007, 
    -8.63346e-007, -3.598109e-007, -2.416232e-008, 3.032369e-009, 
    -1.391494e-007, -2.220993e-007, 4.778823e-007, 8.266942e-007, 
    3.747198e-006, 3.013315e-006, -2.477017e-006, -2.375069e-006, 
    2.711567e-006, 9.790574e-007, 1.10373e-006, 1.114535e-006, 1.476013e-006, 
    2.534864e-006, 3.250988e-006, -9.208397e-007, 1.42607e-007, 
    -1.559107e-006, -5.84696e-007, 1.355284e-007, 3.606146e-008, 
    1.965265e-006, 1.975699e-006, 1.281987e-007, -1.530607e-007, 
    -3.476012e-006, -7.080052e-007, 7.879462e-007, -1.752574e-006, 
    2.512606e-007, 4.654299e-006, 7.683208e-006, 5.786296e-006, 
    8.623465e-008, -2.553716e-007, 8.243369e-007, 2.356421e-006, 
    3.210756e-006, -1.674589e-006, -4.126454e-006, -3.090077e-006, 
    6.40679e-007, -3.902811e-006, 1.177723e-007, -5.614729e-007, 
    -1.024775e-006, 2.046945e-007, 1.123228e-006, 1.185192e-006, 
    2.153396e-006, 1.443106e-006, 3.553196e-007, -2.875872e-006, 
    -3.672339e-006, -2.932992e-006, -1.394945e-006, 3.432342e-008, 
    -4.913356e-006, -3.787574e-006, -1.437911e-009, 3.998654e-006, 
    7.360607e-006, 3.97717e-006, 6.601149e-006, 9.243115e-006, 5.424446e-006, 
    6.237926e-006, 5.03987e-006, 4.588986e-006, 5.50193e-006, 4.478592e-006, 
    -1.045082e-007, -1.375949e-006, 1.023018e-006, 1.370587e-006, 
    -8.408679e-007, 6.71349e-007, 1.139619e-006, 1.60168e-006, 3.056502e-007, 
    -1.047538e-007, 2.168626e-007, -1.653605e-006, -2.238972e-006, 
    -1.850051e-006, -8.023754e-007, -9.157484e-007, -5.838249e-007,
  -1.472804e-006, -1.347882e-006, -1.346268e-006, -1.649134e-006, 
    -1.917852e-006, -3.055927e-006, -2.380284e-006, -8.006368e-007, 
    -1.540106e-006, -2.556862e-006, -9.337539e-007, -6.580824e-007, 
    1.879585e-006, 2.451666e-006, 3.285386e-006, 3.651084e-006, 
    2.248512e-006, 4.744052e-007, 2.603256e-007, 1.224183e-006, 
    -2.689376e-008, 6.918381e-007, 2.306379e-006, 1.302662e-006, 
    6.622845e-007, 2.526276e-007, 2.008107e-006, 3.550378e-006, 
    6.291284e-007, -2.198614e-006, 1.363882e-006, 3.377523e-006, 
    5.264257e-006, 1.867284e-006, -1.933251e-006, 4.64348e-007, 
    -4.570255e-006, -5.689828e-006, -5.902795e-006, -7.562037e-006, 
    -2.379784e-006, 2.972589e-006, 2.306009e-006, -3.35693e-006, 
    -1.949265e-006, 2.745717e-006, 1.830413e-006, -7.266281e-007, 
    -3.496883e-006, -3.572379e-006, -2.13541e-006, 7.184099e-007, 
    -9.717951e-008, 4.975671e-006, 7.650431e-006, 3.303019e-006, 
    6.524351e-008, -3.887453e-007, 1.800981e-006, 1.596213e-006, 
    -2.472299e-006, -3.835258e-006, -3.151916e-006, -1.980188e-006, 
    1.627011e-006, 2.662637e-008, -5.135508e-006, -5.283655e-006, 
    -2.559844e-006, 2.559077e-006, 5.071292e-006, 3.451907e-006, 
    2.56243e-006, 2.073923e-006, 7.570306e-007, 5.232225e-006, 8.070398e-006, 
    6.655282e-006, 3.47264e-006, -1.904191e-006, -2.977697e-006, 
    -1.791686e-006, -3.138666e-007, -1.014469e-006, -1.595363e-006, 
    2.727955e-006, 3.247884e-006, 9.060441e-007, 5.46057e-007, 
    -1.458275e-006, -4.250381e-006, -3.83501e-006, -7.564149e-006, 
    -7.032178e-006, -5.455137e-006, -4.294959e-006,
  -4.779123e-006, -4.799736e-006, -3.693822e-006, -5.736025e-006, 
    -5.593844e-006, -3.994453e-006, -5.217093e-006, -5.005745e-006, 
    -1.12543e-005, -1.098657e-005, -2.184705e-006, -7.990225e-007, 
    2.891497e-006, 2.809167e-006, 3.815247e-006, 2.106579e-006, 
    1.900446e-006, 1.613847e-006, 4.376489e-007, 1.164703e-006, 
    2.195489e-006, 1.379153e-006, 1.121736e-006, 8.546344e-007, 
    1.002529e-006, 1.002403e-006, 1.843947e-006, 5.249978e-006, 
    5.110405e-006, -6.912342e-007, -3.310033e-007, 2.197194e-007, 
    -1.495153e-006, -6.718637e-007, -1.183473e-006, -1.45939e-006, 
    -2.468114e-007, -1.735807e-006, 2.402372e-006, -3.250374e-006, 
    -7.064329e-006, -7.074639e-006, -5.331087e-006, -4.163208e-006, 
    -5.580798e-006, -4.750684e-006, -6.947812e-008, 4.199825e-006, 
    5.7832e-006, 1.30602e-006, -1.706998e-006, 1.340166e-006, -2.084493e-006, 
    1.374305e-006, 5.536331e-006, 8.299874e-006, 4.646354e-006, 
    -2.723755e-006, -4.795111e-007, 1.412558e-006, -1.537996e-006, 
    -1.717555e-006, -2.461869e-006, -5.950978e-006, -1.837014e-006, 
    1.649486e-006, 1.249728e-007, -3.702019e-006, -5.797618e-006, 
    -5.203933e-006, 1.983626e-007, 4.838212e-006, 3.485558e-006, 
    5.173482e-006, 2.767694e-006, -1.754934e-006, 1.641543e-006, 
    9.681458e-006, 4.907753e-006, 1.130928e-006, -1.584805e-006, 
    -1.279957e-006, -2.181605e-006, -4.862231e-007, -1.137152e-006, 
    -6.149035e-006, -2.326393e-006, 1.485323e-006, 3.003131e-006, 
    -2.255487e-006, -3.838986e-006, -5.882805e-006, -1.036247e-005, 
    -1.214775e-005, -1.441148e-005, -7.521432e-006,
  -3.191529e-006, -2.212273e-006, -1.440019e-006, -1.38364e-006, 
    -3.979556e-006, 2.66078e-006, 1.170165e-006, -1.105118e-006, 
    -5.833255e-006, -1.230234e-005, -7.271717e-006, -2.655336e-006, 
    2.13191e-006, 1.384373e-006, 1.021652e-006, 1.681896e-006, 1.107332e-006, 
    3.168252e-007, 2.158704e-007, -2.006182e-007, 1.252618e-006, 
    1.270997e-006, 7.464762e-007, 1.422864e-006, 1.863194e-006, 
    2.222436e-006, 2.187294e-006, 3.408692e-006, 4.605752e-006, 
    3.039267e-006, 1.136388e-006, 1.402872e-006, 2.78756e-006, 2.397772e-006, 
    3.962397e-006, 5.127667e-006, 4.611213e-006, 4.588244e-006, 
    5.636866e-007, -2.804842e-006, -4.915961e-006, -2.063622e-006, 
    -2.499983e-006, -1.458466e-007, 2.584668e-006, 3.475638e-006, 
    -7.082344e-007, -4.064226e-006, 1.849803e-006, 3.042631e-006, 
    4.738751e-006, 7.176204e-006, 9.146512e-006, 8.87581e-006, 9.563497e-006, 
    6.757116e-006, 5.962636e-006, 2.120367e-006, 8.826973e-007, 
    1.485703e-006, -2.566194e-007, 1.984641e-006, -5.872971e-007, 
    -9.29158e-007, 1.935223e-007, 1.511762e-007, 3.841946e-006, 
    1.929129e-006, -1.999188e-006, -3.53649e-006, 3.848745e-007, 
    4.750915e-006, 2.45055e-006, 4.460097e-006, 9.882875e-006, 6.634051e-006, 
    2.857098e-006, 2.207908e-006, 3.74161e-006, 3.796667e-007, 
    -3.545552e-006, -4.747209e-006, -5.446691e-006, -2.372337e-006, 
    -7.725721e-007, -2.497753e-006, -1.00776e-005, -5.033686e-006, 
    -6.600712e-007, -3.24033e-006, -5.073793e-006, -4.875981e-006, 
    -6.601042e-006, -8.602764e-006, -1.013026e-005, -6.323755e-006,
  -2.257349e-006, -2.316581e-006, -3.606152e-006, -4.174382e-006, 
    -6.162354e-007, -2.699668e-006, -2.983157e-006, 1.467941e-006, 
    2.341396e-006, -1.776911e-006, 1.201297e-007, -1.458026e-006, 
    6.408009e-007, 1.258702e-006, 1.984637e-006, 1.694189e-006, 
    2.334444e-006, 2.275707e-006, 1.789434e-006, 1.662773e-006, 
    2.582671e-006, 1.825817e-006, 1.661532e-006, 1.010599e-006, 
    8.607186e-007, 9.581971e-007, 1.016187e-006, 8.383665e-007, 
    1.382135e-006, 2.00848e-006, 2.076032e-006, 2.157492e-006, 2.993696e-006, 
    4.026967e-006, 4.435134e-006, 4.790402e-006, 4.444322e-006, 
    2.706229e-006, 1.94068e-006, 1.007867e-006, 2.373527e-007, 
    -2.058292e-006, -1.807581e-006, -1.401273e-006, 2.455767e-006, 
    4.485795e-006, 8.213945e-006, 7.17261e-006, 4.941161e-006, 7.380608e-006, 
    7.650444e-006, 8.90599e-006, 8.891213e-006, 6.537572e-006, 3.382243e-006, 
    3.388574e-006, 2.544555e-006, 6.792507e-006, 3.563182e-006, 
    3.909663e-007, 4.927861e-007, -4.587782e-007, 2.902056e-006, 
    8.599141e-006, 1.038493e-005, 7.432503e-006, 6.310322e-006, 
    7.185145e-006, 5.657528e-006, 1.445463e-006, 1.255226e-006, 
    7.564253e-006, 1.229649e-005, 8.868479e-006, 1.164469e-005, 8.62695e-006, 
    9.057228e-006, 6.701477e-006, 7.968822e-006, 8.101313e-006, 
    4.047459e-006, 3.638423e-006, 2.142468e-006, -1.818138e-006, 
    -2.637702e-006, -1.9176e-006, -2.018805e-006, -8.88911e-006, 
    -6.010203e-006, -3.16868e-006, -3.117268e-006, -4.966754e-006, 
    -8.484052e-006, -1.074282e-005, -8.743948e-006, -7.086441e-006,
  3.859948e-006, 3.494499e-006, 3.564284e-006, 3.452526e-006, 5.576316e-006, 
    4.711925e-006, 3.612216e-006, 5.292696e-006, 2.891252e-006, 
    3.589991e-006, 4.330329e-006, 5.106433e-006, 3.017537e-006, 
    2.585775e-006, 2.157615e-006, 2.22256e-006, 1.366861e-006, 3.683867e-006, 
    3.392052e-006, 3.038274e-006, 3.933089e-006, 2.909752e-006, 
    2.066842e-006, 1.424107e-006, 1.103732e-006, 7.999961e-007, 
    1.336934e-006, 6.896034e-007, 5.501533e-007, 8.196159e-007, 
    1.134899e-006, 1.221078e-006, 1.398153e-006, 1.99122e-006, 2.638924e-006, 
    3.215599e-006, 4.203173e-006, 4.232478e-006, 1.535618e-006, 6.21174e-007, 
    -4.332032e-007, 2.463639e-008, 9.219402e-007, -6.90241e-007, 
    -1.416673e-006, 2.139739e-006, 7.107657e-006, 5.957911e-006, 
    1.080116e-005, 1.083122e-005, 1.103002e-005, 1.208713e-005, 1.18435e-005, 
    9.935655e-006, 7.644972e-006, 6.247246e-006, 6.068178e-006, 
    7.135975e-006, 9.807627e-006, 9.673153e-006, 4.197464e-006, 
    -7.304698e-007, -2.447705e-006, 2.344757e-006, 8.12926e-006, 
    8.711144e-006, 4.640275e-006, 3.641153e-006, 3.391927e-006, 
    5.610959e-006, 5.515719e-006, 3.692187e-006, 4.736139e-006, 
    8.642603e-006, 1.350547e-005, 1.180637e-005, 7.003848e-006, 
    8.229221e-006, 9.929445e-006, 6.774368e-006, 6.546252e-006, 
    2.943903e-006, 5.542537e-006, 5.718372e-006, 4.263027e-006, 
    -2.655208e-006, -3.470053e-006, 7.236304e-007, 1.486693e-006, 
    -1.566925e-006, -1.615354e-006, -2.335219e-007, 2.078148e-006, 
    1.784589e-006, 3.651454e-006, 5.179078e-006,
  7.904371e-006, 8.839919e-006, 1.004641e-005, 6.683596e-006, 5.716387e-006, 
    5.791515e-006, 6.560537e-006, 6.262639e-006, 4.839203e-006, 
    4.505544e-006, 4.762961e-006, 5.397503e-006, 4.16443e-006, 4.138476e-006, 
    2.35431e-006, 1.710703e-006, 2.562679e-006, 3.147176e-006, 3.017909e-006, 
    3.232858e-006, 2.730691e-006, 2.509407e-006, 3.289979e-006, 
    3.457369e-006, 2.617689e-006, 1.688851e-006, 1.424728e-006, 
    1.526552e-006, 1.29335e-006, 1.51935e-006, 1.206301e-006, 1.293969e-006, 
    1.548779e-006, 1.676558e-006, 1.995939e-006, 2.579692e-006, 
    3.493133e-006, 3.10297e-006, 2.465075e-006, 1.142351e-006, 3.580179e-006, 
    3.472396e-006, 7.82984e-007, -4.390313e-007, 1.223685e-006, 
    3.518715e-006, 4.200814e-006, 4.001889e-006, 7.495095e-006, 
    1.406762e-005, 1.194781e-005, 1.093217e-005, 1.325104e-005, 
    1.492307e-005, 1.128135e-005, 8.723069e-006, 7.706567e-006, 7.22153e-006, 
    9.386178e-006, 7.054394e-006, 6.481692e-006, 7.13698e-006, 4.112168e-006, 
    5.996917e-006, 4.716774e-006, 3.970837e-006, 1.499729e-006, 
    1.055302e-006, 6.437813e-007, 8.465613e-007, 1.471419e-006, 
    1.446086e-006, 2.869147e-006, 3.769301e-006, 7.093869e-006, 
    7.482544e-006, 4.292451e-006, 2.711811e-006, 4.283756e-006, 
    3.726589e-006, 5.945862e-006, 6.339749e-006, 2.236342e-006, 
    6.043098e-006, 7.693277e-006, 6.788898e-006, 3.81151e-007, 7.628842e-009, 
    2.312958e-006, 2.329976e-006, 2.99442e-007, 3.437628e-006, 5.298785e-006, 
    5.552352e-006, 7.08456e-006, 6.712529e-006,
  5.485164e-006, 6.266115e-006, 6.577797e-006, 4.30239e-006, 4.768053e-006, 
    6.107543e-006, 6.622626e-006, 6.468274e-006, 5.106804e-006, 
    3.400248e-006, 3.652949e-006, 4.82952e-006, 4.979896e-006, 3.676417e-006, 
    3.507536e-006, 3.946129e-006, 2.868773e-006, 1.969364e-006, 1.69779e-006, 
    1.9526e-006, 2.741368e-006, 2.397275e-006, 2.570006e-006, 1.455024e-006, 
    9.949517e-007, 1.429942e-006, 1.933353e-006, 2.191267e-006, 
    2.832389e-006, 2.238704e-006, 2.26776e-006, 2.435398e-006, 1.564178e-006, 
    1.323151e-006, 1.76969e-006, 1.948131e-006, 2.38548e-006, 1.700646e-006, 
    2.444589e-006, 1.491775e-006, 9.809191e-007, 2.090314e-006, 
    7.344315e-007, -7.463677e-007, -1.004035e-006, 4.139329e-007, 
    4.200687e-006, 5.952937e-006, 7.168379e-006, 6.359864e-006, 
    9.441053e-006, 9.338855e-006, 9.314888e-006, 1.087144e-005, 
    8.370902e-006, 7.636027e-006, 5.360249e-006, 5.045091e-006, 
    7.190243e-006, 1.010974e-005, 8.352654e-006, 1.412338e-005, 
    1.396828e-005, 1.06971e-005, 7.253195e-006, 3.548888e-006, 3.27781e-006, 
    3.190638e-006, 1.894735e-006, 1.552007e-006, 1.322529e-006, 
    1.449191e-006, 2.009474e-006, 5.964703e-007, 1.859595e-006, 4.73092e-006, 
    8.086043e-006, 5.069051e-006, 2.169163e-006, 4.571975e-006, 
    3.183435e-006, 7.677081e-007, -1.859e-006, 2.18779e-006, 3.980153e-006, 
    3.748934e-006, 8.926254e-007, -3.713649e-007, 1.9978e-006, 8.671777e-007, 
    1.469307e-006, 2.833262e-006, 6.111513e-006, 7.503655e-006, 
    1.028235e-005, 7.948704e-006,
  1.235523e-005, 1.174118e-005, 9.107887e-006, 5.241291e-006, 3.234099e-006, 
    5.345224e-006, 6.400226e-006, 7.607346e-006, 9.506246e-006, 
    8.032275e-006, 5.440716e-006, 3.374794e-006, 3.957181e-006, 
    3.349338e-006, 2.94713e-006, 2.706847e-006, 2.219827e-006, 1.419263e-006, 
    1.503206e-006, 1.750939e-006, 1.511154e-006, 5.746151e-007, 
    8.800889e-007, 1.351463e-006, 2.210018e-006, 3.219696e-006, 
    3.126812e-006, 3.151025e-006, 2.096397e-006, 3.45116e-006, 4.883039e-006, 
    2.92962e-006, 2.45949e-006, 2.644635e-006, 4.181814e-006, 2.833507e-006, 
    1.463099e-006, 5.251941e-007, -7.098652e-007, -1.239227e-006, 
    -1.467464e-006, 1.492279e-006, 2.591488e-006, 2.672949e-006, 
    1.938897e-007, 7.761555e-007, 5.128535e-006, 5.198697e-006, 
    4.747439e-006, 7.47075e-006, 8.185387e-006, 8.111125e-006, 5.737616e-006, 
    4.127553e-006, 4.998023e-006, 9.229338e-006, 1.128371e-005, 
    1.066978e-005, 8.967076e-006, 9.066163e-006, 1.107608e-005, 
    1.576474e-005, 1.145744e-005, 7.288334e-006, 4.912967e-006, 
    3.830643e-006, 3.941781e-006, 3.681136e-006, 2.948124e-006, 
    2.647367e-006, 2.054548e-006, 1.183825e-006, 3.359395e-006, 
    3.506297e-006, 1.794773e-006, 2.561934e-006, 6.619026e-006, 
    8.052642e-006, 3.870629e-006, 5.962229e-007, -4.299691e-007, 
    -9.335054e-007, 5.238271e-007, 3.933337e-006, 3.191133e-006, 
    2.497611e-006, 1.155888e-006, -8.37892e-007, -1.48837e-007, 
    -1.76251e-006, -1.000313e-006, 2.770179e-006, 7.617651e-006, 
    9.268573e-006, 1.169846e-005, 1.118362e-005,
  9.133222e-006, 7.571212e-006, 7.075992e-006, 6.924249e-006, 7.245246e-006, 
    8.257897e-006, 5.777481e-006, 4.876086e-006, 7.544017e-006, 
    7.207496e-006, 5.684846e-006, 5.935433e-006, 6.359744e-006, 
    5.978645e-006, 3.41242e-006, 2.49314e-006, 3.318912e-006, 3.534235e-006, 
    3.135876e-006, 2.300169e-006, 1.054433e-006, 1.628499e-006, 
    2.598069e-006, 2.58031e-006, 2.765459e-006, 2.499224e-006, 2.233984e-006, 
    2.494879e-006, 2.486062e-006, 2.972336e-006, 2.623028e-006, 
    2.238703e-006, 2.579071e-006, 2.706847e-006, 3.057646e-006, 
    2.932477e-006, 1.513141e-006, 9.322439e-007, 4.542894e-007, 
    5.905104e-007, 2.618153e-007, 1.36537e-006, 2.832762e-006, 2.508289e-006, 
    2.166184e-006, 2.245659e-006, 2.165192e-006, 2.160101e-006, 
    1.886416e-006, 4.146923e-006, 7.386683e-006, 6.526512e-006, 6.50143e-006, 
    6.330813e-006, 6.895192e-006, 7.495089e-006, 1.11008e-005, 1.049121e-005, 
    5.656657e-006, 7.192593e-006, 1.025007e-005, 9.798927e-006, 6.34149e-006, 
    3.503068e-006, 2.227899e-006, 2.201202e-006, 2.950357e-006, 
    3.408816e-006, 2.959298e-006, 3.023993e-006, 2.189281e-006, 
    1.392193e-006, 1.441614e-006, 3.90341e-006, 4.627111e-006, 6.019502e-006, 
    7.154969e-006, 6.269841e-006, 4.238937e-006, 1.791421e-006, 
    2.294055e-007, 4.402591e-007, 2.581432e-006, 6.167395e-006, 
    8.597894e-006, 1.003797e-005, 9.767762e-006, 5.009701e-006, 
    6.688642e-007, -1.091332e-006, 5.563634e-007, 2.81004e-006, 
    2.736771e-006, 3.116013e-006, 4.440972e-006, 7.304603e-006,
  -5.617185e-007, -2.233428e-007, 6.442788e-007, 1.113418e-006, 
    1.817747e-006, 2.505436e-006, 2.752051e-006, 3.4606e-006, 6.220913e-006, 
    7.579527e-006, 7.319258e-006, 6.435493e-006, 5.163554e-006, 
    5.248988e-006, 5.410044e-006, 5.442082e-006, 5.254451e-006, 
    4.196964e-006, 2.878459e-006, 2.353813e-006, 2.338664e-006, 
    2.314202e-006, 3.311834e-006, 3.990707e-006, 3.813011e-006, 
    3.437997e-006, 4.134378e-006, 4.263397e-006, 2.918692e-006, 
    1.971227e-006, 1.945524e-006, 2.752049e-006, 3.32922e-006, 2.89932e-006, 
    2.433163e-006, 2.141225e-006, 1.863567e-006, 1.880206e-006, 
    2.396407e-006, 2.23386e-006, 1.650232e-006, 1.535243e-006, 2.216723e-006, 
    2.290855e-006, 2.943154e-006, 3.254837e-006, 2.959795e-006, 
    4.104453e-006, 4.413902e-006, 5.702233e-006, 5.737994e-006, 
    6.331557e-006, 6.526884e-006, 7.119827e-006, 5.748795e-006, 
    4.583649e-006, 4.469034e-006, 4.561048e-006, 4.527024e-006, 
    4.767679e-006, 4.452767e-006, 3.607498e-006, 1.46794e-006, 1.20481e-006, 
    2.137002e-006, 1.099012e-006, 1.836619e-006, 3.289731e-006, 
    3.628733e-006, 2.952096e-006, 2.721128e-006, 3.942154e-006, 
    5.267861e-006, 4.591347e-006, 4.155365e-006, 4.514111e-006, 
    5.324857e-006, 6.812738e-006, 5.86391e-006, 4.478847e-006, 2.258449e-006, 
    2.28465e-006, 3.923404e-006, 3.181698e-006, 2.91122e-007, -1.432491e-007, 
    2.167675e-006, 1.565291e-006, 2.113036e-006, 1.111679e-006, 
    -6.017035e-007, -3.015739e-007, 5.626935e-007, -5.151578e-007, 
    2.587094e-007, 2.095028e-006,
  -5.119242e-006, -5.793396e-006, -3.338799e-006, -3.385758e-007, 
    1.262804e-006, 2.325874e-006, 2.85524e-006, 2.644141e-006, 3.205418e-006, 
    3.141342e-006, 2.09851e-006, 9.802989e-007, 1.092058e-006, 2.4539e-006, 
    4.055651e-006, 4.379006e-006, 3.769424e-006, 3.978289e-006, 
    3.355668e-006, 2.592853e-006, 3.124576e-006, 4.357026e-006, 
    4.937178e-006, 4.896451e-006, 4.676162e-006, 4.778482e-006, 
    4.450408e-006, 3.739622e-006, 3.09316e-006, 2.53623e-006, 2.445953e-006, 
    2.447817e-006, 2.598815e-006, 2.452162e-006, 2.39914e-006, 2.232122e-006, 
    2.616821e-006, 3.478107e-006, 3.198463e-006, 3.345114e-006, 
    2.874487e-006, 2.742735e-006, 2.735905e-006, 2.739507e-006, 
    2.436392e-006, 1.984019e-006, 2.238827e-006, 3.750177e-006, 
    6.255189e-006, 8.711027e-006, 8.462671e-006, 6.347324e-006, 
    4.401978e-006, 4.01281e-006, 4.444819e-006, 4.364477e-006, 3.682625e-006, 
    3.705473e-006, 3.53287e-006, 2.67692e-006, 1.715175e-006, 1.071693e-006, 
    7.158051e-007, 7.009044e-007, 1.14558e-006, 1.459621e-006, 2.012205e-006, 
    2.773406e-006, 3.391556e-006, 3.679893e-006, 4.353674e-006, 4.7606e-006, 
    4.190133e-006, 3.226153e-006, 2.673568e-006, 2.055791e-006, 
    2.000159e-006, 2.796502e-006, 3.640777e-006, 3.45526e-006, 3.569127e-006, 
    4.63543e-006, 5.938039e-006, 4.671939e-006, 2.14942e-006, 1.140452e-007, 
    -5.296843e-007, -1.077426e-006, 1.243516e-007, 1.325263e-006, 
    1.181963e-006, 1.210024e-006, 2.284027e-006, 2.410439e-006, 
    5.775983e-007, -1.915241e-006,
  1.694279e-007, -1.263688e-006, -1.392211e-006, -1.307275e-006, 
    -1.006396e-006, 1.089575e-007, 9.283958e-007, 2.270493e-006, 
    3.291845e-006, 3.604518e-006, 3.852996e-006, 3.252107e-006, 
    2.612973e-006, 2.473146e-006, 2.375544e-006, 2.454769e-006, 
    2.885039e-006, 3.688087e-006, 3.855974e-006, 3.39913e-006, 2.11378e-006, 
    1.803837e-006, 2.063613e-006, 2.197724e-006, 2.445332e-006, 
    2.870387e-006, 3.576703e-006, 3.71752e-006, 3.057771e-006, 1.752926e-006, 
    1.388219e-006, 1.421623e-006, 1.858724e-006, 2.531636e-006, 
    2.839469e-006, 2.583293e-006, 1.869651e-006, 1.737279e-006, 
    1.304152e-006, 1.402251e-006, 1.535244e-006, 2.288002e-006, 
    2.642649e-006, 2.437014e-006, 2.377036e-006, 2.551877e-006, 
    2.644139e-006, 2.301164e-006, 2.135139e-006, 2.936326e-006, 3.64202e-006, 
    3.643012e-006, 2.597076e-006, 1.965392e-006, 1.772918e-006, 
    1.848418e-006, 1.892624e-006, 1.576223e-006, 1.57374e-006, 1.880579e-006, 
    2.159107e-006, 1.596961e-006, 1.076786e-006, 1.038416e-006, 
    1.705243e-006, 2.455639e-006, 2.565039e-006, 2.332828e-006, 
    2.668849e-006, 3.339651e-006, 3.720002e-006, 3.43154e-006, 2.680522e-006, 
    2.248265e-006, 2.917947e-006, 3.125198e-006, 2.855611e-006, 
    2.541321e-006, 2.67779e-006, 2.832016e-006, 2.231252e-006, 2.520832e-006, 
    3.790037e-006, 4.411789e-006, 2.947378e-006, 1.367482e-006, 
    1.193387e-006, 1.445838e-006, 1.261807e-006, 1.346496e-006, 
    1.351837e-006, 5.580841e-008, 6.239152e-007, 2.303399e-006, 2.68077e-006, 
    1.956203e-006,
  -4.697085e-007, -1.371725e-006, -1.715322e-006, -1.069855e-006, 
    2.488559e-008, 1.176249e-006, 2.022884e-006, 2.088449e-006, 
    2.243794e-006, 2.549638e-006, 2.184188e-006, 1.191647e-006, 5.41957e-007, 
    7.479657e-007, 1.512395e-006, 2.368095e-006, 3.023497e-006, 
    3.558946e-006, 3.468917e-006, 2.907392e-006, 2.403236e-006, 
    2.111049e-006, 1.952229e-006, 2.124584e-006, 2.341768e-006, 
    2.388584e-006, 2.494382e-006, 2.480474e-006, 1.941053e-006, 
    1.266029e-006, 1.025872e-006, 7.502015e-007, 8.086877e-007, 
    1.401009e-006, 1.854874e-006, 2.156747e-006, 2.375794e-006, 
    2.294831e-006, 1.904544e-006, 1.565792e-006, 1.276957e-006, 
    1.310982e-006, 1.560452e-006, 1.756899e-006, 1.843326e-006, 
    1.696674e-006, 1.540708e-006, 1.333334e-006, 1.412559e-006, 
    1.341654e-006, 1.42895e-006, 1.926276e-006, 2.470666e-006, 2.507049e-006, 
    2.2243e-006, 1.961666e-006, 1.454034e-006, 1.026865e-006, 9.655223e-007, 
    1.172772e-006, 1.299557e-006, 1.593979e-006, 1.826314e-006, 2.03195e-006, 
    2.360272e-006, 2.598939e-006, 2.626506e-006, 2.336803e-006, 
    2.034558e-006, 1.958935e-006, 2.219332e-006, 2.472776e-006, 
    2.318425e-006, 1.635579e-006, 1.307258e-006, 1.35047e-006, 2.002769e-006, 
    2.839467e-006, 2.867283e-006, 2.694306e-006, 2.634701e-006, 
    2.593102e-006, 2.509532e-006, 1.877723e-006, 1.242188e-006, 
    1.226666e-006, 1.021775e-006, 1.096281e-006, 1.551015e-006, 
    1.892873e-006, 1.718031e-006, 1.574856e-006, 1.961044e-006, 
    2.221941e-006, 1.340411e-006, 3.358236e-007,
  -1.136163e-006, -3.645318e-007, 1.236067e-007, 3.216674e-007, 
    3.604109e-007, 3.041587e-007, 2.544884e-007, 3.970436e-007, 7.71186e-007, 
    1.040277e-006, 1.181217e-006, 1.240697e-006, 1.238711e-006, 
    1.143715e-006, 1.143964e-006, 1.298439e-006, 1.41293e-006, 1.444348e-006, 
    1.407343e-006, 1.346621e-006, 1.361149e-006, 1.355811e-006, 
    1.321289e-006, 1.430315e-006, 1.477254e-006, 1.575478e-006, 
    1.777761e-006, 1.639801e-006, 1.317191e-006, 1.101248e-006, 
    1.063623e-006, 1.125462e-006, 1.226542e-006, 1.115156e-006, 
    8.392358e-007, 6.414227e-007, 6.067776e-007, 7.638605e-007, 1.03531e-006, 
    1.363757e-006, 1.628128e-006, 1.849411e-006, 1.970359e-006, 
    2.022761e-006, 1.900447e-006, 1.562935e-006, 1.313837e-006, 
    1.227783e-006, 1.379154e-006, 1.755533e-006, 2.098509e-006, 
    2.276453e-006, 2.236965e-006, 1.981161e-006, 1.672707e-006, 
    1.470051e-006, 1.521212e-006, 1.698536e-006, 1.965391e-006, 
    2.098508e-006, 2.008729e-006, 1.962038e-006, 2.119742e-006, 
    2.221567e-006, 2.133278e-006, 1.953222e-006, 1.634709e-006, 
    1.406722e-006, 1.274599e-006, 1.051329e-006, 9.245455e-007, 
    9.362184e-007, 9.512437e-007, 9.421788e-007, 1.07691e-006, 1.346248e-006, 
    1.734672e-006, 2.179844e-006, 2.560195e-006, 2.720757e-006, 
    2.495004e-006, 1.969489e-006, 1.492403e-006, 1.143592e-006, 
    7.967672e-007, 6.254043e-007, 6.477558e-007, 8.751222e-007, 
    1.309243e-006, 1.557472e-006, 1.297571e-006, 6.630289e-007, 
    8.523693e-008, -4.785243e-007, -1.119772e-006, -1.50062e-006,
  1.966228e-007, 2.313918e-007, 2.446805e-007, 3.158329e-007, 4.874446e-007, 
    6.74454e-007, 8.417201e-007, 1.013829e-006, 1.112424e-006, 1.051702e-006, 
    8.178777e-007, 5.102934e-007, 3.483674e-007, 2.982006e-007, 
    2.790771e-007, 2.660386e-007, 3.58426e-007, 6.182026e-007, 9.925939e-007, 
    1.379155e-006, 1.664388e-006, 1.845189e-006, 1.905166e-006, 
    1.894984e-006, 1.917212e-006, 1.983645e-006, 2.005377e-006, 
    1.961915e-006, 1.875612e-006, 1.782604e-006, 1.762115e-006, 
    1.774408e-006, 1.720392e-006, 1.583052e-006, 1.438014e-006, 
    1.351711e-006, 1.362639e-006, 1.465581e-006, 1.592738e-006, 
    1.658055e-006, 1.629494e-006, 1.631108e-006, 1.722378e-006, 
    1.862573e-006, 2.001526e-006, 2.093044e-006, 2.06883e-006, 2.030459e-006, 
    2.076902e-006, 2.193628e-006, 2.317804e-006, 2.322771e-006, 
    2.158734e-006, 1.916217e-006, 1.697046e-006, 1.571752e-006, 
    1.540211e-006, 1.561942e-006, 1.626141e-006, 1.741128e-006, 
    1.895107e-006, 2.057654e-006, 2.141598e-006, 2.198595e-006, 
    2.213744e-006, 2.126199e-006, 1.835627e-006, 1.392194e-006, 
    9.451583e-007, 6.630294e-007, 5.803281e-007, 6.186988e-007, 
    7.148114e-007, 8.612155e-007, 9.888686e-007, 1.047852e-006, 
    1.042637e-006, 9.33486e-007, 7.371623e-007, 5.434474e-007, 4.256046e-007, 
    4.00521e-007, 4.08344e-007, 3.789137e-007, 3.385564e-007, 3.160803e-007, 
    2.995653e-007, 2.474117e-007, 1.789904e-007, 1.623507e-007, 
    1.176477e-007, 1.867875e-008, -7.308699e-008, -8.910592e-008, 
    9.860742e-009, 1.181425e-007,
  8.578622e-007, 9.606806e-007, 1.055427e-006, 1.148683e-006, 1.234862e-006, 
    1.296702e-006, 1.320916e-006, 1.303531e-006, 1.242933e-006, 
    1.155016e-006, 1.052199e-006, 9.49753e-007, 8.450725e-007, 7.511958e-007, 
    6.843889e-007, 6.537166e-007, 6.533442e-007, 6.765654e-007, 
    7.139429e-007, 7.639856e-007, 8.261977e-007, 8.971024e-007, 
    9.657715e-007, 1.028729e-006, 1.070701e-006, 1.093549e-006, 
    1.099882e-006, 1.100379e-006, 1.097026e-006, 1.093922e-006, 
    1.088707e-006, 1.081256e-006, 1.065362e-006, 1.043879e-006, 
    1.015442e-006, 9.827836e-007, 9.45779e-007, 9.147348e-007, 8.896513e-007, 
    8.737566e-007, 8.636989e-007, 8.541374e-007, 8.535167e-007, 
    8.777311e-007, 9.220621e-007, 9.862608e-007, 1.068217e-006, 
    1.165447e-006, 1.263174e-006, 1.364005e-006, 1.460862e-006, 
    1.550393e-006, 1.62552e-006, 1.687484e-006, 1.741004e-006, 1.782976e-006, 
    1.813523e-006, 1.84494e-006, 1.869527e-006, 1.873749e-006, 1.848169e-006, 
    1.794525e-006, 1.73343e-006, 1.667244e-006, 1.597953e-006, 1.52382e-006, 
    1.453163e-006, 1.399519e-006, 1.365619e-006, 1.349725e-006, 
    1.345627e-006, 1.341032e-006, 1.327745e-006, 1.294218e-006, 
    1.240822e-006, 1.16433e-006, 1.073929e-006, 9.668893e-007, 8.530196e-007, 
    7.406406e-007, 6.261498e-007, 5.081824e-007, 3.956789e-007, 
    2.939782e-007, 2.023362e-007, 1.301892e-007, 9.032783e-008, 
    9.318546e-008, 1.303138e-007, 1.864419e-007, 2.609472e-007, 
    3.512237e-007, 4.570215e-007, 5.603365e-007, 6.550831e-007, 7.52189e-007,
  -1.197122e-010, -3.240564e-008, -5.748916e-008, -6.642972e-008, 
    -5.475715e-008, -2.892841e-008, 3.853984e-009, 3.688479e-008, 
    7.016422e-008, 1.012083e-007, 1.295205e-007, 1.491403e-007, 
    1.603163e-007, 1.652834e-007, 1.682635e-007, 1.662767e-007, 
    1.615579e-007, 1.538592e-007, 1.536107e-007, 1.625514e-007, 
    1.781976e-007, 1.990592e-007, 2.224044e-007, 2.447562e-007, 
    2.594087e-007, 2.683495e-007, 2.730681e-007, 2.758001e-007, 
    2.730684e-007, 2.653695e-007, 2.522067e-007, 2.395408e-007, 
    2.291099e-007, 2.273714e-007, 2.358156e-007, 2.589122e-007, 
    2.944266e-007, 3.411169e-007, 3.942646e-007, 4.469155e-007, 
    4.968342e-007, 5.470015e-007, 5.971688e-007, 6.530479e-007, 7.15881e-007, 
    7.826884e-007, 8.395614e-007, 8.735856e-007, 8.740822e-007, 
    8.408038e-007, 7.861663e-007, 7.141448e-007, 6.441092e-007, 
    5.782949e-007, 5.104948e-007, 4.506423e-007, 4.15127e-007, 4.049448e-007, 
    4.21584e-007, 4.687708e-007, 5.54701e-007, 6.657142e-007, 7.898905e-007, 
    9.05871e-007, 9.982584e-007, 1.057615e-006, 1.087914e-006, 1.102815e-006, 
    1.109272e-006, 1.120448e-006, 1.139074e-006, 1.159936e-006, 
    1.177569e-006, 1.188993e-006, 1.189242e-006, 1.17136e-006, 1.132866e-006, 
    1.076987e-006, 1.015395e-006, 9.470974e-007, 8.758201e-007, 
    8.028046e-007, 7.34756e-007, 6.699361e-007, 6.08096e-007, 5.460078e-007, 
    4.859066e-007, 4.287854e-007, 3.741479e-007, 3.214971e-007, 2.70088e-007, 
    2.176856e-007, 1.68015e-007, 1.180962e-007, 7.51312e-008, 3.638809e-008,
  -2.593999e-007, -6.419475e-008, 9.574433e-008, 2.077513e-007, 
    2.710815e-007, 2.849891e-007, 2.604022e-007, 2.084965e-007, 
    1.357294e-007, 7.090944e-008, 3.067635e-008, 2.446745e-008, 
    3.663672e-008, 5.575987e-008, 7.264782e-008, 8.158861e-008, 8.58106e-008, 
    9.673806e-008, 1.2207e-007, 1.456634e-007, 1.424349e-007, 1.086589e-007, 
    7.388962e-008, 7.860831e-008, 1.126326e-007, 1.498854e-007, 
    1.613098e-007, 1.424351e-007, 1.223184e-007, 1.091556e-007, 
    6.470043e-008, 1.031117e-008, -6.046935e-008, -1.098914e-007, 
    -1.220607e-007, -1.409355e-007, -1.74463e-007, -2.114676e-007, 
    -1.988017e-007, -1.640325e-007, -1.198257e-007, -9.797054e-008, 
    -1.307531e-007, -1.826588e-007, -2.484722e-007, -3.018681e-007, 
    -3.113059e-007, -3.023647e-007, -3.058415e-007, -3.023642e-007, 
    -1.975591e-007, 2.869001e-008, 2.949241e-007, 4.796984e-007, 
    5.018012e-007, 4.404581e-007, 3.74893e-007, 3.133014e-007, 3.036159e-007, 
    3.825921e-007, 5.348331e-007, 7.007322e-007, 8.179547e-007, 
    8.847612e-007, 8.802906e-007, 8.124905e-007, 7.876547e-007, 
    8.400575e-007, 8.879897e-007, 9.163018e-007, 9.319483e-007, 
    9.135701e-007, 8.812844e-007, 8.030536e-007, 6.42121e-007, 4.225769e-007, 
    2.42273e-007, 1.513756e-007, 1.700021e-007, 2.450045e-007, 2.750551e-007, 
    2.532e-007, 2.032809e-007, 1.824193e-007, 1.81426e-007, 1.849029e-007, 
    1.228145e-007, -8.31551e-009, -1.394455e-007, -2.715692e-007, 
    -4.568406e-007, -6.652083e-007, -7.809408e-007, -7.593342e-007, 
    -6.428567e-007, -4.667747e-007,
  1.861449e-007, 1.238083e-007, -2.768672e-008, -1.14362e-007, 
    -1.019441e-007, -7.09e-008, -3.5634e-008, 4.806088e-008, 2.022878e-007, 
    3.609852e-007, 4.372296e-007, 4.03702e-007, 3.406202e-007, 2.877212e-007, 
    2.673561e-007, 2.703364e-007, 2.705847e-007, 2.750551e-007, 
    2.621408e-007, 2.455012e-007, 2.382989e-007, 1.923537e-007, 
    1.749689e-007, 2.055162e-007, 2.291098e-007, 1.96824e-007, 2.221561e-007, 
    2.042747e-007, 9.201926e-008, 1.875503e-008, -5.177708e-008, 
    -1.193288e-007, -1.146101e-007, -2.818342e-008, 6.569371e-008, 
    1.697535e-007, 2.708332e-007, 2.519582e-007, 1.317557e-007, 
    1.106458e-007, 1.252986e-007, 3.81267e-008, -1.563335e-007, 
    -2.380415e-007, -3.861396e-008, 2.944269e-007, 4.724959e-007, 
    2.586648e-007, 5.79962e-008, 3.390642e-008, 2.427705e-007, 8.184525e-007, 
    1.46864e-006, 1.703333e-006, 1.578163e-006, 1.404812e-006, 1.314413e-006, 
    1.277408e-006, 1.356384e-006, 1.451006e-006, 1.65093e-006, 1.756728e-006, 
    1.796465e-006, 1.742325e-006, 1.456967e-006, 1.14156e-006, 8.333532e-007, 
    5.768043e-007, 4.667836e-007, 4.968349e-007, 7.101694e-007, 
    9.798803e-007, 9.264847e-007, 7.230838e-007, 9.04133e-007, 1.482298e-006, 
    1.983473e-006, 1.983473e-006, 1.54687e-006, 1.170367e-006, 1.049419e-006, 
    9.436208e-007, 6.376501e-007, 1.498856e-007, -3.177624e-007, 
    -6.666983e-007, -8.231602e-007, -1.060089e-006, -1.40058e-006, 
    -1.627574e-006, -1.424422e-006, -8.191864e-007, -1.461506e-007, 
    2.57422e-007, 2.442598e-007, 1.662772e-007,
  5.119839e-007, 5.477465e-007, 4.248118e-007, 2.549386e-007, 6.047844e-008, 
    -2.346474e-008, -6.079972e-009, 7.330982e-009, 5.253128e-008, 
    2.000527e-007, 3.493127e-007, 2.864795e-007, 1.695053e-007, 
    1.004631e-007, -2.743832e-008, -1.061661e-007, -1.651074e-008, 
    7.513131e-008, 1.332458e-007, 2.03033e-007, 2.703364e-007, 2.708332e-007, 
    1.911123e-007, 2.750555e-007, 2.907016e-007, 2.815123e-007, 3.33418e-007, 
    3.5875e-007, 3.952578e-007, 4.183546e-007, 4.277921e-007, 4.039501e-007, 
    3.408687e-007, 2.047713e-007, 9.152245e-008, 1.853998e-007, 
    2.929365e-007, 3.858204e-007, 3.512994e-007, 2.760487e-007, 
    3.888008e-007, 2.574225e-007, -6.161827e-010, 1.8987e-007, 5.733268e-007, 
    9.612545e-007, 8.768152e-007, 3.560185e-007, 6.001496e-007, 
    1.430144e-006, 1.655897e-006, 1.325836e-006, 1.27716e-006, 1.394879e-006, 
    1.256049e-006, 7.305352e-007, 6.292066e-007, 2.904526e-007, 
    -2.467359e-007, 3.291934e-007, 1.426914e-006, 1.990921e-006, 
    2.190596e-006, 1.329062e-006, -4.372223e-007, -1.745542e-006, 
    -1.780562e-006, -3.721543e-007, 8.162151e-007, 1.011918e-006, 
    1.01614e-006, 8.817815e-007, 7.454364e-007, 1.046191e-006, 1.294544e-006, 
    1.576424e-006, 1.936286e-006, 1.815091e-006, 1.599272e-006, 
    1.458207e-006, 1.432627e-006, 1.118462e-006, 1.004717e-006, 
    1.155466e-006, 7.874069e-007, 1.369722e-007, -3.490545e-007, 
    -5.2464e-007, -1.645287e-007, 3.505547e-007, 4.702606e-007, 5.07762e-007, 
    4.943508e-007, 5.256434e-007, 4.861552e-007, 3.93768e-007,
  4.312692e-007, 5.112388e-007, 7.948577e-007, 6.483294e-007, -1.675903e-008, 
    -3.011228e-007, -2.072456e-007, -2.452437e-007, 2.918591e-008, 
    1.938436e-007, 1.590744e-007, 1.888766e-007, 1.496371e-007, 
    3.772129e-010, -1.717299e-007, 2.082486e-007, 3.155367e-007, 
    1.002149e-007, 3.191781e-008, 2.373055e-007, 3.118116e-007, 
    4.275439e-007, 5.984116e-007, 6.714267e-007, 4.687708e-007, 
    6.023852e-007, 5.353293e-007, 4.384717e-007, 4.998146e-007, 
    4.389683e-007, 2.700883e-007, 3.721614e-007, 3.450905e-007, 
    1.101491e-007, 3.234838e-007, -9.648011e-008, -5.355678e-007, 
    -4.419387e-007, -7.934386e-008, 3.920297e-007, 3.962518e-007, 
    7.258163e-007, 1.312425e-006, 1.377244e-006, 1.79994e-006, 2.524882e-006, 
    2.903867e-006, 2.658743e-006, 1.858551e-006, 1.631308e-006, 
    1.246362e-006, 1.319129e-006, 1.452742e-006, 1.208363e-006, 
    1.090146e-006, 5.936899e-007, -5.277252e-008, -9.309588e-009, 
    1.071024e-006, 1.758215e-006, 1.060095e-006, -2.445995e-008, 
    -3.123005e-007, 4.630565e-007, 6.41372e-007, 3.638706e-008, 
    -7.934432e-008, 4.287858e-007, 3.165305e-007, 1.245544e-007, 
    -2.147726e-008, 3.090804e-007, 4.690196e-007, 7.427043e-007, 
    1.281381e-006, 9.751625e-007, 1.521212e-007, 1.428543e-008, 
    8.226739e-007, 2.125035e-006, 3.027052e-006, 2.618264e-006, 
    1.541655e-006, 8.974284e-007, 1.021356e-006, 1.27691e-006, 1.229972e-006, 
    1.388918e-006, 1.313419e-006, 8.887364e-007, 1.926032e-007, 
    -8.008874e-008, 4.990698e-007, -5.128004e-008, -2.298448e-007, 
    -3.414289e-008,
  1.930998e-007, 7.81695e-007, 9.801283e-007, 1.933472e-007, -6.632206e-007, 
    -1.190969e-006, -1.119445e-006, -5.92936e-007, 3.840833e-007, 
    4.267986e-007, 6.811117e-007, 8.666314e-007, 1.030048e-006, 
    1.055877e-006, 7.658009e-007, -2.536863e-007, -4.963276e-007, 
    -1.456533e-007, 3.920304e-007, 1.950862e-007, 6.49502e-008, 
    7.886497e-007, 2.320241e-006, 2.998988e-006, 2.386548e-006, 
    1.694638e-006, 1.808882e-006, 1.668812e-006, 2.020402e-007, 
    -1.121928e-006, -8.748175e-007, -1.203216e-007, 1.373519e-006, 
    1.535196e-006, 7.146382e-007, 1.913586e-007, -1.831577e-007, 
    -4.118892e-007, -1.776934e-007, 5.790371e-007, 6.160417e-007, 
    2.79415e-008, 1.322606e-006, 1.572945e-006, 2.097465e-006, 3.466882e-006, 
    4.500277e-006, 4.280981e-006, 2.609319e-006, 1.968569e-006, 
    2.416349e-006, 1.777587e-006, 6.997352e-007, 4.064314e-007, 
    2.054748e-006, 2.074866e-006, 9.624182e-008, -6.570144e-007, 
    -4.173535e-007, -3.175155e-007, 3.381347e-007, 1.216311e-006, 
    1.323848e-006, 1.840918e-006, 2.390275e-006, 1.67477e-006, 1.900771e-006, 
    1.248598e-006, 1.25133e-006, 1.273183e-006, 3.552705e-007, 6.073496e-007, 
    1.508125e-006, 1.942993e-006, 1.670549e-006, 1.990179e-006, 
    2.074371e-006, 2.496569e-006, 2.486385e-006, 2.525624e-006, 
    2.768016e-006, 1.755734e-006, 8.594297e-007, 4.47661e-007, 9.180408e-007, 
    2.381335e-006, 1.773615e-006, 1.38246e-006, 1.471868e-006, 8.422926e-007, 
    8.904735e-007, 1.72171e-006, 3.091375e-006, 2.221396e-006, 4.600788e-007, 
    -2.445722e-008,
  9.873274e-007, 3.773739e-007, 7.464259e-007, 1.220532e-006, 1.785039e-006, 
    2.033641e-006, 1.855075e-006, 1.813601e-006, 2.690782e-006, 
    2.515694e-006, 2.031157e-006, 3.038723e-006, 3.462165e-006, 
    1.635283e-006, 1.353403e-006, 1.692901e-006, 1.216312e-006, 
    7.066919e-007, -3.018686e-007, -1.205874e-006, -3.81342e-007, 
    8.666302e-007, 1.623113e-006, 3.238398e-006, 3.267953e-006, 
    2.668182e-006, 2.851963e-006, 4.370638e-006, 3.500163e-006, 
    2.909577e-006, 9.927926e-007, 1.13038e-006, 2.570083e-006, 2.787141e-006, 
    3.319359e-006, 2.640611e-006, 1.496949e-006, 4.553567e-007, 
    1.828002e-006, 1.71078e-006, 1.786776e-006, 1.83123e-006, 1.484778e-006, 
    9.560363e-007, 2.658644e-007, 2.872239e-007, 6.229939e-007, 
    1.715499e-006, 3.745533e-006, 4.666177e-006, 3.416217e-006, 
    1.122929e-006, 1.120695e-006, 1.773117e-006, 1.967329e-006, 2.38158e-006, 
    2.541022e-006, 2.89567e-006, 2.968935e-006, 1.482545e-006, 3.038613e-007, 
    4.640497e-007, -7.323251e-009, -1.67759e-007, 1.413253e-006, 
    2.13422e-006, 2.682086e-006, 2.436962e-006, 2.122795e-006, 2.97862e-006, 
    3.538406e-006, 2.681341e-006, 2.225366e-006, 2.296892e-006, 2.88822e-006, 
    2.292173e-006, 2.2656e-006, 2.73747e-006, 2.641606e-006, 2.599882e-006, 
    2.531834e-006, 2.223131e-006, 1.740333e-006, 2.038855e-006, 
    3.250816e-006, 4.383553e-006, 3.927329e-006, 2.353271e-006, 
    1.927843e-006, 2.13025e-006, 2.483405e-006, 3.669289e-006, 2.782422e-006, 
    2.164275e-006, 1.793484e-006, 1.928834e-006,
  2.002594e-006, 1.560527e-006, 1.088903e-006, 2.189107e-006, 4.698214e-006, 
    3.609684e-006, 2.254424e-006, 1.993404e-006, 1.906233e-006, 
    4.052497e-006, 3.947443e-006, 4.241493e-006, 4.306065e-006, 4.9791e-006, 
    3.68866e-006, 2.93044e-006, 4.46203e-006, 3.130612e-006, 2.572315e-006, 
    2.081818e-006, 1.316894e-006, 2.530841e-006, 3.686177e-006, 
    3.381199e-006, 4.146623e-006, 4.209951e-006, 4.232304e-006, 
    5.261229e-006, 5.523737e-006, 5.182999e-006, 5.29103e-006, 4.522877e-006, 
    4.798548e-006, 3.260498e-006, 3.130113e-006, 3.001716e-006, 
    2.813963e-006, 2.073623e-006, 2.454843e-006, 2.524631e-006, 
    1.693146e-006, 2.783665e-006, 2.589452e-006, 1.052646e-006, 
    1.115477e-006, 3.635512e-006, 4.934645e-006, 3.799425e-006, 
    3.989663e-006, 3.245599e-006, 2.563374e-006, 5.600668e-008, 
    4.059348e-007, 1.537926e-006, 2.522644e-006, 3.332522e-006, 
    3.026801e-006, 2.649057e-006, 4.413851e-006, 3.425407e-006, 
    1.657882e-006, -7.264134e-008, -1.435599e-006, 2.75797e-007, 
    1.948951e-006, 3.009914e-006, 3.271677e-006, 3.525989e-006, 
    2.857672e-006, 3.91615e-006, 4.148361e-006, 3.129368e-006, 3.777072e-006, 
    4.077084e-006, 4.101918e-006, 4.72007e-006, 3.649669e-006, 4.534052e-006, 
    4.337109e-006, 3.765899e-006, 2.470988e-006, 2.768514e-006, 
    2.757835e-006, 3.033754e-006, 3.372011e-006, 3.116455e-006, 
    3.023324e-006, 3.27714e-006, 4.092978e-006, 1.951185e-006, 9.878249e-007, 
    2.234556e-006, 3.80936e-006, 4.2482e-006, 3.526486e-006, 2.817439e-006,
  2.925223e-006, 3.594783e-006, 3.647432e-006, 4.018224e-006, 4.741428e-006, 
    3.955639e-006, 4.13495e-006, 3.730384e-006, 3.720201e-006, 5.0772e-006, 
    8.305785e-006, 8.412078e-006, 5.29451e-006, 5.000955e-006, 5.010393e-006, 
    5.84759e-006, 5.329279e-006, 5.677965e-006, 7.226692e-006, 6.204721e-006, 
    5.602714e-006, 6.062415e-006, 7.679439e-006, 7.814791e-006, 
    5.921351e-006, 5.778298e-006, 7.374461e-006, 7.787721e-006, 
    7.448224e-006, 6.68876e-006, 6.003555e-006, 5.577136e-006, 5.495427e-006, 
    5.194422e-006, 6.008771e-006, 4.178658e-006, 1.89158e-006, 3.041205e-006, 
    3.939247e-006, 4.503008e-006, 4.916021e-006, 5.629041e-006, 
    4.988789e-006, 6.849696e-006, 8.480127e-006, 8.322424e-006, 
    7.183977e-006, 6.136423e-006, 3.848103e-006, 5.281347e-006, 
    5.275886e-006, 3.377972e-006, 3.436584e-006, 4.105397e-006, 
    3.761927e-006, 3.531204e-006, 1.583374e-006, 1.026319e-006, 
    2.087283e-006, 3.240635e-006, 2.958254e-006, 3.118939e-006, 
    1.395125e-006, 1.434113e-006, 3.26646e-006, 4.362195e-006, 3.246098e-006, 
    1.29181e-006, 1.06978e-006, 3.051387e-006, 4.742174e-006, 3.469118e-006, 
    3.684938e-006, 2.737721e-006, 2.757091e-006, 2.438952e-006, 
    4.002331e-006, 3.997862e-006, 4.149357e-006, 6.139158e-006, 
    6.576009e-006, 5.531685e-006, 4.10639e-006, 5.395091e-006, 4.6098e-006, 
    2.321975e-006, 1.887607e-006, 3.199653e-006, 3.658859e-006, 
    2.782669e-006, 4.220383e-006, 6.078559e-006, 4.835554e-006, 
    4.241741e-006, 2.398468e-006, 2.375372e-006,
  6.708135e-006, 7.30443e-006, 7.830937e-006, 8.086241e-006, 6.752092e-006, 
    4.932661e-006, 4.804759e-006, 3.295521e-006, 2.620747e-006, 
    5.608428e-006, 8.660187e-006, 1.117004e-005, 9.372212e-006, 
    8.780888e-006, 5.880873e-006, 8.553645e-006, 1.091275e-005, 
    9.480496e-006, 8.603814e-006, 7.396569e-006, 7.608664e-006, 
    8.214147e-006, 8.221597e-006, 6.651262e-006, 9.155154e-006, 
    1.019178e-005, 9.140751e-006, 1.26152e-005, 1.477339e-005, 1.348693e-005, 
    1.051538e-005, 7.095568e-006, 5.259493e-006, 5.458423e-006, 5.30519e-006, 
    5.177539e-006, 5.990396e-006, 4.999716e-006, 6.310025e-006, 
    6.316483e-006, 4.977363e-006, 3.090629e-006, 3.595535e-006, 
    7.273882e-006, 9.726366e-006, 6.408123e-006, 3.864992e-006, 
    4.452349e-006, 6.127737e-006, 5.791217e-006, 7.236134e-006, 
    7.875891e-006, 6.56583e-006, 3.404548e-006, 2.418588e-006, 1.222521e-006, 
    2.179671e-006, 1.222023e-006, 2.022465e-006, 1.978256e-006, 2.31999e-006, 
    4.151845e-006, 3.962348e-006, 3.921867e-006, 5.529704e-006, 
    4.739944e-006, 2.580015e-006, 1.185515e-006, 4.31501e-006, 5.478543e-006, 
    3.387162e-006, 1.933306e-006, 1.745799e-006, 2.853205e-006, 
    3.807127e-006, 3.622103e-006, 2.646078e-006, 1.42791e-006, 3.210336e-006, 
    1.979748e-006, 1.036897e-007, 6.679493e-007, 2.973655e-006, 
    4.270054e-006, 3.43584e-006, 2.108642e-006, 1.56301e-006, 2.135217e-006, 
    2.660729e-006, 4.963207e-006, 6.523362e-006, 6.910295e-006, 
    7.054838e-006, 5.112221e-006, 4.974387e-006, 6.170205e-006,
  1.814595e-006, 4.903854e-006, 5.438806e-006, 4.347052e-006, 3.950183e-006, 
    4.197787e-006, 4.821399e-006, 5.318352e-006, 6.126489e-006, 
    1.010585e-005, 7.816037e-006, 5.965063e-006, 6.33188e-006, 7.433579e-006, 
    7.491693e-006, 1.033558e-005, 1.368114e-005, 1.207727e-005, 
    8.496523e-006, 7.858258e-006, 9.131063e-006, 1.10101e-005, 9.689862e-006, 
    9.564192e-006, 8.509436e-006, 7.764131e-006, 8.988263e-006, 
    9.795418e-006, 9.999561e-006, 8.204217e-006, 7.90718e-006, 8.830559e-006, 
    6.361681e-006, 4.613526e-006, 3.80663e-006, 1.166392e-006, 1.291068e-006, 
    1.060842e-006, 1.221277e-006, 2.976138e-006, 5.129357e-006, 
    5.495678e-006, 4.89963e-006, 3.210831e-006, 3.849349e-006, 1.67502e-006, 
    2.615032e-006, 6.066639e-006, 7.542598e-006, 5.83592e-006, 3.926336e-006, 
    5.174807e-006, 6.338838e-006, 5.614142e-006, 9.302927e-006, 
    7.147968e-006, 4.68729e-006, 5.672751e-006, 2.333651e-006, 1.80913e-006, 
    1.934299e-006, 1.572946e-006, 1.183778e-006, 7.77969e-007, 1.557548e-006, 
    1.953671e-006, 2.441686e-006, 3.427893e-006, 3.288569e-006, 
    3.722935e-006, 2.736973e-006, 1.936038e-006, 2.972911e-006, 
    3.105035e-006, 2.128512e-006, 2.196317e-006, 1.101082e-006, 
    -4.344289e-006, -2.44267e-006, -4.071726e-007, -1.510852e-006, 
    -4.963276e-007, 1.157949e-006, 1.062335e-006, 1.213331e-006, 
    2.297142e-006, 5.321333e-006, 6.714841e-006, 7.654855e-006, 
    7.033233e-006, 4.847974e-006, 5.170088e-006, 3.87716e-006, 3.508852e-006, 
    2.986069e-006, 1.816334e-006,
  2.284731e-006, 2.913304e-006, 1.079719e-006, 6.751525e-007, 2.069899e-006, 
    2.595414e-006, 1.633296e-006, 9.023934e-007, 2.157818e-006, 3.4649e-006, 
    3.007432e-006, 3.968562e-006, 5.767135e-006, 6.745391e-006, 
    6.929175e-006, 9.076928e-006, 6.877268e-006, 5.027287e-006, 
    8.405132e-006, 9.647887e-006, 9.472056e-006, 8.956726e-006, 
    7.632014e-006, 6.617003e-006, 5.095837e-006, 2.072895e-006, 
    1.782315e-006, 1.633056e-006, -2.160035e-006, -3.39187e-006, 
    -1.506374e-006, -7.225772e-007, -2.893428e-006, -2.765777e-006, 
    -3.003697e-006, -4.137428e-006, -4.870317e-006, -2.936391e-006, 
    7.066228e-008, -2.688357e-007, 8.208553e-008, -2.946654e-007, 
    -1.98222e-006, -5.817601e-007, 1.100583e-006, 4.141402e-007, 
    1.941509e-006, 1.290075e-006, 1.906732e-006, -4.759659e-007, 
    2.264609e-006, 2.12851e-006, 1.232951e-006, 3.128376e-006, 1.863767e-006, 
    -1.409522e-006, -1.975019e-006, -7.610724e-007, 7.388917e-008, 
    2.255416e-006, 1.412513e-006, -8.003117e-007, 6.637274e-007, 
    1.42468e-006, 1.044391e-007, 9.673749e-008, 7.501549e-007, 1.10679e-006, 
    1.144539e-006, 2.201705e-007, -2.333143e-006, -2.214681e-006, 
    -2.72008e-006, -4.305315e-006, -3.646683e-006, -6.383765e-006, 
    -9.631476e-006, -1.32825e-005, -6.738426e-006, -3.077459e-006, 
    -3.655872e-006, -2.444905e-006, -2.909324e-006, -2.819172e-006, 
    -1.232196e-006, 3.193702e-006, 8.083516e-006, 8.644052e-006, 
    7.80437e-006, 6.749116e-006, 3.699595e-006, 2.203513e-006, 3.67302e-006, 
    4.357978e-006, 3.053883e-006, 1.500437e-006,
  -7.923554e-007, -2.893426e-006, -2.479177e-006, -1.748771e-006, 
    -3.020585e-006, -5.451213e-006, -4.096697e-006, -1.614661e-006, 
    -1.285593e-006, -7.059371e-007, 8.542156e-007, 2.212459e-006, 
    -7.061826e-007, -1.298249e-006, -7.506351e-007, -7.079216e-007, 
    3.796205e-006, 6.424274e-006, 6.107872e-006, 6.374856e-006, 
    1.279153e-006, -1.641722e-006, -3.442525e-006, -5.57438e-006, 
    -7.957078e-006, -7.090333e-006, -4.742411e-006, -6.166714e-006, 
    -8.528803e-006, -9.12261e-006, -9.831409e-006, -1.108211e-005, 
    -1.21247e-005, -1.242247e-005, -1.018978e-005, -1.004152e-005, 
    -1.053052e-005, -9.193889e-006, -9.899706e-006, -9.572132e-006, 
    -7.525454e-006, -6.892902e-006, -4.990023e-006, -2.060453e-006, 
    -1.914919e-006, -4.566078e-006, -5.580598e-006, -2.335875e-006, 
    -3.168108e-006, -3.160905e-006, -9.992455e-007, 1.378976e-008, 
    -7.305225e-007, -8.395509e-007, -3.885845e-006, -5.512062e-006, 
    -2.246221e-006, -2.166496e-006, 1.736364e-006, 1.790753e-006, 
    3.776258e-007, -2.423543e-006, -1.485514e-006, -1.459439e-006, 
    -1.988681e-006, -9.875712e-007, -1.434852e-006, -1.955401e-006, 
    -2.36543e-006, -5.881113e-006, -7.899474e-006, -6.874277e-006, 
    -9.57958e-006, -8.670608e-006, -9.27808e-006, -9.918086e-006, 
    -9.559712e-006, -1.079105e-005, -6.213656e-006, -3.14079e-006, 
    -4.049261e-006, -6.540489e-006, -4.722049e-006, -1.975262e-006, 
    6.279733e-007, 6.411858e-006, 6.101669e-006, 7.741037e-006, 
    8.015464e-006, 4.919006e-006, 2.88376e-006, 2.379602e-006, 8.698626e-007, 
    2.04557e-006, 1.07575e-006, 1.045701e-006,
  -5.173059e-006, -6.352982e-006, -6.620956e-006, -6.142379e-006, 
    -5.41545e-006, -4.625193e-006, -3.836923e-006, -5.040685e-006, 
    -3.4105e-006, -2.688288e-006, -2.604595e-006, -6.614247e-006, 
    -1.104386e-005, -1.088045e-005, -9.078394e-006, -7.680173e-006, 
    -5.873902e-006, -2.21741e-006, -4.604328e-006, -7.692834e-006, 
    -8.909763e-006, -6.988012e-006, -7.234134e-006, -7.531167e-006, 
    -6.552906e-006, -5.679451e-006, -7.436051e-006, -7.79889e-006, 
    -7.91487e-006, -7.03893e-006, -8.378544e-006, -9.476512e-006, 
    -8.861341e-006, -8.760014e-006, -8.567294e-006, -8.820364e-006, 
    -1.03758e-005, -9.450934e-006, -1.122243e-005, -1.043838e-005, 
    -7.591266e-006, -4.614018e-006, -2.600127e-006, 1.364715e-007, 
    -3.728946e-007, -3.261737e-006, -5.574148e-006, -5.772084e-006, 
    -6.481629e-006, -4.431477e-006, 1.22153e-006, -2.31675e-006, 
    -5.116433e-006, -6.540242e-006, -6.075074e-006, -2.404917e-006, 
    -2.134462e-006, -3.346669e-006, -1.774846e-006, -3.347415e-006, 
    -2.826129e-006, -1.567223e-006, -3.107511e-006, -3.581612e-006, 
    -1.96136e-006, -3.808609e-006, -4.742167e-006, -4.419806e-006, 
    -4.826854e-006, -5.584081e-006, -5.894273e-006, -7.361296e-006, 
    -7.337203e-006, -5.121651e-006, -4.274022e-006, -4.687529e-006, 
    -6.692728e-006, -7.520238e-006, -1.949938e-006, -1.660856e-006, 
    -3.788244e-006, -5.822585e-007, 3.737594e-006, 8.708372e-006, 
    8.713589e-006, 7.219998e-006, 9.901214e-006, 6.622955e-006, 
    4.228339e-006, 1.30945e-006, 1.368313e-006, 4.069407e-007, 
    -2.208213e-006, -5.414946e-006, -6.759026e-006, -6.993976e-006,
  -4.569315e-006, -4.272035e-006, -2.719333e-006, -1.718969e-006, 
    -8.318525e-007, -1.491725e-006, -2.036364e-006, -1.88164e-006, 
    -1.17011e-006, -1.937769e-006, -5.871429e-006, -1.053773e-005, 
    -9.956082e-006, -9.00936e-006, -7.700792e-006, -5.555521e-006, 
    -3.119183e-006, -7.845583e-006, -9.340667e-006, -6.258855e-006, 
    -2.276771e-006, -4.080057e-006, -4.222613e-006, -3.986925e-006, 
    -3.969046e-006, -3.761422e-006, -3.150972e-006, -1.887353e-006, 
    -1.925846e-006, -1.812349e-006, -3.664813e-006, -4.657232e-006, 
    -3.413233e-006, -2.362203e-006, -1.153968e-006, -1.937272e-006, 
    -3.496181e-006, -4.112841e-006, -4.099182e-006, -4.660707e-006, 
    -2.888461e-006, 3.112233e-006, 2.774228e-006, 8.375737e-007, 
    -2.509971e-006, -4.0659e-006, -4.496795e-006, -2.22412e-006, 
    -2.497307e-006, 8.907191e-007, -1.868724e-006, -6.056696e-006, 
    -5.283076e-006, -3.180025e-006, -1.678491e-006, 1.102067e-006, 
    2.132165e-007, -1.914665e-006, -3.02282e-006, -2.408146e-006, 
    -1.173092e-006, -2.021958e-006, -3.507354e-006, -3.649664e-006, 
    -5.113701e-006, -6.880235e-006, -2.559145e-006, -2.046547e-006, 
    -4.658718e-006, -5.620339e-006, -4.906574e-006, -3.591052e-006, 
    -3.430368e-006, -3.884605e-006, -3.275646e-006, -2.168239e-006, 
    -2.36394e-006, -1.332531e-006, 1.618893e-006, 5.333752e-006, 
    1.029187e-005, 1.310272e-005, 1.050049e-005, 4.996989e-006, 
    2.482913e-006, 6.448612e-006, 6.517155e-006, 2.341108e-006, 
    -5.745533e-007, -3.19715e-006, -6.370112e-006, -5.504102e-006, 
    -4.59042e-006, -6.69124e-006, -3.803396e-006, -3.343939e-006,
  -2.045055e-006, -8.328457e-007, -2.668501e-007, -4.374683e-007, 
    -6.999772e-007, -9.82851e-007, 1.49887e-007, 6.035842e-006, 1.19002e-005, 
    1.317396e-006, -3.48848e-006, -1.837187e-006, -1.785777e-006, 
    -2.427768e-006, -2.687299e-006, 6.617393e-007, -2.829354e-006, 
    -2.675375e-006, -6.227419e-007, 5.61653e-007, -3.984796e-007, 
    -1.401575e-006, -1.62544e-007, -7.572453e-009, -2.089841e-007, 
    2.576717e-007, -1.786848e-007, -1.282688e-007, -3.525311e-007, 
    -1.138567e-006, -1.536678e-006, -3.676815e-007, 1.16987e-006, 
    1.427412e-006, 4.173621e-007, -1.24064e-006, -1.526991e-006, 
    -1.381208e-006, -1.231453e-006, -4.709973e-007, 4.518824e-007, 
    -3.245839e-006, -3.442785e-006, -5.937487e-006, -3.68766e-006, 
    -2.453347e-006, -8.922043e-007, 5.521006e-006, 5.065032e-006, 
    3.621359e-006, -3.793955e-006, -3.756702e-006, 1.975059e-008, 
    4.180649e-006, 2.594177e-006, 4.050513e-006, 1.880409e-006, 
    -5.403532e-006, -3.775578e-006, -6.771334e-007, 2.199042e-006, 
    -4.290214e-007, -2.632158e-006, -7.071218e-006, -1.06912e-005, 
    -3.894291e-006, -1.607954e-006, -5.120657e-006, -5.596997e-006, 
    -4.177661e-006, -3.288558e-006, -3.375731e-006, -1.700841e-006, 
    -1.260757e-006, -1.49868e-006, -7.570179e-009, 2.527031e-007, 
    4.973306e-007, 1.366566e-006, 9.920837e-006, 1.627742e-005, 
    1.515139e-005, 1.633156e-005, 9.170803e-006, 6.13643e-006, 3.97009e-007, 
    4.101639e-007, -4.206457e-006, -8.326631e-006, -4.658221e-006, 
    -5.980701e-006, -6.416809e-006, -3.180774e-006, -2.612543e-006, 
    -3.023566e-006, -3.10428e-006,
  -2.805086e-007, 1.456647e-007, -2.713205e-007, -2.147681e-008, 
    -5.991459e-007, 1.388669e-006, 4.814691e-006, 1.445748e-005, 
    2.224831e-005, 2.674391e-006, -2.29465e-006, -1.156948e-006, 
    -2.857287e-007, -1.441804e-006, -1.203189e-007, -2.116332e-006, 
    1.570712e-006, 2.362458e-006, 9.582727e-007, 1.051652e-006, 
    1.646208e-006, 2.09225e-006, 1.818566e-006, 2.681018e-007, 1.496373e-007, 
    -2.084867e-007, 8.084362e-008, -1.051893e-006, -8.676154e-007, 
    -9.244877e-007, -7.3276e-007, -4.354822e-007, 2.034137e-006, 
    3.808541e-007, 8.283864e-007, -6.594951e-007, -1.12317e-006, 
    -5.862312e-007, 9.046298e-007, 2.233065e-006, 9.667165e-007, 
    -4.279982e-006, -5.714965e-006, -5.246075e-006, -8.928055e-008, 
    -1.145277e-006, 2.743091e-007, 9.965279e-006, 1.466586e-005, 
    9.317826e-006, 7.672737e-006, 1.39131e-005, 9.70178e-006, 7.203103e-006, 
    2.818688e-006, -3.004436e-006, -2.183137e-006, -9.468349e-007, 
    -2.030141e-006, 1.287102e-006, 1.461704e-007, -5.118667e-006, 
    -7.604178e-006, -7.67571e-006, -4.211437e-006, -2.778937e-006, 
    -4.02219e-006, -2.816441e-006, -1.515072e-006, -3.062062e-006, 
    -1.438083e-006, -1.306207e-006, -7.744825e-007, -2.949128e-007, 
    6.271512e-008, 4.777125e-007, 2.899562e-007, 7.91877e-007, 3.28946e-007, 
    1.933066e-005, 1.098129e-005, 1.207603e-005, 2.347344e-005, 
    2.048948e-005, 8.878749e-006, 2.467525e-006, -7.560961e-006, 
    -5.598235e-006, -8.63485e-006, -1.018457e-005, -7.406988e-006, 
    -6.174168e-006, -3.663818e-006, -2.917023e-006, -1.487503e-006, 
    -7.521307e-007,
  -2.710722e-007, -3.579953e-007, 5.219179e-007, 2.527036e-007, 
    7.439421e-007, 1.256281e-005, 1.367915e-005, 9.614609e-006, 
    3.797701e-006, -1.568715e-006, -1.992896e-006, -6.719092e-007, 
    1.398359e-006, -4.428486e-006, -3.788977e-006, 1.404322e-006, 
    9.088508e-007, 2.04581e-006, -1.289069e-006, -2.803527e-006, 
    -1.575176e-006, 9.549422e-008, 9.605064e-007, -3.166315e-008, 
    -8.877341e-007, -1.777333e-006, -7.27794e-007, -1.130869e-006, 
    -7.844169e-007, -4.300177e-007, -3.932616e-007, 2.874727e-007, 
    5.25315e-008, -1.286835e-006, -4.685123e-007, -1.073498e-006, 
    -5.450047e-007, 1.104803e-006, 2.256413e-006, 3.324221e-007, 
    -1.112741e-006, -4.396955e-006, -6.039561e-006, -4.161102e-007, 
    7.797062e-007, 7.946171e-006, 1.27128e-005, 1.720998e-005, 7.546081e-006, 
    8.307283e-006, 7.236387e-006, 1.500038e-005, 1.035942e-005, 
    3.574925e-006, -2.428256e-006, -1.542952e-005, -1.294128e-005, 
    -2.562367e-006, -5.13182e-006, -6.874016e-006, -5.263944e-006, 
    -2.84176e-006, -1.09163e-006, -1.909206e-006, -6.666996e-007, 
    -2.153834e-006, -1.290173e-007, 5.643842e-007, -4.486465e-007, 
    -8.083589e-008, -1.096102e-006, -1.27889e-006, -4.185927e-007, 
    1.801836e-007, 5.029619e-008, -5.601544e-007, -6.146297e-008, 
    6.77138e-007, -6.14387e-006, 2.544752e-006, 8.623436e-006, 1.171021e-005, 
    1.935574e-005, 1.320082e-005, 1.392825e-005, 1.047691e-006, 
    -1.479498e-005, -1.805809e-005, -1.348443e-005, -7.9253e-006, 
    -6.177645e-006, -2.307317e-006, -1.785528e-006, -1.56375e-006, 
    -8.199331e-007, -6.237324e-007,
  -8.909619e-007, 1.151175e-007, 6.239907e-007, -9.499036e-008, 
    3.333764e-006, 1.53605e-005, 1.979211e-005, 4.939873e-006, 3.980727e-006, 
    3.438508e-007, -3.515048e-006, 3.194196e-006, 1.529667e-005, 
    -6.498085e-007, -2.992761e-006, 2.971683e-007, 3.509354e-006, 
    2.801795e-006, 2.815123e-007, -1.43858e-006, -1.862271e-006, 
    2.895174e-006, 1.739092e-006, 1.726403e-008, -1.719715e-006, 
    -2.553684e-006, -2.733987e-006, -1.986693e-006, -1.163652e-006, 
    -3.624662e-007, 1.173514e-007, -1.626581e-006, -1.241387e-006, 
    -2.369901e-006, -2.773225e-006, 4.526278e-007, 1.751016e-006, 
    2.919266e-006, 2.284974e-006, -2.465767e-006, -1.708043e-006, 
    1.230714e-006, -1.620447e-007, 2.598146e-006, 7.518262e-006, 
    1.364289e-005, 1.38597e-005, 9.357813e-006, 1.002986e-005, 1.269642e-005, 
    5.247832e-006, 7.758423e-006, 9.177253e-006, -6.730734e-006, 
    -1.857019e-005, -1.105057e-005, -3.530695e-006, -2.525114e-006, 
    -4.425761e-006, 1.633809e-006, 4.617763e-006, 5.548336e-006, 
    7.255694e-007, -9.361629e-007, 3.746445e-007, -7.263034e-007, 
    2.762945e-007, 2.719753e-008, -1.362584e-006, -1.747282e-006, 
    -1.917901e-006, -1.440816e-006, -5.189304e-007, -1.647442e-006, 
    -1.446277e-006, -3.070863e-007, -3.808443e-007, -2.127097e-007, 
    -1.241303e-005, 3.354631e-006, 1.806804e-005, 1.852575e-005, 
    1.188927e-005, 3.035733e-006, -8.715309e-006, -2.360355e-005, 
    -2.515948e-005, -1.241179e-005, -5.915632e-006, -2.714368e-006, 
    -1.05562e-006, -5.181846e-007, -9.319401e-007, -1.356623e-006, 
    -1.102807e-006, -1.054131e-006,
  -1.190474e-006, -6.469054e-008, -5.993948e-007, 1.163662e-006, 
    8.253148e-006, 1.191163e-005, 1.533517e-005, 1.042076e-005, 
    5.804883e-006, 3.706551e-006, -7.735554e-006, 2.2815e-006, 1.204425e-005, 
    -1.911681e-006, -2.546469e-006, 2.023713e-006, 1.197496e-005, 
    6.856899e-006, 2.401202e-006, -2.498302e-006, -3.031015e-006, 
    2.003339e-006, 1.90375e-006, -5.780385e-007, -1.376739e-006, 
    -2.789619e-006, -2.425782e-006, -1.660109e-006, -5.219085e-007, 
    -4.979211e-008, -8.321022e-007, 2.707427e-006, 3.106776e-006, 
    -2.780678e-006, -3.41646e-006, -3.691721e-007, -2.338188e-007, 
    1.057118e-006, 5.058822e-006, 2.343086e-006, -1.562506e-006, 
    -4.767244e-006, -6.003829e-007, 5.203867e-006, -7.267881e-007, 
    4.624468e-006, 1.461719e-005, 1.676717e-005, 2.33433e-005, 2.541928e-005, 
    3.089271e-005, 2.17968e-005, 1.485039e-005, 1.532524e-005, 7.38143e-006, 
    8.954979e-006, 1.177329e-005, 1.268028e-005, 1.179092e-005, 
    1.017017e-005, 9.569416e-006, 2.036872e-006, -3.704135e-007, 
    -3.458263e-007, -1.002081e-007, -1.891576e-006, -1.330299e-006, 
    -2.408398e-006, -2.678852e-006, -3.065043e-006, -2.343578e-006, 
    -2.67314e-006, -2.872072e-006, -2.848726e-006, -4.789463e-007, 
    -6.287004e-007, -9.716755e-007, -6.878497e-006, -2.699803e-005, 
    1.522366e-005, 1.969574e-005, 7.120652e-006, 2.777961e-006, 
    3.383902e-007, -1.472892e-005, -2.284633e-005, -1.831488e-005, 
    -6.951761e-006, -3.168357e-006, -1.469624e-006, -9.474388e-008, 
    -5.395441e-007, -7.705112e-007, -9.401365e-007, -1.531464e-006, 
    -9.446067e-007,
  -2.288195e-006, -1.686436e-006, 1.970734e-007, 5.149474e-006, 
    1.230005e-005, 1.407576e-005, 1.925764e-005, 1.555719e-005, 
    5.527967e-006, -3.454697e-006, -1.310544e-005, -1.16424e-005, 
    1.290318e-007, -5.638722e-007, -1.140522e-005, -4.215908e-006, 
    5.808608e-006, 1.613139e-005, 1.374373e-005, 5.971782e-006, 
    1.012086e-007, 5.466374e-006, 3.90125e-006, -4.910798e-006, 
    -4.739188e-006, -3.466378e-006, 1.10892e-007, 1.753e-006, 3.61192e-006, 
    2.987319e-006, 3.802172e-006, 6.202499e-006, 6.855662e-006, 
    6.697708e-006, -3.681453e-006, 4.090249e-006, 2.132236e-006, 
    5.002454e-006, 6.464749e-006, 2.958752e-006, -7.938459e-006, 
    -4.561611e-006, -4.256381e-006, 1.578395e-005, 2.214438e-006, 
    7.990871e-006, 2.387179e-005, 2.377071e-005, 3.824024e-005, 
    4.551822e-005, 5.19339e-005, 4.458638e-005, 1.786761e-005, 2.708099e-005, 
    2.753622e-005, 1.94387e-005, 1.660028e-005, 2.51133e-005, 2.349927e-005, 
    1.329421e-005, 6.910293e-006, -1.314404e-006, -2.126268e-006, 
    3.365494e-008, -4.223211e-007, -1.822285e-006, -2.557658e-006, 
    -3.691884e-006, -3.603472e-006, -3.289801e-006, -3.174564e-006, 
    -2.345564e-006, -3.180028e-006, -1.122177e-006, 8.472599e-007, 
    -7.471635e-007, 4.707905e-006, -1.819208e-007, 1.75499e-006, 
    1.059859e-005, 2.566856e-006, -8.666248e-007, -6.752824e-006, 
    -2.259876e-006, -1.688263e-005, -1.47622e-005, -1.206062e-005, 
    -4.994741e-006, -1.39959e-006, -1.277151e-006, -6.676937e-007, 
    -1.135094e-006, -1.512091e-006, -2.257896e-006, -2.239269e-006, 
    -2.220643e-006,
  -9.128153e-007, -8.020493e-007, 2.204008e-006, 5.886091e-006, 
    2.799567e-006, 1.196699e-006, 1.187711e-005, 1.897752e-005, 
    -6.329632e-006, -2.420481e-005, 5.159916e-006, -9.0635e-006, 
    -9.825941e-006, -5.094334e-006, -7.597722e-006, 2.162538e-006, 
    -1.71797e-006, 1.416691e-005, 2.697943e-005, 9.542091e-006, 
    -4.218637e-006, 4.116555e-007, 4.360467e-006, 5.694372e-006, 
    1.155713e-006, -1.3606e-006, 4.638041e-007, 5.428126e-006, 8.506957e-006, 
    8.627405e-006, 1.058841e-005, 4.415349e-006, 6.305803e-006, 
    5.785514e-006, 1.325585e-006, -1.46142e-006, 3.626337e-006, 
    4.863368e-006, 6.675598e-006, -7.712442e-007, 1.161012e-005, 
    1.983433e-005, 9.623807e-006, 3.63314e-005, 3.500445e-005, 2.166419e-005, 
    1.565629e-005, 4.382571e-006, 2.635506e-005, 3.307576e-005, 
    3.733374e-005, 7.903787e-005, 6.82102e-005, 4.487597e-005, 4.511636e-005, 
    4.759891e-005, 4.167644e-005, 3.773037e-005, 3.16867e-005, 2.637171e-005, 
    1.40487e-005, 4.385049e-006, -2.888213e-006, -2.34606e-006, 
    -1.953415e-006, -2.391012e-006, -3.053617e-006, -3.118188e-006, 
    -3.323327e-006, -3.376476e-006, -3.349902e-006, -2.773475e-006, 
    -1.828243e-006, -7.027088e-007, 2.709905e-006, 1.496339e-005, 
    1.11931e-005, -6.128961e-006, 1.124183e-006, -1.988927e-006, 
    8.49404e-006, -1.529719e-006, -1.201268e-005, -1.086853e-005, 
    -5.655849e-006, -4.330148e-006, -2.291175e-006, 3.160923e-006, 
    4.081558e-006, 4.503756e-006, 1.697369e-006, 1.212586e-006, 
    -8.325997e-007, -1.124166e-006, -1.570703e-006, -1.717729e-006,
  6.65151e-006, 7.187452e-006, 9.602687e-006, 7.496405e-006, 1.416734e-006, 
    -5.556518e-006, -3.622343e-006, 1.125573e-005, -9.499352e-006, 
    2.538298e-006, 5.061567e-006, -2.085282e-006, -3.397949e-005, 
    -4.598387e-005, -2.319328e-005, -5.301481e-006, -8.533279e-006, 
    6.205963e-006, 2.028235e-005, 1.259782e-005, 7.389754e-007, 
    -7.590788e-007, 1.761691e-006, 1.233779e-005, 8.578732e-006, 
    7.747003e-006, 1.597741e-005, 2.034295e-005, 1.293211e-005, 
    6.225593e-006, 8.679563e-006, 7.760915e-006, 1.059287e-005, 
    3.573681e-006, 4.158544e-006, 2.067165e-006, 7.506096e-006, 
    5.829701e-006, 1.426869e-005, 1.615697e-005, 2.438587e-005, 
    2.037696e-005, 7.100534e-006, 4.07019e-005, 5.256248e-005, 4.703613e-005, 
    4.974863e-005, 4.812441e-005, 3.969284e-005, 5.881624e-005, 
    5.220484e-005, 8.014874e-005, 8.858901e-005, 7.412447e-005, 
    7.054248e-005, 6.600458e-005, 6.361518e-005, 5.768452e-005, 
    5.412611e-005, 4.768782e-005, 3.947479e-005, 2.818046e-005, 
    1.988697e-005, 8.84968e-006, 5.358336e-006, 1.712022e-006, 8.584329e-007, 
    8.788011e-007, -4.056792e-007, 4.156236e-007, -3.617206e-007, 
    4.116505e-007, 6.845898e-007, -1.998887e-008, 1.964596e-006, 
    -1.065309e-006, -3.582358e-006, 5.890321e-006, -7.155395e-006, 
    -1.767396e-006, -7.511335e-007, -8.864568e-006, -1.192303e-005, 
    -1.424165e-005, -1.18824e-006, 3.712754e-006, 1.880155e-006, 
    7.575141e-006, 9.76288e-006, 1.140598e-005, 1.432462e-005, 1.058642e-005, 
    6.816663e-006, 7.675215e-006, 7.047382e-006, 6.361433e-006,
  7.84584e-006, 5.824004e-006, 9.402767e-006, 4.945083e-006, 2.507259e-007, 
    -3.670022e-006, -1.94732e-005, -1.95192e-005, 5.317837e-006, 
    1.214955e-005, 6.729253e-006, -3.876157e-006, -3.85308e-005, 
    -7.542115e-005, -7.482978e-005, -5.417755e-005, 3.836409e-006, 
    4.804519e-006, -1.853325e-006, 6.234281e-006, -1.189522e-005, 
    -1.11067e-005, -4.593647e-006, 8.023417e-006, 1.402089e-005, 
    5.602473e-006, 1.514891e-005, 3.096095e-006, 1.350665e-006, 
    -6.415794e-006, -5.586589e-007, 2.033475e-005, 3.148728e-005, 
    6.870396e-007, -6.811199e-006, 4.87057e-006, 9.816766e-006, 
    2.298915e-005, 7.257993e-006, 1.205443e-005, 1.787404e-005, 
    1.016843e-005, 4.6637e-006, 1.976875e-005, 1.172359e-005, 5.305519e-005, 
    4.988597e-005, 7.367096e-005, 5.259925e-005, 5.717167e-005, 
    5.106666e-005, 5.1618e-005, 4.419001e-005, 3.792955e-005, 3.144233e-005, 
    2.549924e-005, 2.209756e-005, 1.810926e-005, 1.675524e-005, 
    1.251512e-005, 1.016421e-005, 1.021984e-005, 9.59747e-006, 7.431338e-006, 
    5.764643e-006, 3.753732e-006, 3.172089e-006, 3.002712e-006, 
    3.715484e-006, 3.153959e-006, 4.191078e-006, 6.552662e-006, 
    4.347043e-006, 5.083164e-006, -3.573903e-006, -3.401306e-006, 
    8.974352e-006, 9.012852e-006, 3.441528e-008, -2.942597e-006, 
    -8.640305e-006, -9.998303e-006, -5.353115e-006, -7.747732e-006, 
    -3.22498e-006, 2.17442e-008, 4.556168e-006, 8.028634e-006, 1.021463e-005, 
    8.237253e-006, 1.483945e-005, 9.000934e-006, 8.836269e-006, 
    7.757919e-006, 8.333849e-006, 7.43059e-006,
  6.471706e-006, 7.616618e-006, 1.875196e-006, -1.296264e-005, -1.19668e-006, 
    1.669065e-006, 1.955665e-006, 7.880364e-006, 1.466312e-005, 
    9.883575e-006, 6.393719e-006, 1.181788e-006, -4.296613e-006, 
    -7.603172e-006, 7.173658e-007, -9.170821e-006, 1.43549e-005, 
    8.767471e-006, -1.840254e-005, -1.963313e-005, -1.249648e-005, 
    -7.527939e-006, -7.782728e-006, 6.465925e-007, 5.015107e-006, 
    1.505577e-005, 2.284882e-005, -4.194801e-006, -1.694225e-005, 
    -1.557183e-005, -3.453169e-007, 2.276487e-005, 4.166504e-006, 
    -6.488321e-006, 6.013986e-006, 1.594836e-005, 1.307814e-005, 
    8.99101e-006, -1.381704e-006, -1.654561e-005, -1.246941e-005, 
    -2.456395e-005, -3.704344e-005, -3.987961e-005, -1.995577e-005, 
    5.220019e-006, 7.307412e-006, 3.418091e-005, 3.990445e-005, 
    3.611235e-005, 4.283452e-005, 4.392205e-005, 3.649333e-005, 
    3.009253e-005, 2.813899e-005, 2.775057e-005, 2.670127e-005, 2.32519e-005, 
    2.046836e-005, 2.065984e-005, 1.489086e-005, 1.043492e-005, 
    6.979089e-006, 6.192059e-006, 5.346417e-006, 3.911684e-006, 
    2.748893e-006, 3.356116e-006, 3.241874e-006, 3.973024e-006, 4.91577e-006, 
    4.344562e-006, 5.572665e-006, 9.335465e-006, 7.567691e-006, 
    1.507216e-005, 8.330873e-006, 3.086656e-006, 6.894647e-006, 
    -7.588387e-007, -3.299736e-006, -2.720078e-006, -5.936993e-006, 
    -1.193992e-005, -1.238025e-005, -1.369949e-005, -1.274731e-005, 
    -8.937084e-006, -7.301933e-006, -4.988771e-006, 4.278008e-007, 
    -3.43682e-006, -4.715344e-006, -1.050394e-006, 8.684525e-006, 
    8.324903e-006,
  7.121571e-007, 5.385555e-007, -1.361836e-006, -1.18352e-006, 1.284361e-006, 
    2.102436e-006, 2.33688e-006, 3.259014e-006, 3.136576e-006, 3.254292e-006, 
    1.350382e-005, 5.543108e-006, 3.170235e-007, -8.760435e-007, 
    5.812086e-006, 1.642245e-005, 2.099836e-005, 3.791283e-007, 
    -1.539156e-006, 1.175392e-005, 2.427562e-005, 1.731429e-005, 
    7.221024e-007, 1.227749e-006, 2.053515e-006, 1.435691e-005, 
    1.021835e-005, -1.298847e-005, -1.685035e-005, -1.907758e-005, 
    -1.267331e-005, -1.14278e-005, -1.759118e-005, -4.069298e-007, 
    -1.858542e-006, 9.453914e-006, 1.738581e-005, 1.048932e-005, 
    8.954521e-007, -6.442628e-006, -1.303837e-005, -1.984002e-005, 
    -1.632384e-005, -9.423857e-006, -8.963405e-006, -1.008695e-005, 
    -1.450715e-005, -1.466286e-005, -1.322514e-005, -9.925352e-007, 
    -1.322594e-006, 2.959998e-006, 1.134613e-006, 3.427151e-006, 
    1.120631e-005, 1.57976e-005, 1.450766e-005, 1.422354e-005, 1.299394e-005, 
    1.887469e-005, 2.070207e-005, 2.453439e-005, 1.943324e-005, 
    1.359942e-005, 1.268202e-005, 1.15391e-005, 8.411098e-006, 7.8297e-006, 
    5.206595e-006, 1.563756e-006, -2.112114e-006, -3.146004e-006, 
    -3.061308e-006, 2.076613e-006, 6.172195e-006, 1.29172e-005, 2.5974e-006, 
    -8.282041e-008, 3.996866e-006, -1.293291e-006, -2.271305e-006, 
    -7.097792e-006, -9.782236e-006, -1.268498e-005, -2.284633e-005, 
    -2.2594e-005, -2.089154e-005, -1.927029e-005, -1.639462e-005, 
    -8.508676e-006, -5.81679e-006, -4.277746e-006, -1.510602e-006, 
    4.100182e-006, 1.54985e-006, 8.28883e-007,
  8.333518e-007, 4.938538e-007, 2.397064e-008, 7.243253e-007, 6.803669e-007, 
    4.084208e-007, 1.747209e-007, 3.557699e-007, 4.995661e-007, 
    2.569835e-006, 1.760063e-005, 6.564836e-006, 2.612551e-006, 
    2.287951e-006, 7.476039e-006, 6.776434e-006, 7.702049e-006, 
    6.103401e-007, 1.365134e-005, 2.259651e-005, 8.052464e-006, 
    -1.321603e-006, -6.561095e-006, -5.216765e-006, -5.945685e-006, 
    -3.417204e-006, -2.82414e-006, -2.212694e-006, -8.685261e-006, 
    -1.629503e-005, -1.90058e-005, -2.351391e-005, -1.959241e-005, 
    -2.094667e-005, -3.43448e-005, -5.294496e-006, 4.802278e-006, 
    -4.978938e-008, -8.164956e-006, -1.000824e-005, -9.769567e-006, 
    -7.480747e-006, -1.354205e-005, -1.792696e-005, -1.242768e-005, 
    -7.728846e-006, -5.582082e-006, -2.405258e-005, -2.044948e-005, 
    -1.753058e-005, -2.243579e-005, -1.703786e-005, -1.876364e-005, 
    -2.455424e-005, -2.374014e-005, -3.207237e-005, -3.492867e-005, 
    -4.012372e-005, -4.380877e-005, -3.793449e-005, -3.702851e-005, 
    -2.045048e-005, -1.568931e-005, -1.114891e-005, -8.141615e-006, 
    -4.426511e-006, -3.195913e-006, 2.394248e-006, 3.370529e-006, 
    -1.907461e-006, -2.988781e-007, 3.086408e-006, 1.749668e-007, 
    -2.02196e-006, 9.843516e-007, 3.952163e-006, 4.980739e-007, 
    -1.59529e-006, -1.010916e-006, -3.415465e-006, -9.673706e-006, 
    -7.792184e-006, -5.264948e-006, -1.117624e-005, -1.55686e-005, 
    -1.165457e-005, -1.200822e-005, -5.301456e-006, -1.765164e-006, 
    1.138575e-006, 9.403884e-007, 2.906846e-006, 1.227489e-006, 
    1.120448e-006, 1.098841e-006, 6.686939e-007,
  8.331035e-007, 8.509849e-007, 7.109139e-007, 7.511474e-007, 6.798703e-007, 
    4.978277e-007, 2.139606e-007, 1.809296e-007, 1.332458e-007, 
    8.797938e-007, 2.830605e-006, 1.790503e-006, 1.442064e-006, 
    1.428655e-006, 2.355655e-007, 5.269179e-006, 4.533558e-006, 
    -1.120934e-006, 6.219378e-006, 1.502298e-005, 9.463533e-007, 
    -4.314255e-006, -6.357703e-006, -4.651516e-006, -4.305067e-006, 
    -4.185856e-006, -1.553396e-007, 1.81924e-007, -3.964326e-006, 
    -1.038697e-005, -8.863082e-006, -1.100586e-005, -8.458515e-006, 
    -1.409339e-005, -2.297771e-005, -4.396461e-006, 1.698121e-006, 
    -1.438566e-006, -6.077553e-006, -4.79928e-006, -1.579137e-006, 
    -8.619434e-006, -9.280806e-006, -7.064513e-006, -7.147213e-006, 
    -9.188176e-006, -6.93065e-006, -7.806837e-006, -6.725264e-006, 
    -7.730099e-006, -1.016991e-005, -1.205838e-005, -1.014632e-005, 
    -1.118741e-005, -1.158503e-005, -1.673462e-005, -2.554443e-005, 
    -1.801363e-005, -1.602383e-005, -1.26271e-005, -1.374892e-005, 
    -1.098674e-005, -7.109451e-006, -6.201972e-006, -8.435905e-006, 
    -3.069756e-006, -8.439631e-006, -2.254172e-006, -3.054109e-006, 
    -4.496047e-006, 1.206377e-006, 3.641974e-006, 2.988975e-007, 
    -4.691254e-006, -3.220512e-006, -1.903249e-006, -1.533201e-006, 
    -2.971412e-006, -5.250545e-006, -5.195408e-006, -4.466498e-006, 
    -3.418944e-006, -5.411477e-006, -4.478664e-006, -6.408115e-006, 
    -6.583701e-006, -5.113702e-006, -4.207714e-006, -8.77304e-007, 
    6.324349e-007, 1.261265e-006, 1.152982e-006, 9.167989e-007, 
    2.358154e-007, 4.451767e-007, 9.997487e-007,
  1.320372e-006, 9.813704e-007, 1.201907e-006, 7.163778e-007, 4.561045e-007, 
    5.99404e-007, 4.605749e-007, 1.781977e-007, 2.007978e-007, 1.811779e-007, 
    9.170467e-007, 8.100067e-007, 2.182404e-006, 8.494949e-007, 
    1.056621e-006, 2.696739e-006, 1.893568e-006, -6.671962e-007, 
    4.249439e-006, 7.781759e-006, 3.3817e-006, 1.488755e-006, -7.934523e-008, 
    7.337594e-007, -2.17445e-006, -8.462573e-007, 5.971684e-007, 
    3.686841e-007, -8.673678e-007, -2.645325e-006, -5.502152e-007, 
    -4.139165e-006, -5.597729e-006, -1.093384e-005, -5.251775e-006, 
    2.116354e-006, 3.42865e-007, 1.851622e-007, -2.810222e-006, 
    -2.962959e-006, -5.65371e-007, -2.595652e-006, -1.933298e-006, 
    -1.252067e-006, -4.353989e-006, -7.908909e-006, -8.882454e-006, 
    -7.420154e-006, -4.764272e-006, -5.332249e-006, -3.108502e-006, 
    -7.49193e-006, -1.191509e-005, -1.2795e-005, -1.132301e-005, 
    -1.336025e-005, -1.286852e-005, -6.947786e-006, -9.532643e-006, 
    -1.152443e-005, -8.613242e-006, -1.0986e-005, -8.415302e-006, 
    -8.8755e-006, -3.771594e-006, -3.972764e-006, -1.102548e-005, 
    -1.128203e-005, -2.695797e-007, -2.470915e-008, -1.35687e-006, 
    -1.925104e-006, -2.598885e-006, -4.892907e-006, 2.010789e-006, 
    -4.471567e-007, -1.459193e-006, -2.16998e-006, -4.075588e-006, 
    -1.234187e-006, -1.161419e-006, -2.718092e-006, -2.756092e-006, 
    -1.19147e-006, -4.160773e-006, -3.817051e-006, -4.166982e-006, 
    -4.019461e-006, -2.314024e-006, -6.86317e-007, 5.420347e-007, 
    1.180961e-007, 8.740817e-007, 1.71128e-006, 9.339351e-007, 1.354148e-006,
  1.132866e-006, 8.147258e-007, 7.935319e-008, 5.410409e-007, 6.758963e-007, 
    5.922014e-007, 6.3467e-007, 5.067685e-007, 2.579189e-007, 1.960791e-007, 
    1.398605e-006, 1.954912e-006, 1.794974e-006, 1.367807e-006, 
    1.702587e-006, 2.240768e-006, -3.659443e-007, 9.398946e-007, 
    7.600879e-007, 3.188978e-006, 2.799312e-006, 1.118212e-006, 
    2.345572e-006, 3.742059e-006, 3.212322e-006, 1.358866e-006, 
    8.725929e-007, 6.56526e-007, 1.194456e-006, 4.385537e-006, 6.067133e-006, 
    2.087418e-007, -1.682696e-006, -8.084971e-007, -1.603734e-006, 
    -1.028042e-006, -7.417162e-006, -2.677112e-006, 5.362814e-006, 
    -3.618867e-006, -3.916146e-006, 1.061762e-007, 3.901005e-006, 
    3.103793e-006, -3.47567e-007, -5.183984e-006, -7.656833e-006, 
    -9.13503e-006, -8.334337e-006, -7.552027e-006, -6.206452e-006, 
    -4.794816e-006, -9.24356e-006, -9.688607e-006, -1.128179e-005, 
    -9.927271e-006, -2.753361e-006, -4.282792e-007, -2.307566e-006, 
    -6.897371e-006, -3.837171e-006, -3.434094e-006, -4.358959e-006, 
    -8.534016e-006, -6.51466e-006, -4.648788e-006, -8.143854e-006, 
    -9.433548e-006, -5.196725e-007, 2.993524e-006, -9.768919e-007, 
    -1.392877e-006, -9.225732e-008, -7.168601e-007, 5.390881e-006, 
    7.415199e-006, 3.718711e-006, 1.727918e-006, 1.081706e-006, 
    -6.915343e-007, -2.814451e-006, -2.79235e-006, -2.812217e-006, 
    -1.709033e-006, -2.281735e-006, -2.07362e-006, -3.365547e-006, 
    -2.886725e-006, -2.074859e-006, -6.277064e-007, -5.052686e-007, 
    -3.262064e-007, 4.210867e-007, 1.127898e-006, 1.384944e-006, 1.028061e-006,
  1.635447e-007, 2.420243e-007, 4.695155e-007, -4.690094e-007, 
    -3.803476e-007, 1.908636e-007, 3.835851e-007, 5.931948e-007, 
    4.682738e-007, 3.734031e-007, 3.654557e-007, 7.280503e-007, 
    2.091507e-006, 2.117087e-006, 2.017747e-006, 2.338618e-006, 2.98649e-007, 
    -6.632235e-007, 1.276662e-006, -9.5735e-008, 8.472603e-007, 
    3.329794e-006, 9.540513e-007, 4.498791e-006, 3.314645e-006, 
    1.210849e-006, 1.769572e-007, 1.289573e-006, 4.4218e-006, 5.929298e-006, 
    8.414067e-006, 4.517414e-006, -4.29769e-007, 8.016967e-006, 
    3.252062e-006, -1.349421e-006, -1.586839e-006, -3.899997e-006, 
    2.226116e-006, -4.595749e-007, -2.680343e-006, -3.030273e-006, 
    9.1332e-007, 2.175946e-006, 1.470873e-006, -1.649183e-006, 
    -6.020437e-006, -6.637842e-006, -5.205844e-006, -6.674596e-006, 
    -6.380549e-006, -3.405285e-006, -1.637758e-006, -1.252314e-006, 
    -2.303592e-006, -2.632163e-006, -7.363269e-008, 7.608342e-007, 
    -1.002472e-006, -2.895911e-006, -3.146252e-006, -6.162809e-007, 
    -2.914385e-007, -2.621484e-006, -3.819785e-006, -2.092741e-006, 
    5.139682e-007, -1.49297e-006, -5.385647e-006, -3.982952e-006, 
    -1.975517e-006, 4.934158e-006, 1.652923e-006, 5.85505e-006, 
    9.864456e-006, 1.102476e-005, 9.475529e-006, 7.239114e-006, 
    4.627685e-006, 8.666302e-007, -1.674265e-006, -3.03623e-006, 
    -6.196022e-006, -5.073964e-006, -1.097093e-006, -9.59757e-007, 
    -2.121051e-006, -3.05844e-007, -1.336011e-006, 1.980643e-007, 
    1.834137e-007, -1.203223e-007, 3.522932e-007, 4.176098e-007, 
    7.675387e-007, 5.445178e-007,
  1.069205e-007, 4.433571e-008, -2.387865e-007, -3.324153e-007, 
    -6.314319e-007, -5.387958e-007, -4.819243e-007, 1.680148e-007, 
    6.093383e-007, 3.724097e-007, 5.782937e-007, 3.902908e-007, 
    5.380607e-007, 1.998376e-006, 1.837691e-006, 1.372279e-006, 
    -1.934042e-006, -3.586583e-006, -2.430253e-006, -8.216698e-007, 
    -1.702577e-006, -2.709153e-006, 1.183279e-006, 1.53023e-006, 
    3.961354e-006, 7.752711e-006, 2.930688e-006, 2.977629e-006, 
    4.073114e-006, 7.956856e-006, 9.896741e-006, 6.439419e-006, 
    3.856811e-006, 3.89828e-006, 5.75844e-006, 3.719251e-007, -2.628425e-006, 
    -4.817652e-006, -2.795565e-006, 9.918076e-007, -3.410969e-007, 
    -1.412005e-006, -2.542009e-006, -3.710507e-006, -4.76998e-006, 
    -3.103785e-006, -5.003187e-006, -5.491944e-006, -5.346161e-006, 
    -7.310631e-006, -6.567059e-006, -4.896228e-007, -3.464083e-008, 
    6.289556e-007, 1.376249e-006, 3.77385e-006, 4.564852e-006, 4.435457e-006, 
    6.982464e-007, -6.393802e-007, -5.301063e-007, -2.332401e-006, 
    -1.636021e-006, -2.026183e-006, -3.235411e-006, -1.480798e-006, 
    8.673769e-007, 1.961366e-006, -2.875798e-006, -3.265712e-006, 
    -3.038567e-007, 2.579771e-006, 9.323296e-006, 1.218705e-005, 8.99e-006, 
    1.083998e-005, 1.13434e-005, 8.85018e-006, 8.960202e-006, 4.186364e-006, 
    1.684459e-006, -3.567706e-006, -6.810447e-006, -4.971644e-006, 
    -5.888562e-006, -6.161999e-006, -1.477571e-006, 2.425044e-006, 
    3.643214e-006, 2.41958e-006, 8.167099e-007, 5.16206e-007, 3.776252e-007, 
    3.565151e-007, 3.445941e-007, 2.628859e-007,
  -1.045436e-006, -6.982389e-007, -7.792016e-007, -7.195968e-007, 
    -1.588334e-006, -3.755959e-006, -2.677612e-006, -8.614061e-007, 
    -1.580638e-006, -8.814823e-009, -6.150399e-007, -3.793532e-007, 
    1.019534e-007, 4.960893e-007, 3.097084e-006, 3.933042e-006, 
    3.359096e-006, 4.086687e-007, -1.903743e-006, -2.098205e-006, 
    -2.759321e-006, -6.191552e-006, -1.783543e-006, 7.804533e-007, 
    4.541178e-007, -1.200409e-006, 2.462298e-006, 3.620863e-006, 
    2.371645e-006, 1.965098e-006, 7.316848e-006, 8.155283e-006, 
    8.951753e-006, 8.370862e-006, 7.670013e-006, 4.876543e-006, 
    4.000845e-006, -9.436044e-007, -6.146343e-006, 1.317647e-006, 
    4.232566e-006, 3.304474e-006, 1.63107e-006, -6.483097e-007, 
    -6.927658e-007, -2.633893e-006, -4.096193e-006, -2.698962e-006, 
    -2.610792e-006, -5.477279e-006, -5.527694e-006, 2.137458e-006, 
    3.128884e-006, 3.474594e-006, 5.808608e-006, 5.507354e-006, 
    4.767016e-006, 4.78067e-006, 2.729525e-006, -2.06269e-006, 
    -2.815448e-006, -2.756835e-006, -2.417089e-006, -2.630922e-006, 
    -3.143272e-006, -1.267214e-006, -7.461713e-007, -1.92098e-007, 
    -4.948406e-007, -1.12069e-006, -2.791356e-006, 8.927091e-007, 
    7.311639e-006, 1.08154e-005, 1.013292e-005, 1.06264e-005, 1.078759e-005, 
    2.723074e-006, 3.006196e-006, 4.286201e-006, 3.250076e-006, 
    2.873327e-006, -2.576031e-006, -4.708629e-006, -4.970887e-006, 
    -6.571525e-006, -5.621296e-007, 4.185869e-006, 8.414569e-006, 
    6.904089e-006, 4.868583e-006, 2.575295e-006, 2.599036e-007, 
    2.482338e-007, -6.003879e-007, -7.521312e-007,
  -2.082308e-006, -4.595888e-006, -3.949178e-006, -6.004791e-006, 
    -4.89093e-006, -6.054463e-006, -4.883976e-006, -3.227217e-006, 
    -5.595753e-006, -1.922854e-006, -4.548547e-007, 1.094022e-007, 
    1.970693e-007, 8.773086e-007, 1.021849e-006, 3.078958e-006, 4.27403e-006, 
    3.48203e-006, 1.977261e-006, 3.593044e-006, 1.368798e-006, 8.740244e-010, 
    2.661127e-007, 1.163414e-006, 1.204888e-006, 8.276397e-007, 
    8.696115e-007, 2.60982e-006, 3.662831e-006, 3.134337e-006, 4.266079e-006, 
    5.675481e-006, 5.195416e-006, 5.643451e-006, 8.845211e-006, 
    1.067706e-005, 1.144572e-005, 1.355175e-005, 9.307896e-006, 
    2.460067e-006, 3.767142e-006, 4.867346e-006, 4.356982e-006, 5.88187e-006, 
    8.611758e-006, 1.225759e-005, 1.269766e-005, 8.789844e-006, 
    4.640598e-006, 4.495327e-006, 4.423055e-006, 4.894675e-006, 
    6.575523e-006, 1.112782e-005, 1.156642e-005, 1.195956e-005, 
    1.146335e-005, 8.454805e-006, 6.542985e-006, 1.773617e-006, 2.77075e-006, 
    -9.898049e-007, -2.634397e-006, -2.755593e-006, -1.118824e-007, 
    1.406943e-007, -2.996339e-007, 1.717238e-006, 1.105545e-006, 
    2.777951e-006, 2.328929e-006, 1.814095e-006, 4.326193e-006, 
    1.166998e-005, 1.475874e-005, 1.433158e-005, 1.114025e-005, 
    9.352356e-006, 8.365896e-007, -3.998095e-006, -3.379697e-006, 
    -3.073725e-006, -3.42316e-006, -3.936751e-006, -6.750837e-006, 
    -6.302558e-006, -4.508707e-006, 6.565584e-006, 1.265221e-005, 
    1.254716e-005, 1.03167e-005, 5.621343e-006, 2.008059e-006, 
    -1.262833e-007, -2.016001e-006, -2.29639e-006,
  -5.248903e-007, -2.019227e-006, -5.062542e-006, -5.587804e-006, 
    -3.668534e-006, -4.357466e-006, -2.012275e-006, -8.505594e-008, 
    -2.424535e-006, -2.357476e-006, 2.194576e-006, 1.96435e-006, 
    2.028672e-006, 2.17942e-006, 3.467875e-006, 2.670415e-006, 2.388042e-006, 
    3.33948e-006, 4.157553e-006, 4.667418e-006, 1.808133e-006, 1.613676e-006, 
    9.67711e-007, 1.253565e-006, 1.389662e-006, 1.347442e-006, 1.058608e-006, 
    9.53306e-007, 1.051656e-006, 1.472365e-006, 2.080331e-006, 3.117205e-006, 
    3.91218e-006, 4.653761e-006, 4.067398e-006, 4.443655e-006, 1.280892e-006, 
    4.179416e-006, 7.259732e-006, 6.279737e-006, 5.304697e-006, 
    5.795941e-006, 3.39809e-006, 9.806317e-007, 2.261295e-007, 4.923975e-006, 
    8.517884e-006, 9.505085e-006, 1.071059e-005, 9.274612e-006, 
    6.439921e-006, 1.117426e-005, 1.087425e-005, 9.572388e-006, 1.18915e-005, 
    1.568585e-005, 1.643511e-005, 1.497208e-005, 1.194491e-005, 
    9.476284e-006, 5.263479e-006, 3.16216e-006, 8.204443e-007, 
    -1.726159e-006, -6.882947e-007, 7.633153e-007, 1.309198e-006, 
    6.473338e-007, 1.500176e-006, 3.519036e-006, 6.538009e-006, 
    6.002565e-006, 6.769729e-006, 1.014683e-005, 1.362277e-005, 
    1.856127e-005, 1.857691e-005, 1.684068e-005, 1.147875e-005, 
    6.651513e-006, 3.545356e-007, -3.363552e-006, -5.530175e-006, 
    -2.642082e-006, -5.589784e-006, -9.571373e-006, -8.177372e-006, 
    -3.799159e-006, 5.424412e-006, 9.342912e-006, 1.375912e-005, 
    1.06187e-005, 4.851949e-006, 2.212952e-006, -1.043451e-006, -2.434721e-006,
  3.23964e-006, 9.689484e-007, 3.475725e-007, -2.350644e-007, -6.657065e-007, 
    -1.589824e-006, 3.244364e-006, 3.112733e-006, 5.057579e-006, 
    4.175683e-006, 3.920128e-006, 5.985679e-006, 3.998852e-006, 
    3.640231e-006, 3.139056e-006, 2.273301e-006, 3.14055e-006, 3.838421e-006, 
    4.573295e-006, 5.366286e-006, 4.544239e-006, 2.180914e-006, 
    1.454979e-006, 9.113352e-007, 4.831747e-007, 5.109901e-007, 7.98831e-007, 
    7.491603e-007, 6.955162e-007, 6.232456e-007, 5.805292e-007, 8.48005e-007, 
    1.259774e-006, 1.2784e-006, 1.934796e-006, 2.365441e-006, 1.952676e-006, 
    -4.126305e-007, 3.148001e-006, 5.5898e-006, 7.088867e-006, 5.241371e-006, 
    4.334888e-006, 3.804649e-006, 2.782675e-006, 4.831891e-007, 
    -3.733949e-007, -1.612432e-006, 1.334774e-006, 3.22624e-006, 
    8.087991e-006, 6.981085e-006, 9.574876e-006, 8.467468e-006, 
    5.581613e-006, 4.716603e-006, 6.844231e-006, 1.166204e-005, 
    1.508781e-005, 9.527939e-006, 8.823368e-006, 7.366772e-006, 
    4.278259e-006, 5.942216e-006, 5.526985e-006, 2.198805e-006, 
    2.404184e-006, 3.071007e-006, 4.743414e-006, 4.201262e-006, 
    5.464382e-006, 8.894629e-006, 7.746747e-006, 7.266679e-006, 
    1.112558e-005, 1.415747e-005, 1.332226e-005, 1.362725e-005, 1.13501e-005, 
    6.991268e-006, 6.48413e-006, 3.300251e-006, 2.83161e-006, -4.632857e-007, 
    -2.11806e-006, -3.067518e-006, -3.125635e-006, -1.549088e-006, 
    4.398215e-006, 5.92757e-006, 9.531661e-006, 8.88644e-006, 7.330258e-006, 
    1.004973e-006, -2.42627e-006, -7.983908e-008,
  -4.16723e-006, -1.940252e-006, 6.063583e-007, 2.942115e-006, 4.58338e-007, 
    3.200897e-006, 3.33203e-006, 1.920142e-006, 1.613178e-006, 2.397228e-006, 
    2.673891e-006, 3.451978e-006, 3.117699e-006, 3.846116e-006, 
    5.833186e-006, 4.496306e-006, 3.989419e-006, 3.746531e-006, 
    3.731878e-006, 3.127883e-006, 3.711761e-006, 3.265472e-006, 
    2.198548e-006, 1.453489e-006, 1.081953e-006, 1.522531e-006, 
    1.633545e-006, 6.185269e-007, 5.181923e-007, 7.081824e-007, 
    7.061957e-007, 7.543758e-007, 5.301134e-007, 6.006455e-007, 1.14727e-006, 
    1.018872e-006, 1.391153e-006, 8.457673e-007, -3.155292e-007, 
    -1.039225e-007, -6.145638e-008, 1.307959e-006, 2.54302e-006, 
    3.857058e-006, 3.434609e-006, 3.843648e-006, 4.392008e-006, 
    7.464405e-008, 2.214201e-006, 2.512224e-006, 2.14715e-006, 4.753609e-006, 
    5.958616e-006, 7.601713e-006, 9.854772e-006, 5.854054e-006, 
    1.593318e-006, 4.764777e-006, 6.068636e-006, 7.162129e-006, 
    8.683044e-006, 8.220362e-006, 7.221483e-006, 9.13057e-006, 9.741278e-006, 
    7.305436e-006, 5.0402e-006, 4.497543e-006, 3.968554e-006, 4.525114e-006, 
    4.758316e-006, 6.324428e-006, 8.788582e-006, 9.521473e-006, 1.01965e-005, 
    1.164042e-005, 1.367542e-005, 1.398288e-005, 1.119563e-005, 
    7.576135e-006, 6.645059e-006, 4.248461e-006, 3.189485e-006, 
    3.925852e-006, 2.655775e-006, 3.703823e-006, -1.083423e-006, 
    3.479563e-006, 3.439574e-006, 2.103934e-006, 2.832348e-006, 
    6.212686e-006, 4.823152e-006, 1.611195e-006, -2.914312e-007, 
    -4.224592e-006,
  -2.464276e-006, -8.882271e-007, 1.447283e-006, 4.77645e-006, 4.755833e-006, 
    3.297755e-006, 1.878916e-006, 1.491981e-006, 2.181408e-006, 
    3.547846e-006, 2.993273e-006, 1.54786e-006, 1.990177e-006, 1.877425e-006, 
    3.65389e-006, 4.709887e-006, 3.454963e-006, 3.3365e-006, 3.960113e-006, 
    3.088644e-006, 1.542399e-006, 1.811864e-006, 3.378223e-006, 
    3.549337e-006, 1.735618e-006, 1.327823e-006, 1.249094e-006, 
    1.127899e-006, 9.237526e-007, 5.561906e-007, 5.18193e-007, 2.301033e-007, 
    2.924398e-007, 5.316037e-007, 2.243917e-007, 5.750653e-007, 
    7.958513e-007, -2.91685e-007, -1.14627e-006, -1.679979e-006, 
    -9.046198e-007, 9.744163e-007, 5.894726e-007, 7.402195e-007, 
    9.42382e-007, 1.830991e-006, 3.349178e-006, 1.685708e-006, 5.884107e-006, 
    7.541363e-006, 5.430124e-006, 4.553687e-006, 7.96431e-006, 4.553931e-006, 
    8.658462e-006, 1.158927e-005, 9.124124e-006, 5.233182e-006, 
    5.642461e-006, 4.809488e-006, 3.167872e-006, 5.422422e-006, 
    5.805625e-006, 8.65473e-006, 1.015479e-005, 6.631644e-006, 4.235782e-006, 
    2.925223e-006, 2.32322e-006, 3.062067e-006, 2.061206e-006, 1.157699e-006, 
    2.609071e-006, 6.846215e-006, 6.991502e-006, 7.931771e-006, 
    9.306901e-006, 9.689364e-006, 9.74574e-006, 9.889287e-006, 7.401788e-006, 
    3.070272e-006, 1.909721e-006, 5.993879e-006, 6.868326e-006, 
    3.031531e-006, -8.437637e-007, -1.568456e-006, -2.904599e-006, 
    -2.722802e-006, -1.107517e-006, 2.960998e-006, 4.000853e-006, 
    2.735989e-006, -3.669302e-007, -1.312656e-006,
  2.403689e-006, 8.797961e-007, 4.918638e-007, 1.196195e-006, 1.1423e-006, 
    5.519687e-007, 7.908839e-007, 1.59579e-006, 3.192452e-006, 4.339343e-006, 
    3.638243e-006, 2.981351e-006, 4.071619e-006, 3.930803e-006, 
    3.689654e-006, 4.014499e-006, 3.351398e-006, 2.734245e-006, 
    2.518922e-006, 2.84948e-006, 2.515198e-006, 1.958142e-006, 2.774475e-006, 
    2.799808e-006, 1.456219e-006, 1.305223e-006, 1.648446e-006, 
    1.037748e-006, 4.034541e-007, 1.019866e-006, 1.004468e-006, 
    1.106293e-006, 7.362462e-007, 6.893076e-007, 1.135846e-006, 
    9.011528e-007, 6.339255e-007, -3.639561e-007, -5.345773e-007, 
    2.40617e-006, 5.244001e-007, 1.612681e-006, 9.463492e-007, 3.632194e-007, 
    8.149727e-007, 1.526514e-006, 1.681481e-006, 4.934152e-006, 
    4.471225e-006, 4.939873e-006, 4.991769e-006, 6.814433e-006, 
    5.196918e-006, 4.959988e-006, 6.361199e-006, 6.142149e-006, 
    7.040941e-006, 7.674735e-006, 4.524132e-006, 3.293539e-006, 
    3.531211e-006, 5.001457e-006, 7.575632e-006, 6.985054e-006, 
    4.945829e-006, 5.049384e-006, 4.772472e-006, 2.494332e-006, 
    2.120313e-006, 1.866e-006, 1.244869e-006, 1.807637e-006, 1.877673e-006, 
    2.159802e-006, 3.467129e-006, 5.8158e-006, 6.86286e-006, 6.28395e-006, 
    6.270287e-006, 6.98033e-006, 4.346301e-006, 9.97019e-007, 2.558663e-006, 
    5.40751e-006, 5.035228e-006, 6.417071e-006, 4.457575e-006, 5.152215e-007, 
    -3.276626e-006, -7.145714e-006, -5.627786e-006, -5.504626e-007, 
    -1.75025e-006, 1.674038e-006, 3.859284e-006, 2.857425e-006,
  1.193959e-006, 3.740079e-006, 5.940979e-006, 3.93156e-006, 4.228334e-006, 
    3.004203e-006, 8.30617e-007, 8.085135e-007, 2.809495e-006, 1.848864e-006, 
    8.800407e-007, 2.845751e-006, 3.70058e-006, 3.116705e-006, 7.446888e-007, 
    1.832223e-006, 2.414362e-006, 2.332657e-006, 2.403935e-006, 2.33241e-006, 
    2.225121e-006, 1.723448e-006, 1.510113e-006, 1.298268e-006, 
    1.875937e-006, 1.998621e-006, 2.090263e-006, 1.715749e-006, 
    9.823643e-007, 1.221028e-006, 1.166142e-006, 1.694889e-006, 
    1.547367e-006, 2.072882e-006, 2.827128e-006, 1.749775e-006, 
    8.167128e-007, 1.665253e-007, -6.654582e-007, -7.024628e-007, 
    -2.8672e-007, 1.419958e-006, 2.098458e-006, 2.406911e-006, 1.835702e-006, 
    1.176079e-006, 1.371531e-006, 2.377858e-006, 4.553176e-006, 
    4.054986e-006, 2.289196e-006, 3.954403e-006, 6.38975e-006, 7.492436e-006, 
    8.017205e-006, 9.08388e-006, 1.072599e-005, 1.01965e-005, 9.562955e-006, 
    1.09813e-005, 1.142163e-005, 1.299668e-005, 7.464125e-006, 2.672405e-006, 
    2.638126e-006, 2.907591e-006, 2.081822e-006, 1.173343e-006, 
    1.045939e-006, 1.013157e-006, 1.633542e-006, 1.649685e-006, 
    3.650413e-006, 6.30282e-006, 7.32057e-006, 6.776178e-006, 4.77694e-006, 
    1.929826e-006, 2.9215e-006, 5.353118e-006, 5.734591e-006, 6.211183e-006, 
    5.101792e-006, 5.116444e-006, 3.760688e-006, 1.470627e-006, 
    -5.134643e-007, 1.998051e-007, -1.374992e-006, -3.378707e-006, 
    -1.303717e-006, 3.047175e-006, 5.023569e-006, 2.893197e-006, 
    1.059605e-006, 5.55694e-007,
  3.20885e-006, 3.812351e-006, 2.541776e-006, 2.608329e-006, 2.428522e-006, 
    2.11758e-006, 1.632052e-006, 2.642597e-006, 4.485377e-006, 3.586338e-006, 
    1.555558e-006, 1.587596e-006, 4.193809e-006, 4.268812e-006, 
    3.212568e-006, 2.346562e-006, 2.656508e-006, 3.014632e-006, 
    2.409397e-006, 2.194325e-006, 2.136707e-006, 2.346562e-006, 
    1.564003e-006, 2.200783e-006, 2.570329e-006, 2.101687e-006, 
    1.463171e-006, 1.510611e-006, 1.858552e-006, 2.218415e-006, 
    2.503028e-006, 1.34198e-006, 1.148761e-006, 1.601259e-006, 2.238035e-006, 
    1.453986e-006, 6.413759e-007, 7.054507e-007, 1.059354e-006, 
    1.482299e-006, 1.574932e-006, 1.850357e-006, 2.062201e-006, 2.78441e-006, 
    3.88635e-006, 4.14091e-006, 3.492213e-006, 2.635148e-006, 3.529467e-006, 
    3.867724e-006, 4.710882e-006, 5.466616e-006, 5.924579e-006, 
    6.466981e-006, 6.635117e-006, 1.050222e-005, 1.501951e-005, 1.66862e-005, 
    1.082955e-005, 9.5041e-006, 7.282828e-006, 4.815936e-006, 4.305817e-006, 
    3.178296e-006, 1.623359e-006, 1.433621e-006, 2.229591e-006, 
    2.035874e-006, 1.577166e-006, 1.774855e-006, 1.879661e-006, 
    2.724558e-006, 3.83221e-006, 5.256761e-006, 5.006422e-006, 3.976255e-006, 
    4.255651e-006, 3.759194e-006, 3.54561e-006, 5.833433e-006, 8.220103e-006, 
    8.564071e-006, 6.714339e-006, 7.7609e-006, 9.127096e-006, 5.098071e-006, 
    -1.83544e-006, -2.571309e-006, -3.388883e-006, -2.219145e-006, 
    9.153118e-007, 1.537683e-006, 2.934357e-007, 1.246121e-006, 
    2.287215e-006, 2.822166e-006,
  -1.04717e-006, -1.133598e-006, 6.823557e-007, 1.746794e-006, 1.869976e-006, 
    9.793839e-007, 1.122185e-006, 2.056737e-006, 2.350786e-006, 
    1.424429e-006, 1.34297e-006, 9.813684e-007, 1.601257e-006, 1.674521e-006, 
    1.946218e-006, 1.855321e-006, 1.566735e-006, 1.458701e-006, 
    1.652914e-006, 1.771875e-006, 2.108395e-006, 1.915174e-006, 
    1.663345e-006, 1.599517e-006, 2.216177e-006, 3.197666e-006, 
    3.594785e-006, 1.916418e-006, 1.401584e-006, 1.831482e-006, 
    1.818817e-006, 1.865259e-006, 1.868239e-006, 2.073875e-006, 
    1.745304e-006, 1.367062e-006, 1.345953e-006, 1.439084e-006, 
    1.805653e-006, 2.583246e-006, 4.022202e-006, 4.003326e-006, 
    3.203133e-006, 3.135333e-006, 2.475461e-006, 2.607833e-006, 
    4.072615e-006, 5.29004e-006, 5.605199e-006, 5.964564e-006, 6.704158e-006, 
    5.430111e-006, 5.220253e-006, 5.101044e-006, 5.646177e-006, 
    5.804874e-006, 6.513425e-006, 6.339576e-006, 6.174175e-006, 
    5.288301e-006, 3.932544e-006, 2.892941e-006, 2.271811e-006, 
    1.838684e-006, 1.93728e-006, 2.544252e-006, 2.913055e-006, 1.627336e-006, 
    1.070778e-006, 1.298766e-006, 1.0298e-006, 8.894808e-007, 1.223763e-006, 
    1.316399e-006, 1.181543e-006, 1.27567e-006, 1.830738e-006, 3.61391e-006, 
    4.863867e-006, 5.831449e-006, 7.324298e-006, 8.797524e-006, 
    9.051339e-006, 1.053376e-005, 1.121127e-005, 6.578754e-006, 
    1.372355e-007, 6.657247e-007, 6.408125e-006, 4.449874e-006, 
    -6.281989e-007, -3.463399e-006, -1.707793e-006, 6.870741e-007, 
    1.036915e-007, 8.456846e-008,
  -2.209717e-006, -4.626185e-006, -4.621215e-006, -2.086033e-006, 
    2.149536e-007, 1.642977e-006, 2.657252e-006, 3.562746e-006, 
    2.563623e-006, 9.667165e-007, 3.279529e-007, 4.33005e-007, 9.118303e-007, 
    2.242752e-006, 2.799308e-006, 2.282984e-006, 2.004581e-006, 
    1.405556e-006, 1.594057e-006, 1.925608e-006, 2.459316e-006, 2.52364e-006, 
    2.087779e-006, 1.684453e-006, 2.212948e-006, 2.126025e-006, 
    1.940261e-006, 1.286099e-006, 1.221279e-006, 1.357874e-006, 
    1.048179e-006, 1.635781e-006, 2.144407e-006, 2.265603e-006, 
    2.265602e-006, 2.122799e-006, 2.24499e-006, 2.527118e-006, 2.554437e-006, 
    2.292674e-006, 1.962364e-006, 1.76716e-006, 2.017003e-006, 1.400343e-006, 
    1.52129e-006, 2.101194e-006, 2.699723e-006, 2.974155e-006, 3.463159e-006, 
    4.479417e-006, 5.191445e-006, 4.608315e-006, 3.772608e-006, 
    3.178796e-006, 2.88102e-006, 2.331416e-006, 2.147138e-006, 1.790255e-006, 
    9.888208e-007, 9.185369e-007, 1.484037e-006, 2.548973e-006, 2.33092e-006, 
    1.920394e-006, 1.605978e-006, 1.918903e-006, 1.992167e-006, 1.37824e-006, 
    1.679739e-006, 1.452745e-006, 1.335522e-006, 1.08568e-006, 6.423693e-007, 
    6.582641e-007, 1.044205e-006, 9.036366e-007, 1.561275e-006, 
    2.703698e-006, 2.943358e-006, 3.261248e-006, 3.374497e-006, 
    3.828983e-006, 6.078065e-006, 6.876518e-006, 5.27638e-006, 4.165498e-006, 
    5.244589e-006, 6.472697e-006, 6.622706e-006, 6.275754e-006, 
    5.502383e-006, 4.166999e-006, 2.976636e-006, 2.572569e-006, 
    1.900025e-006, 3.520454e-007,
  1.565491e-006, 2.378019e-007, -2.64011e-006, -5.250542e-006, 
    -4.961461e-006, -1.27591e-006, 8.991665e-007, 1.526005e-006, 
    2.587217e-006, 3.155696e-006, 2.719587e-006, 1.549102e-006, 
    1.591322e-006, 2.423551e-006, 2.343831e-006, 2.267835e-006, 
    2.077845e-006, 1.68098e-006, 1.164903e-006, 9.076102e-007, 1.304478e-006, 
    1.390159e-006, 1.370539e-006, 1.13212e-006, 1.52104e-006, 1.693398e-006, 
    1.979252e-006, 1.702339e-006, 1.262507e-006, 1.210103e-006, 
    1.407296e-006, 1.616408e-006, 1.761198e-006, 1.955658e-006, 
    1.800438e-006, 1.439333e-006, 1.283616e-006, 1.192719e-006, 
    1.275171e-006, 1.482049e-006, 1.490742e-006, 1.331051e-006, 
    1.641989e-006, 1.814097e-006, 1.680235e-006, 1.294047e-006, 
    1.401335e-006, 1.640003e-006, 1.886617e-006, 1.681975e-006, 
    1.434616e-006, 1.128645e-006, 1.15944e-006, 1.368056e-006, 1.29678e-006, 
    1.510611e-006, 1.899779e-006, 1.776348e-006, 1.658381e-006, 1.33602e-006, 
    1.116724e-006, 1.966089e-006, 2.81322e-006, 2.527615e-006, 2.256911e-006, 
    1.604736e-006, 9.962719e-007, 9.463533e-007, 1.059105e-006, 
    1.336764e-006, 1.472861e-006, 1.322856e-006, 1.081705e-006, 
    7.215936e-007, 2.956695e-007, 4.096642e-007, 1.273683e-006, 
    1.642487e-006, 1.64199e-006, 1.614919e-006, 1.568476e-006, 1.90425e-006, 
    2.117584e-006, 1.752506e-006, 1.332543e-006, 1.142303e-006, 
    1.428157e-006, 2.842774e-006, 4.491587e-006, 5.18573e-006, 5.254523e-006, 
    5.480525e-006, 5.7408e-006, 3.823021e-006, 1.378734e-006, 1.389908e-006,
  1.051401e-006, 5.59914e-007, 1.106418e-007, -5.600123e-008, 4.429385e-007, 
    1.582877e-006, 2.649056e-006, 3.39312e-006, 3.635512e-006, 3.146507e-006, 
    2.273796e-006, 1.669056e-006, 1.485525e-006, 1.698364e-006, 2.2358e-006, 
    2.759326e-006, 2.802541e-006, 2.453606e-006, 1.870225e-006, 
    1.468391e-006, 1.27244e-006, 1.294543e-006, 1.560529e-006, 1.882642e-006, 
    1.85284e-006, 1.869232e-006, 1.997134e-006, 1.959633e-006, 1.745055e-006, 
    1.382212e-006, 1.099338e-006, 9.480912e-007, 1.117716e-006, 
    1.246114e-006, 1.360108e-006, 1.440078e-006, 1.358122e-006, 
    1.259277e-006, 1.099338e-006, 9.639855e-007, 1.173844e-006, 
    1.602501e-006, 1.858305e-006, 1.927595e-006, 1.759956e-006, 
    1.609455e-006, 1.677255e-006, 1.942495e-006, 2.070645e-006, 
    2.231578e-006, 2.051523e-006, 1.80168e-006, 1.677503e-006, 1.651426e-006, 
    1.674026e-006, 1.45473e-006, 1.174838e-006, 1.014402e-006, 1.064072e-006, 
    9.160542e-007, 1.006206e-006, 1.555313e-006, 2.002598e-006, 
    2.087534e-006, 1.838436e-006, 1.583377e-006, 1.284609e-006, 
    9.769001e-007, 8.929574e-007, 9.734235e-007, 1.426171e-006, 
    1.861285e-006, 1.765917e-006, 1.465907e-006, 1.069287e-006, 
    5.810259e-007, 2.278684e-007, 2.112297e-007, 4.223298e-007, 
    3.865666e-007, 3.480723e-007, 4.70759e-007, 6.947721e-007, 6.818573e-007, 
    5.00311e-007, 5.889733e-007, 9.883245e-007, 1.500676e-006, 2.290439e-006, 
    2.83582e-006, 2.905358e-006, 3.105281e-006, 4.372376e-006, 5.602466e-006, 
    4.473455e-006, 2.294408e-006,
  4.831081e-006, 4.604583e-006, 4.259871e-006, 3.851333e-006, 3.48973e-006, 
    3.411997e-006, 3.402561e-006, 3.229459e-006, 2.871086e-006, 
    2.377858e-006, 2.111374e-006, 2.023706e-006, 2.041339e-006, 
    2.132485e-006, 2.151608e-006, 2.009054e-006, 1.882891e-006, 1.86799e-006, 
    2.010794e-006, 2.103926e-006, 1.871964e-006, 1.581888e-006, 
    1.404813e-006, 1.404068e-006, 1.555563e-006, 1.690418e-006, 
    1.686196e-006, 1.590828e-006, 1.393388e-006, 1.093378e-006, 
    8.902255e-007, 8.313655e-007, 8.482534e-007, 9.503262e-007, 
    1.076738e-006, 1.169871e-006, 1.178563e-006, 1.169622e-006, 
    1.156707e-006, 1.170615e-006, 1.285851e-006, 1.404315e-006, 
    1.435111e-006, 1.54985e-006, 1.903504e-006, 2.336631e-006, 2.515445e-006, 
    2.384066e-006, 2.093742e-006, 1.789014e-006, 1.57394e-006, 1.660864e-006, 
    1.703332e-006, 1.455724e-006, 1.169125e-006, 1.105298e-006, 
    1.339744e-006, 1.621624e-006, 1.745551e-006, 1.850357e-006, 
    2.084057e-006, 2.22512e-006, 2.30062e-006, 2.116591e-006, 1.696875e-006, 
    1.39761e-006, 1.233697e-006, 1.023343e-006, 8.447767e-007, 6.878181e-007, 
    5.010568e-007, 5.549489e-007, 6.855826e-007, 7.099213e-007, 
    7.238284e-007, 7.337626e-007, 6.028811e-007, 2.867282e-007, -4.7306e-008, 
    -1.630385e-007, 5.344418e-009, 2.469915e-007, 4.243152e-007, 
    5.077618e-007, 5.137224e-007, 6.304479e-007, 1.15025e-006, 2.006819e-006, 
    2.880525e-006, 3.667057e-006, 4.322212e-006, 4.701943e-006, 
    4.836797e-006, 4.89491e-006, 4.914033e-006, 4.883485e-006,
  3.288567e-006, 3.218532e-006, 3.369033e-006, 3.542633e-006, 3.57318e-006, 
    3.44205e-006, 3.240387e-006, 3.044437e-006, 2.91579e-006, 2.834578e-006, 
    2.783666e-006, 2.744178e-006, 2.699475e-006, 2.656759e-006, 
    2.620251e-006, 2.574057e-006, 2.551954e-006, 2.61578e-006, 2.744675e-006, 
    2.826135e-006, 2.806515e-006, 2.642602e-006, 2.351284e-006, 
    2.001604e-006, 1.652172e-006, 1.391898e-006, 1.199673e-006, 
    1.018126e-006, 8.278885e-007, 6.513101e-007, 5.189381e-007, 
    4.096628e-007, 3.686846e-007, 3.530381e-007, 3.696773e-007, 
    4.645481e-007, 6.398859e-007, 8.360846e-007, 1.018127e-006, 
    1.174092e-006, 1.283119e-006, 1.379232e-006, 1.50912e-006, 1.642982e-006, 
    1.768896e-006, 1.903007e-006, 2.018242e-006, 2.057482e-006, 
    1.981983e-006, 1.780073e-006, 1.48056e-006, 1.179556e-006, 9.756586e-007, 
    9.197788e-007, 9.65724e-007, 1.029551e-006, 1.146773e-006, 1.214077e-006, 
    1.228481e-006, 1.245369e-006, 1.288086e-006, 1.365324e-006, 
    1.466652e-006, 1.544138e-006, 1.575678e-006, 1.585861e-006, 
    1.605977e-006, 1.579652e-006, 1.455724e-006, 1.275668e-006, 
    1.142303e-006, 1.08245e-006, 1.081457e-006, 1.090398e-006, 1.09437e-006, 
    1.084685e-006, 1.070529e-006, 1.071274e-006, 1.14578e-006, 1.244376e-006, 
    1.287589e-006, 1.311679e-006, 1.354148e-006, 1.414497e-006, 
    1.539916e-006, 1.806894e-006, 2.272308e-006, 2.882013e-006, 
    3.596773e-006, 4.283717e-006, 4.814943e-006, 5.070498e-006, 
    5.041939e-006, 4.760306e-006, 4.276018e-006, 3.690154e-006,
  1.847626e-006, 1.860292e-006, 1.866997e-006, 1.863769e-006, 1.864266e-006, 
    1.866749e-006, 1.864017e-006, 1.85756e-006, 1.834712e-006, 1.802922e-006, 
    1.76691e-006, 1.733383e-006, 1.706064e-006, 1.68719e-006, 1.683961e-006, 
    1.689922e-006, 1.700104e-006, 1.71426e-006, 1.740088e-006, 1.776348e-006, 
    1.814842e-006, 1.843651e-006, 1.85284e-006, 1.836946e-006, 1.800438e-006, 
    1.75176e-006, 1.699359e-006, 1.643231e-006, 1.584372e-006, 1.535446e-006, 
    1.50614e-006, 1.497944e-006, 1.514087e-006, 1.541158e-006, 1.572698e-006, 
    1.616408e-006, 1.661608e-006, 1.702586e-006, 1.736362e-006, 
    1.761695e-006, 1.773119e-006, 1.768649e-006, 1.750022e-006, 
    1.718233e-006, 1.68098e-006, 1.640499e-006, 1.607468e-006, 1.593063e-006, 
    1.594801e-006, 1.606723e-006, 1.617402e-006, 1.619389e-006, 
    1.605481e-006, 1.57692e-006, 1.538674e-006, 1.504153e-006, 1.482298e-006, 
    1.479566e-006, 1.498441e-006, 1.534949e-006, 1.582384e-006, 
    1.629322e-006, 1.67651e-006, 1.716743e-006, 1.748284e-006, 1.772374e-006, 
    1.810123e-006, 1.866003e-006, 1.944482e-006, 2.042582e-006, 
    2.144903e-006, 2.240519e-006, 2.327442e-006, 2.407909e-006, 
    2.475212e-006, 2.50725e-006, 2.503027e-006, 2.473474e-006, 2.426535e-006, 
    2.366186e-006, 2.300124e-006, 2.240271e-006, 2.189111e-006, 
    2.155086e-006, 2.141427e-006, 2.140433e-006, 2.141675e-006, 
    2.127023e-006, 2.098462e-006, 2.063444e-006, 2.01601e-006, 1.959882e-006, 
    1.913688e-006, 1.878918e-006, 1.853586e-006, 1.841169e-006 ;
}
