netcdf CGMR_SRA1B_1_tas-change_2070-2099 {
dimensions:
	time = 12 ;
	latitude = 48 ;
	longitude = 96 ;
	bounds = 2 ;
data:
 air_temperature_anomaly =
  2.341751, 2.305161, 2.272995, 2.248322, 2.232758, 2.22937, 2.234711, 
    2.246628, 2.270981, 2.295395, 2.327682, 2.360825, 2.396698, 2.433167, 
    2.464066, 2.49025, 2.510361, 2.521103, 2.529373, 2.5271, 2.509796, 
    2.497726, 2.471695, 2.446182, 2.418121, 2.392929, 2.36525, 2.337982, 
    2.310486, 2.281723, 2.250854, 2.214218, 2.175537, 2.136139, 2.101257, 
    2.067993, 2.04129, 2.018387, 2.001053, 1.983597, 1.970978, 1.957123, 
    1.9534, 1.964996, 1.969162, 1.9646, 1.949036, 1.959259, 1.962585, 
    1.960754, 1.946701, 1.941498, 1.961288, 1.914093, 1.943893, 1.944931, 
    1.953278, 1.958023, 1.972595, 2.005753, 2.032318, 2.055222, 2.1064, 
    2.153595, 2.212524, 2.284195, 2.339539, 2.390961, 2.433609, 2.459198, 
    2.48764, 2.504898, 2.517654, 2.52652, 2.544556, 2.556396, 2.570511, 
    2.599365, 2.614136, 2.631271, 2.644424, 2.660172, 2.672424, 2.67717, 
    2.671692, 2.668442, 2.655289, 2.637985, 2.615967, 2.585693, 2.55835, 
    2.53009, 2.49826, 2.459854, 2.418564, 2.379196,
  2.211731, 2.176895, 2.170517, 2.177292, 2.172028, 2.171829, 2.16864, 
    2.14859, 2.112244, 2.066483, 2.028854, 1.999237, 1.990128, 2.010498, 
    2.059647, 2.123642, 2.194672, 2.265442, 2.328461, 2.365311, 2.383148, 
    2.395004, 2.391617, 2.387329, 2.382828, 2.360565, 2.339218, 2.28804, 
    2.242599, 2.18895, 2.144669, 2.114471, 2.114532, 2.109909, 2.102692, 
    2.102814, 2.116745, 2.130539, 2.145325, 2.157043, 2.171204, 2.189606, 
    2.214355, 2.204254, 2.184784, 2.182404, 2.157501, 2.180176, 2.203033, 
    2.244324, 2.265839, 2.263702, 2.32132, 2.327698, 2.412598, 2.28479, 
    2.242157, 2.262665, 2.257141, 2.288116, 2.283752, 2.336761, 2.353729, 
    2.390015, 2.443848, 2.498871, 2.508026, 2.546265, 2.61203, 2.676086, 
    2.717361, 2.726974, 2.717484, 2.757721, 2.774109, 2.764557, 2.757111, 
    2.750092, 2.778473, 2.775757, 2.773651, 2.79953, 2.809601, 2.827576, 
    2.851532, 2.869202, 2.857208, 2.839172, 2.845673, 2.795166, 2.727829, 
    2.649765, 2.556519, 2.461151, 2.365387, 2.275665,
  2.258743, 2.17598, 2.13147, 2.102615, 2.131332, 2.198318, 2.217133, 
    2.190186, 2.230286, 2.271103, 2.311417, 2.369156, 2.466095, 2.585693, 
    2.62645, 2.618317, 2.597733, 2.593765, 2.579498, 2.554962, 2.510376, 
    2.479309, 2.417587, 2.323334, 2.248657, 2.187454, 2.197998, 2.250992, 
    2.293762, 2.332764, 2.3396, 2.315323, 2.292725, 2.274231, 2.271301, 
    2.261673, 2.267456, 2.2883, 2.313004, 2.33017, 2.322693, 2.338379, 
    2.331482, 2.324646, 2.335968, 2.318726, 2.333099, 2.347778, 2.276093, 
    2.14209, 2.010834, 1.927185, 1.915894, 1.922638, 1.914368, 1.976288, 
    2.1073, 2.15271, 2.254456, 2.348541, 2.482269, 2.574951, 2.605164, 
    2.742523, 2.848846, 2.91156, 2.879578, 2.807907, 2.701584, 2.682449, 
    2.754715, 2.815002, 2.811829, 2.773865, 2.764496, 2.733063, 2.73349, 
    2.711609, 2.625946, 2.596191, 2.533478, 2.426086, 2.346466, 2.303497, 
    2.318085, 2.372284, 2.408112, 2.408875, 2.435974, 2.451721, 2.470215, 
    2.50116, 2.533417, 2.492844, 2.459854, 2.376328,
  2.482895, 2.275284, 2.06752, 1.915833, 1.868973, 1.953735, 2.103729, 
    2.187714, 2.179642, 2.136078, 2.141556, 2.125473, 2.147736, 2.219803, 
    2.286148, 2.312912, 2.307312, 2.369537, 2.385818, 2.338547, 2.306473, 
    2.278931, 2.284851, 2.218643, 2.094864, 1.987778, 1.912262, 1.944611, 
    2.047531, 2.117996, 2.121628, 2.156921, 2.25737, 2.313293, 2.266235, 
    2.179321, 2.129639, 2.130676, 2.129578, 2.145386, 2.204712, 2.221252, 
    2.221527, 2.192993, 2.113068, 1.994904, 1.082855, 0.8957825, 0.9254761, 
    0.979187, 1.030334, 1.028625, 0.9282837, 0.8403931, 0.8907166, 0.920929, 
    0.9367676, 1.538055, 1.780518, 1.947296, 2.169678, 2.401764, 2.559082, 
    2.596924, 2.53891, 2.380249, 2.347595, 2.415009, 2.474976, 2.483826, 
    2.42627, 2.312988, 2.212708, 2.100311, 2.024292, 2.009735, 1.987274, 
    2.043915, 2.115265, 2.119812, 1.706421, 1.72229, 1.69632, 1.618073, 
    1.701569, 1.743469, 1.74176, 1.762024, 1.71344, 2.479156, 2.511169, 
    2.549591, 2.581879, 2.608307, 2.618515, 2.574173,
  2.321777, 2.244568, 2.188782, 2.225784, 2.304077, 2.260178, 2.171768, 
    2.087784, 2.053345, 1.97348, 1.89827, 1.883774, 1.831192, 1.875412, 
    2.066544, 2.216476, 2.220596, 2.21611, 2.156097, 2.112274, 2.05426, 
    2.03688, 1.95816, 1.8004, 1.632507, 1.546768, 1.549744, 1.703796, 
    1.774307, 1.828018, 1.835434, 1.83374, 1.917786, 2.050659, 2.171432, 
    2.239471, 2.289795, 2.465378, 2.488953, 2.391617, 2.307846, 2.267563, 
    2.234131, 2.146454, 2.013885, 1.90863, 1.084656, 0.8503113, 0.6000366, 
    0.4362488, 0.3918152, 0.3330383, 0.2655334, 0.2478943, 0.32547, 
    0.4508972, 0.5824585, 0.6856995, 0.825531, 0.9524231, 1.049591, 1.060059, 
    1.004211, 0.8954163, 0.8186646, 0.7725525, 0.6322021, 0.5087585, 
    0.5269775, 0.6066895, 1.415649, 1.110321, 1.041443, 0.8077087, 0.5775146, 
    0.474762, 1.109802, 1.086151, 1.174744, 1.28598, 1.219696, 1.23584, 
    1.239868, 1.225494, 1.231354, 1.202942, 1.191437, 1.240387, 1.335449, 
    1.398224, 1.527374, 2.003601, 2.12146, 2.212067, 2.240509, 2.262024,
  1.047119, 0.9476318, 1.606537, 1.612274, 1.705048, 1.668243, 1.60199, 
    1.599426, 1.673462, 1.640137, 1.783325, 1.895935, 1.838898, 1.742065, 
    1.673462, 1.81897, 1.74353, 1.591827, 1.404388, 1.328949, 1.360321, 
    1.378143, 1.340149, 1.509613, 1.616699, 1.654083, 1.61441, 1.594177, 
    1.672699, 1.698975, 1.663177, 1.514618, 1.47467, 1.501129, 1.52594, 
    1.43631, 1.34079, 1.340393, 1.243347, 1.274048, 1.386108, 1.399902, 
    1.313782, 1.188141, 0.7401428, 0.5007629, 0.3675537, 0.2330933, 
    0.1566162, 0.08877563, 0.0736084, 0.1006775, 0.1239319, 0.137085, 
    0.1641541, 0.227417, 0.3023682, 0.3329163, 0.3284302, 0.329071, 0.32901, 
    0.3452148, 0.3479919, 0.3273926, 0.307251, 0.2817383, 0.2735596, 
    0.3437195, 0.4213257, 0.4539185, 0.4003296, 0.3487244, 0.3323975, 
    0.3479614, 0.3622742, 0.3453369, 0.3718262, 0.4780273, 1.392822, 
    1.606812, 1.287903, 1.232117, 1.10022, 1.05661, 1.085968, 1.094757, 
    1.10141, 1.153015, 1.245361, 1.365906, 1.436768, 1.388062, 1.38974, 
    1.380371, 1.322632, 1.212738,
  1.058777, 1.147949, 1.258881, 1.423798, 1.560455, 1.610382, 1.602325, 
    1.602478, 1.592865, 1.549133, 1.528168, 1.526489, 1.483948, 1.470673, 
    1.521271, 1.47464, 1.340057, 1.147339, 0.8456421, 0.5639038, 0.3579712, 
    0.2712402, 0.3670349, 0.4813538, 0.4744873, 0.394043, 0.2687378, 
    0.213562, 0.2177429, 0.2157898, 0.3106384, 0.2898254, 0.3479309, 
    1.388763, 1.343262, 1.340576, 1.017548, 0.6291199, 0.436615, 0.3467102, 
    0.145813, 0.1380615, 0.2461853, 0.2544556, 0.1382446, 0.04467773, 
    -0.1136475, -0.262146, -0.331665, -0.2941284, -0.1669006, -0.04064941, 
    -0.05804443, -0.1547852, -0.2175903, -0.1907959, 0.008026123, 0.2329102, 
    0.3744507, 0.5325012, 0.6930847, 0.8335571, 0.9251099, 0.9463196, 
    0.9223022, 0.9298401, 0.9423523, 0.9545288, 0.9503479, 0.9515381, 
    0.9940186, 1.026276, 1.068451, 1.092285, 1.118744, 1.073669, 0.9666748, 
    1.013458, 1.368103, 1.693298, 1.22171, 0.6929321, 0.412384, 0.4035339, 
    0.5451965, 0.6412354, 0.6361694, 0.6804199, 0.7162476, 0.775116, 
    0.7978821, 0.8144836, 0.8716431, 0.9302368, 0.9710693, 1.017426,
  1.165527, 1.172119, 1.149567, 1.116302, 1.11673, 1.138824, 1.232056, 
    1.363281, 1.446228, 1.492645, 1.530151, 1.627106, 1.718475, 1.674957, 
    1.56546, 1.485107, 1.460266, 1.429565, 1.32959, 1.169128, 1.051544, 
    0.9526978, 0.8823242, 0.867157, 0.8883362, 0.8286133, 0.670929, 
    0.5388184, 0.4943542, 0.5076599, 0.4735413, 0.4489441, 0.4671021, 
    0.5312805, 0.651001, 0.8057556, 0.9630737, 0.8654175, 0.7555237, 
    0.7130432, 0.6942444, 0.6918945, 0.7268677, 0.7459717, 0.679718, 
    0.469635, 0.08004761, -0.2209473, -0.3483887, -0.4688416, -0.5793457, 
    -0.6149597, -0.6022644, -0.6141663, -0.4963989, -0.242981, 0.06872559, 
    0.2938538, 0.4216614, 0.6226196, 0.8890991, 1.096497, 1.221649, 1.328918, 
    1.424255, 1.491058, 1.543182, 1.561798, 1.563873, 1.630157, 1.772247, 
    1.902252, 1.92804, 1.931, 1.914886, 1.842987, 1.726196, 1.622101, 
    1.539032, 1.457825, 1.394958, 1.243713, 0.9247131, 0.8189087, 0.9397278, 
    1.079803, 1.207489, 1.284576, 1.24942, 1.19458, 1.159576, 1.15976, 
    1.188995, 1.199768, 1.162323, 1.151459,
  1.24234, 1.183807, 1.156281, 1.096832, 1.038452, 1.004181, 1.045135, 
    1.111572, 1.144501, 1.148346, 1.198029, 1.32489, 1.432709, 1.509796, 
    1.518585, 1.497681, 1.501343, 1.523285, 1.460175, 1.32309, 1.219482, 
    1.068329, 0.9560242, 0.9293213, 0.9987183, 1.039093, 0.9914551, 
    0.9546509, 0.9418335, 0.8848572, 0.753418, 0.5855713, 0.4995117, 
    0.4732666, 0.4298401, 0.4301147, 0.5766602, 0.8433228, 1.023773, 
    1.084076, 1.055634, 1.123779, 1.259918, 1.225281, 1.118988, 1.055481, 
    0.8377991, 0.4025574, -0.08520508, -0.4661255, -0.6682434, -0.6954041, 
    -0.5701599, -0.4899597, -0.4472351, -0.2721252, 0.003692627, 0.1653137, 
    0.1523743, 0.367157, 0.8235779, 1.120148, 1.278564, 1.462402, 1.677124, 
    1.808899, 1.87796, 1.927185, 1.943665, 1.980957, 2.029449, 2.03772, 
    2.011444, 1.971588, 1.893799, 1.723846, 1.40921, 1.278168, 1.352051, 
    1.486694, 1.588074, 1.623413, 1.403534, 1.03421, 0.7997131, 0.8534241, 
    1.028473, 1.158173, 1.20993, 1.251587, 1.363647, 1.400116, 1.387421, 
    1.375671, 1.347443, 1.312744,
  1.378021, 1.45578, 1.576324, 1.662415, 1.689819, 1.708405, 1.734406, 
    1.730957, 1.738983, 1.764038, 1.726715, 1.732147, 1.728241, 1.770325, 
    1.893066, 1.97937, 2.111176, 2.24765, 2.17276, 1.739349, 1.440338, 
    1.304321, 1.138916, 1.055054, 1.141388, 1.295807, 1.368256, 1.390411, 
    1.383057, 1.370728, 1.328949, 1.195007, 1.062866, 0.9378967, 0.8462524, 
    0.8572083, 1.020813, 1.249329, 1.389862, 1.385315, 1.384552, 1.477295, 
    1.542053, 1.419464, 1.315826, 1.374664, 1.361633, 1.04953, 0.555542, 
    0.2490234, 0.1841736, 0.218689, 0.2655029, 0.2757874, 0.2723389, 
    0.328125, 0.444397, 0.5187683, 0.5533447, 0.7034912, 0.9830017, 1.174011, 
    1.28418, 1.445923, 1.630554, 1.65686, 1.644318, 1.733063, 1.788086, 
    1.777985, 1.781433, 1.794861, 1.789001, 1.72168, 1.550842, 1.21582, 
    1.131714, 1.304291, 1.439148, 1.446411, 1.462646, 1.414215, 1.306488, 
    1.023743, 0.967804, 1.20752, 1.53598, 1.715027, 1.671906, 1.610962, 
    1.621002, 1.613464, 1.572693, 1.533569, 1.484863, 1.412842,
  1.773529, 1.922821, 2.130493, 2.314301, 2.394684, 2.415588, 2.437134, 
    2.46109, 2.469238, 2.519897, 2.620758, 2.621979, 2.595154, 2.61676, 
    2.624725, 2.619904, 2.726746, 2.888763, 2.891357, 2.637421, 2.42099, 
    2.324188, 2.100739, 1.826111, 1.747711, 1.852539, 1.980377, 1.987305, 
    1.905548, 1.822876, 1.775696, 1.698181, 1.522003, 1.318817, 1.204376, 
    1.202209, 1.299927, 1.398376, 1.477814, 1.568237, 1.682404, 1.780853, 
    1.775024, 1.705383, 1.685883, 1.736328, 1.679565, 1.428497, 1.094666, 
    0.9387207, 0.9632568, 1.042053, 1.041748, 0.9651794, 0.9379578, 
    0.9899597, 1.040436, 1.149658, 1.2276, 1.295563, 1.430511, 1.544067, 
    1.589325, 1.622803, 1.676605, 1.662384, 1.628662, 1.634491, 1.636414, 
    1.608673, 1.58078, 1.559326, 1.500122, 1.383667, 1.220703, 1.166931, 
    1.463013, 1.585541, 1.772034, 1.829041, 1.744659, 1.567505, 1.329498, 
    1.176331, 1.242554, 1.506073, 1.789551, 2.017731, 2.076202, 2.055176, 
    2.046326, 1.98877, 1.905518, 1.880554, 1.859924, 1.77536,
  1.956299, 2.095245, 2.265106, 2.381439, 2.444611, 2.548004, 2.773834, 
    2.964966, 2.99942, 3.072205, 3.242371, 3.348907, 3.366089, 3.301178, 
    3.116028, 2.951904, 2.920898, 2.959961, 2.939911, 2.953186, 3.069275, 
    3.055206, 2.806, 2.544861, 2.437958, 2.429749, 2.367889, 2.220123, 
    2.039978, 1.903778, 1.89389, 1.88678, 1.748169, 1.604736, 1.551575, 
    1.528534, 1.572357, 1.5625, 1.487488, 1.614655, 1.973114, 2.096344, 
    2.084564, 2.034393, 2.089722, 2.218353, 2.282745, 2.096405, 1.799133, 
    1.698059, 1.81366, 1.87149, 1.800537, 1.661011, 1.562164, 1.545624, 
    1.614899, 1.708069, 1.75592, 1.757996, 1.769196, 1.804504, 1.774536, 
    1.715088, 1.733978, 1.731812, 1.696564, 1.658264, 1.604797, 1.501129, 
    1.378326, 1.316589, 1.300079, 1.227753, 1.198059, 1.259369, 1.486206, 
    1.829498, 2.302612, 1.989563, 1.849152, 1.651672, 1.583649, 1.630676, 
    1.822571, 2.007019, 2.073975, 2.102539, 2.110352, 2.11261, 2.065643, 
    2.028137, 1.987091, 1.920258, 1.90274, 1.908264,
  2.068695, 2.165039, 2.352356, 2.487701, 2.650848, 3.045959, 3.522125, 
    3.817444, 4.014648, 4.244843, 4.459045, 4.371552, 3.976563, 3.611908, 
    3.297729, 3.099701, 2.971344, 2.8927, 2.901215, 2.947601, 2.87793, 
    2.651947, 2.382202, 2.211395, 2.150177, 2.169861, 2.157166, 2.078522, 
    2.039703, 2.033661, 2.064392, 2.073303, 1.991364, 1.894775, 1.875671, 
    1.890259, 1.908386, 1.752228, 1.691254, 2.109833, 2.621613, 2.622833, 
    2.539978, 2.506531, 2.523651, 2.667969, 3.330597, 2.742584, 2.617645, 
    2.542664, 2.641602, 2.554352, 2.345123, 2.133453, 1.986847, 1.957947, 
    1.96582, 1.935272, 1.921173, 1.893494, 1.83316, 1.788666, 1.787445, 
    1.811401, 1.817169, 1.766083, 1.662506, 1.573181, 1.514191, 1.5112, 
    1.482819, 1.451019, 1.491791, 1.45697, 1.410278, 1.405396, 1.555145, 
    2.367554, 3.409119, 2.272217, 1.97168, 1.821106, 2.025909, 2.315216, 
    2.449768, 2.459045, 2.370514, 2.206055, 2.142853, 2.13678, 2.084503, 
    2.053711, 2.015167, 1.967377, 1.980804, 2.028381,
  1.989899, 2.077576, 2.217926, 2.396301, 2.692657, 3.113464, 3.447388, 
    4.065552, 4.344269, 4.026947, 3.568115, 3.184113, 2.80658, 2.51297, 
    2.36145, 2.362091, 2.323517, 2.230927, 2.156982, 2.033661, 1.900726, 
    1.841797, 1.826233, 1.845703, 1.80835, 1.835663, 1.924408, 1.931763, 
    2.035034, 2.182343, 2.2659, 2.227264, 2.128265, 2.013092, 2.025909, 
    2.006897, 1.942322, 1.996552, 2.401428, 4.380859, 3.165436, 3.053925, 
    3.156128, 3.095642, 2.943146, 2.931702, 3.062836, 3.651489, 2.852875, 
    2.596924, 2.466034, 2.381042, 2.290161, 2.218353, 2.129944, 2.06958, 
    2.000244, 1.943939, 1.936218, 1.904572, 1.880035, 1.879425, 1.846954, 
    1.856445, 1.874817, 1.865173, 1.881042, 1.852783, 1.761597, 1.761658, 
    1.7211, 1.650513, 1.661987, 1.583344, 1.5047, 1.407684, 1.424652, 
    2.83963, 4.432617, 3.41864, 1.925262, 1.965576, 2.352203, 2.636719, 
    2.635742, 2.497589, 2.406311, 2.338806, 2.290863, 2.201569, 2.117523, 
    2.092896, 2.040771, 1.975067, 1.929962, 1.935852,
  1.913147, 1.900513, 1.977142, 2.149933, 2.380219, 2.567383, 2.849884, 
    3.126251, 3.069855, 2.730591, 2.122131, 1.96817, 1.915894, 1.958588, 
    1.919403, 1.875061, 1.785736, 1.671295, 1.598816, 1.530853, 1.551178, 
    1.599091, 1.557495, 1.626648, 1.631165, 1.753052, 1.934937, 2.020508, 
    2.236511, 2.368347, 2.178436, 2.190094, 2.045074, 1.871552, 1.898041, 
    1.920258, 2.033203, 3.354187, 4.455292, 5.429993, 4.406158, 3.103058, 
    3.578461, 3.392761, 3.109955, 3.072144, 2.8638, 2.632813, 2.302917, 
    2.005249, 1.937317, 1.904938, 1.913422, 1.904816, 1.897644, 1.912628, 
    1.897675, 1.928955, 1.960541, 1.959381, 1.999664, 2.055664, 2.086578, 
    2.069397, 2.069122, 2.022583, 1.945587, 1.868683, 1.798187, 1.716278, 
    1.648254, 1.633392, 1.56842, 1.392365, 1.30365, 1.180847, 1.181793, 
    3.013489, 4.018494, 2.347046, 1.554291, 2.272186, 2.296356, 2.543365, 
    2.509308, 2.330811, 2.254883, 2.255005, 2.246613, 2.088531, 1.97818, 
    1.972198, 1.892975, 1.884979, 1.875214, 1.883453,
  1.767517, 1.726685, 1.733337, 1.839661, 2.146423, 4.10614, 4.645569, 
    3.593292, 2.508545, 2.236786, 2.28833, 2.414642, 2.337769, 2.286072, 
    2.175964, 2.060822, 2.05899, 2.016479, 1.992188, 1.95697, 1.981049, 
    2.039734, 2.082275, 2.147583, 2.179108, 2.246399, 2.367462, 2.40332, 
    2.323822, 1.937805, 2.197449, 3.989044, 3.46225, 2.81778, 3.279358, 
    3.614838, 3.887543, 4.340179, 4.707367, 4.727844, 3.505676, 2.251953, 
    2.004883, 2.025848, 2.267883, 2.430847, 2.160492, 1.749023, 1.668213, 
    1.783997, 1.876312, 1.91452, 1.96875, 1.990631, 1.911987, 1.916595, 
    1.909363, 1.951782, 1.977173, 2.017059, 2.031464, 1.991791, 2.028015, 
    1.982361, 1.938202, 1.817627, 1.64505, 1.518372, 1.485352, 1.382141, 
    1.302673, 1.271301, 1.18222, 1.150513, 1.059784, 1.000305, 1.139252, 
    2.655884, 4.135468, 2.513, 2.368103, 3.011658, 2.826294, 2.479889, 
    2.351685, 2.300201, 2.365814, 2.243378, 2.240479, 2.188995, 2.124084, 
    2.01535, 1.878265, 1.865051, 1.837036, 1.807465,
  1.557434, 1.55423, 1.696014, 1.887299, 2.632629, 4.443146, 4.249268, 
    2.68573, 2.559113, 2.241455, 2.213135, 2.406464, 2.362671, 2.297791, 
    2.364136, 2.418365, 2.494659, 2.498901, 2.466217, 2.463531, 2.406311, 
    2.404144, 2.319061, 2.21817, 2.164398, 2.101166, 2.007629, 2.013214, 
    2.040253, 2.011536, 2.850861, 4.661316, 4.339203, 3.966858, 4.305328, 
    4.332275, 4.670959, 4.608917, 4.166473, 3.727448, 2.934296, 1.757904, 
    1.418945, 1.548004, 1.826813, 1.989777, 1.967438, 1.933899, 1.995941, 
    2.103333, 2.094635, 1.991333, 1.928101, 1.901611, 1.871735, 1.836334, 
    1.798828, 1.805786, 1.791473, 1.826385, 1.819397, 1.768555, 1.700958, 
    1.58432, 1.511536, 1.350189, 1.284515, 1.158722, 1.087738, 1.093597, 
    1.06485, 1.088287, 1.008545, 1.031128, 0.8671265, 1.104675, 1.585083, 
    2.843689, 5.076294, 3.246307, 2.640564, 3.09082, 3.076813, 3.135345, 
    2.446411, 2.34314, 2.422607, 2.342896, 2.246674, 2.118561, 2.051239, 
    1.957092, 1.887817, 1.843567, 1.701752, 1.644379,
  1.60379, 1.778595, 2.023376, 2.468536, 3.347321, 2.922424, 1.935364, 
    1.575562, 2.262482, 2.888855, 2.367645, 2.517517, 2.875275, 2.333344, 
    2.249359, 2.355652, 2.276001, 2.2276, 2.141876, 2.087952, 2.040161, 
    2.007294, 1.988556, 1.961975, 1.948303, 1.96167, 1.954437, 2.051453, 
    2.228912, 2.315826, 2.892273, 4.297546, 4.479279, 4.70163, 4.749023, 
    4.519653, 4.542969, 4.137177, 3.176544, 2.936768, 2.361969, 1.786407, 
    1.89447, 2.141602, 2.173035, 2.145752, 2.157166, 2.196869, 2.167725, 
    2.152618, 2.101776, 2.014771, 1.955933, 1.89975, 1.849213, 1.798309, 
    1.770111, 1.794739, 1.810883, 1.794556, 1.722534, 1.588623, 1.480072, 
    1.360565, 1.327942, 1.168365, 1.08783, 1.003784, 1.00769, 1.018097, 
    1.049957, 1.052277, 0.8720093, 0.9806824, 1.01828, 1.558899, 2.261658, 
    3.39035, 6.031891, 3.611145, 2.14798, 3.146027, 3.117828, 3.03833, 
    2.999023, 2.461517, 2.293427, 2.258026, 2.091217, 1.874939, 1.786835, 
    1.706268, 1.675323, 1.654297, 1.601959, 1.592834,
  1.955475, 2.161316, 2.340973, 2.541382, 2.39212, 1.80249, 1.481323, 
    2.082764, 2.582092, 2.904694, 2.431549, 2.381226, 2.490112, 2.670776, 
    2.215881, 2.180664, 2.080353, 2.067383, 2.081116, 2.031982, 2.046753, 
    2.00174, 2.03476, 2.041534, 2.045959, 2.087097, 2.226685, 2.35788, 
    2.492004, 2.501343, 2.502991, 2.808533, 4.053589, 4.482361, 4.61972, 
    4.279572, 3.988922, 3.353668, 2.786499, 2.9198, 2.012299, 2.038086, 
    2.21463, 2.238403, 2.233124, 2.226715, 2.248444, 2.254578, 2.197479, 
    2.181976, 2.148102, 2.107117, 2.042053, 2.063995, 2.041473, 2.019989, 
    1.989258, 1.954926, 1.979248, 1.927399, 1.864441, 1.777679, 1.734253, 
    1.552155, 1.427521, 1.346527, 1.278198, 1.248901, 1.264984, 1.301758, 
    1.266022, 1.303009, 1.275848, 1.505707, 1.500244, 1.774994, 2.429169, 
    3.81958, 5.539978, 3.504364, 2.120331, 3.102783, 2.936188, 2.985016, 
    3.606964, 4.048737, 2.17865, 2.033875, 1.880798, 1.724731, 1.686707, 
    1.654938, 1.714996, 1.728699, 1.796021, 1.877533,
  2.362061, 2.548126, 2.725586, 2.689575, 2.402008, 2.103516, 2.189209, 
    2.785858, 3.072571, 3.167816, 3.383209, 2.422058, 2.45578, 2.957428, 
    2.307281, 2.249023, 2.18869, 2.188477, 2.22168, 2.203705, 2.21701, 
    2.209717, 2.236786, 2.223511, 2.281982, 2.384918, 2.502228, 2.585236, 
    2.579102, 2.532227, 2.370697, 2.350891, 2.491089, 3.247223, 3.609253, 
    3.730988, 3.428558, 2.449097, 3.091736, 1.990753, 1.983673, 2.229675, 
    2.307007, 2.274658, 2.31012, 2.343292, 2.300446, 2.27597, 2.228363, 
    2.184113, 2.161591, 2.175049, 2.201874, 2.249481, 2.235413, 2.203125, 
    2.146149, 2.1763, 2.218811, 2.199005, 2.146362, 2.055725, 1.974426, 
    1.886536, 1.812561, 1.777283, 1.730927, 1.77478, 1.774078, 1.812042, 
    1.789246, 1.795654, 1.794586, 1.843018, 1.811615, 2.32019, 4.172394, 
    5.762238, 4.214844, 3.109436, 2.795044, 2.949341, 2.805725, 3.013611, 
    4.030853, 4.134003, 2.125214, 2.063599, 1.942322, 1.912567, 1.931854, 
    1.958984, 2.107941, 2.168549, 2.260864, 2.321167,
  2.626526, 2.714264, 2.730988, 2.520172, 2.603302, 2.636871, 2.619263, 
    2.819458, 2.758057, 2.940613, 3.398499, 2.470581, 2.361145, 2.450928, 
    2.40683, 2.344818, 2.282013, 2.335144, 2.359772, 2.360596, 2.359894, 
    2.397461, 2.389709, 2.369995, 2.366211, 2.405151, 2.471497, 2.585602, 
    2.566925, 2.506592, 2.473267, 2.436737, 2.411591, 2.365753, 2.329926, 
    2.901154, 2.917755, 2.43634, 2.510101, 2.081238, 2.12851, 2.314636, 
    2.267822, 2.205475, 2.212433, 2.240875, 2.235474, 2.19342, 2.129242, 
    2.022247, 2.04422, 2.104614, 2.231781, 2.306183, 2.33548, 2.301239, 
    2.319611, 2.370758, 2.393616, 2.344452, 2.312134, 2.28598, 2.241821, 
    2.231049, 2.159973, 2.143616, 2.121948, 2.177521, 2.162415, 2.201813, 
    2.202911, 2.256165, 2.411072, 2.3703, 2.431122, 3.285278, 3.143372, 
    3.421234, 3.261017, 2.812195, 3.012573, 3.003235, 3.01062, 3.083618, 
    3.344208, 3.474609, 2.134644, 2.229492, 2.218872, 2.202515, 2.249481, 
    2.315125, 2.359039, 2.455658, 2.537506, 2.595245,
  2.742126, 2.744476, 2.621338, 2.406891, 2.697021, 2.725952, 2.658508, 
    2.54303, 2.631378, 2.895111, 2.954285, 2.448822, 2.499207, 2.505249, 
    2.472534, 2.437561, 2.372345, 2.420074, 2.421234, 2.458069, 2.467316, 
    2.478394, 2.475128, 2.478424, 2.456177, 2.429016, 2.394531, 2.414063, 
    2.45462, 2.42395, 2.318726, 2.362762, 2.494141, 2.473297, 2.454041, 
    2.376282, 2.294708, 2.349731, 2.727081, 2.12265, 2.12558, 2.242371, 
    2.157013, 2.084198, 2.020844, 2.02356, 2.068024, 2.099213, 2.135742, 
    2.071808, 2.137482, 2.189667, 2.271667, 2.369659, 2.412964, 2.406036, 
    2.420258, 2.463562, 2.465698, 2.480286, 2.44693, 2.492249, 2.485657, 
    2.471313, 2.429108, 2.424225, 2.445374, 2.462128, 2.499542, 2.54071, 
    2.645264, 2.679108, 2.73761, 2.639984, 2.584961, 2.700012, 2.897064, 
    3.289978, 3.279358, 3.083008, 3.138275, 3.252594, 3.273376, 3.287262, 
    3.017365, 2.679901, 2.668152, 2.372375, 2.400177, 2.396088, 2.418152, 
    2.505219, 2.545837, 2.63559, 2.677887, 2.700134,
  2.649353, 2.646027, 2.519012, 2.46225, 3.085663, 2.99826, 2.942322, 
    2.645203, 2.393372, 2.461731, 2.257965, 2.492889, 2.526764, 2.606567, 
    2.517334, 2.47168, 2.47287, 2.470184, 2.506836, 2.509003, 2.487701, 
    2.521576, 2.504547, 2.518799, 2.510895, 2.462372, 2.452728, 2.422791, 
    2.464203, 2.497375, 2.407013, 2.323242, 2.392822, 2.40213, 2.441864, 
    2.437103, 2.328583, 2.879944, 2.837036, 2.672913, 2.080078, 2.235687, 
    2.244141, 2.186523, 2.12558, 2.177948, 2.28067, 2.347137, 2.479034, 
    2.534454, 2.546936, 2.565033, 2.606232, 2.618347, 2.68573, 2.704437, 
    2.694153, 2.705383, 2.701965, 2.699219, 2.701691, 2.689819, 2.705719, 
    2.705719, 2.6987, 2.640961, 2.648163, 2.658264, 2.714233, 2.705658, 
    2.746246, 2.750519, 2.660614, 2.650848, 2.592773, 2.74173, 3.233582, 
    3.396667, 3.1409, 2.916809, 3.319061, 3.42395, 3.417816, 4.092834, 
    3.477478, 2.720398, 2.830292, 2.411713, 2.478241, 2.479736, 2.525665, 
    2.61499, 2.658752, 2.694855, 2.702606, 2.685486,
  2.474548, 2.494202, 2.461975, 2.79895, 3.086639, 3.0401, 2.879059, 
    2.521606, 2.467194, 2.318024, 2.036255, 3.32605, 2.59726, 2.641815, 
    2.602875, 2.511993, 2.514893, 2.428131, 2.436462, 2.485168, 2.508331, 
    2.560089, 2.571686, 2.552979, 2.574615, 2.516998, 2.52121, 2.946472, 
    2.668304, 2.449738, 2.723694, 2.508331, 2.493683, 2.179108, 2.247009, 
    2.943298, 2.751282, 2.522919, 2.44754, 2.06842, 2.171295, 2.235687, 
    2.267517, 2.285339, 2.377991, 2.497223, 2.583984, 2.642975, 2.665558, 
    2.727875, 2.762787, 2.744843, 2.742493, 2.780396, 2.847382, 2.919525, 
    2.944397, 2.95517, 2.983215, 2.996613, 2.993469, 2.962646, 2.96405, 
    2.925385, 2.971863, 2.992004, 3.049866, 3.068176, 3.023285, 3.025726, 
    2.971161, 2.827393, 2.64389, 2.46524, 2.54364, 2.679108, 2.596497, 
    2.969208, 2.933868, 3.44577, 3.526428, 4.553314, 4.598511, 4.446167, 
    3.493225, 2.436707, 2.425018, 2.457275, 2.500458, 2.523895, 2.57254, 
    2.540436, 2.593872, 2.617523, 2.591858, 2.504364,
  2.436127, 2.649597, 2.624786, 3.113556, 3.23938, 3.058197, 2.875183, 
    2.657166, 2.565247, 2.705658, 2.168945, 3.223877, 2.765961, 2.533325, 
    2.574677, 2.590363, 2.526184, 2.469727, 2.448151, 2.445984, 2.439056, 
    2.42923, 2.468048, 2.47641, 2.516846, 2.43457, 2.379547, 2.853119, 
    2.316803, 2.424927, 2.563477, 2.368622, 2.434631, 2.213745, 2.105988, 
    2.122406, 2.017578, 2.050507, 2.12558, 2.181, 2.183258, 2.214142, 
    2.230072, 2.228729, 2.323761, 2.407806, 2.516418, 2.585632, 2.57962, 
    2.608856, 2.632629, 2.613098, 2.608521, 2.622528, 2.648712, 2.657837, 
    2.71405, 2.726288, 2.751587, 2.7341, 2.751556, 2.722595, 2.757965, 
    2.79068, 2.847015, 2.893036, 2.928467, 3.017914, 3.078766, 3.059509, 
    2.942047, 2.742126, 2.600189, 2.362305, 2.225372, 2.635284, 3.153534, 
    3.522919, 3.049347, 3.656647, 4.175018, 4.448364, 3.867462, 2.362, 
    2.223389, 2.24649, 2.284943, 2.353302, 2.383209, 2.444916, 2.498199, 
    2.544708, 2.596893, 2.50885, 2.501282, 2.395905,
  3.527344, 2.870453, 3.573761, 3.832764, 3.258179, 3.098053, 3.199677, 
    2.979309, 3.125641, 3.616364, 3.252533, 2.213867, 2.848969, 2.552673, 
    2.544342, 2.575989, 2.566345, 2.520721, 2.469147, 2.481049, 2.495941, 
    2.487732, 2.390747, 2.367188, 2.471527, 2.511993, 2.912445, 2.936462, 
    2.370453, 2.304626, 2.271759, 2.585266, 2.369415, 2.406128, 2.151245, 
    2.024323, 2.054626, 2.108856, 2.109894, 2.138672, 2.167053, 2.219086, 
    2.240387, 2.253723, 2.311523, 2.396423, 2.474274, 2.555847, 2.592438, 
    2.613953, 2.653961, 2.680481, 2.682373, 2.664581, 2.682922, 2.635284, 
    2.640045, 2.596619, 2.543793, 2.494812, 2.450012, 2.415375, 2.416779, 
    2.44812, 2.458069, 2.506836, 2.59845, 2.687775, 2.83905, 2.938354, 
    2.961243, 2.690887, 2.396637, 2.309906, 2.443176, 2.848511, 3.923187, 
    5.054993, 4.221344, 5.048248, 4.25, 4.057281, 2.514526, 2.319458, 
    2.311432, 2.286469, 2.326813, 2.353577, 2.375641, 2.38678, 2.451477, 
    2.489075, 2.510223, 2.566345, 3.576965, 3.563599,
  3.199738, 3.176361, 3.363678, 3.515869, 3.476837, 3.492706, 3.151581, 
    3.176361, 3.368866, 3.587646, 3.476166, 3.538483, 3.748932, 3.099365, 
    2.625519, 2.627197, 2.727936, 2.678864, 2.69162, 2.684052, 2.755798, 
    3.045197, 2.535278, 2.411316, 2.410614, 2.380005, 2.472534, 3.226166, 
    2.425537, 2.295502, 2.3013, 2.23465, 2.28775, 2.624298, 2.311279, 
    2.209229, 2.246155, 2.272125, 2.26535, 2.256439, 2.273193, 2.296021, 
    2.28418, 2.29422, 2.288605, 2.324554, 2.360046, 2.37674, 2.432617, 
    2.45813, 2.523132, 2.575256, 2.624786, 2.677795, 2.72995, 2.729614, 
    2.730286, 2.712646, 2.6474, 2.62323, 2.579224, 2.542267, 2.542145, 
    2.556763, 2.55896, 2.581238, 2.609558, 2.646545, 2.782806, 2.855682, 
    2.840485, 2.75351, 2.79837, 2.74649, 3.377747, 3.586975, 4.096954, 
    5.106293, 4.206329, 3.786865, 2.3237, 2.270325, 2.362122, 2.419342, 
    2.330475, 2.318115, 2.324097, 2.361328, 2.405212, 2.397339, 2.432312, 
    2.428589, 2.698761, 3.336243, 3.517456, 3.324097,
  4.169006, 3.552643, 3.080536, 3.106232, 3.079163, 3.040894, 3.000305, 
    3.021545, 3.244781, 3.639252, 4.016449, 4.566528, 4.313141, 3.755676, 
    2.708405, 2.674622, 2.753754, 2.72583, 2.742432, 2.772644, 3.844086, 
    3.699677, 2.652405, 2.524567, 2.383545, 2.249939, 2.21402, 3.085083, 
    3.097992, 2.622589, 2.298187, 2.278564, 2.308594, 2.632019, 2.258209, 
    2.267975, 2.288147, 2.287354, 2.312775, 2.295105, 2.305389, 2.302094, 
    2.324585, 2.33725, 2.361969, 2.370758, 2.393951, 2.395721, 2.463074, 
    2.476501, 2.539246, 2.577789, 2.631317, 2.696289, 2.740631, 2.791016, 
    2.76413, 2.774628, 2.727722, 2.682739, 2.649078, 2.62265, 2.583527, 
    2.563568, 2.555908, 2.531769, 2.515839, 2.594086, 2.633087, 2.689819, 
    2.772766, 2.876282, 4.157043, 3.926361, 2.605804, 2.724487, 2.664063, 
    2.562836, 2.454498, 2.466522, 2.417236, 2.439331, 2.351624, 2.314667, 
    2.29068, 2.326111, 2.34259, 2.415222, 2.411072, 2.449402, 2.501892, 
    2.777069, 3.913269, 4.299042, 4.209442, 3.94696,
  4.073975, 3.864014, 3.6091, 3.334381, 3.063232, 2.892578, 2.822662, 
    2.73645, 2.8591, 3.149811, 4.201019, 4.677673, 4.077271, 3.905396, 
    3.708801, 2.736511, 2.734375, 2.714264, 2.721069, 2.751953, 4.414368, 
    4.507111, 2.7901, 2.672699, 2.50351, 2.299347, 3.066864, 2.622253, 
    2.096344, 1.928436, 2.184509, 2.206238, 2.094604, 2.09726, 2.129822, 
    2.165619, 2.234283, 2.297791, 2.323425, 2.318726, 2.357086, 2.346008, 
    2.357147, 2.332153, 2.307281, 2.294067, 2.311737, 2.306, 2.355988, 
    2.406311, 2.443817, 2.489044, 2.550934, 2.62619, 2.630157, 2.643494, 
    2.602356, 2.565765, 2.497833, 2.412201, 2.328583, 2.281311, 2.302734, 
    2.319641, 2.317627, 2.303009, 2.22879, 2.160889, 2.234497, 3.632629, 
    4.021423, 3.6138, 2.695831, 2.246735, 2.419464, 2.477722, 2.495239, 
    2.515961, 2.47876, 2.424866, 2.349487, 2.309174, 2.204865, 2.13913, 
    2.113922, 2.072571, 2.142303, 2.227661, 2.275146, 2.375977, 2.406708, 
    2.849213, 4.525146, 4.503693, 4.413147, 4.179688,
  4.009583, 3.794067, 3.785614, 3.678558, 3.419861, 3.25769, 3.198975, 
    3.088806, 3.039124, 2.853394, 2.508667, 4.164642, 4.026825, 4.079712, 
    4.387299, 3.889252, 2.709686, 2.739441, 2.813141, 2.633789, 4.121735, 
    4.322784, 3.773376, 3.735687, 2.601685, 3.281952, 3.263031, 2.642517, 
    1.609253, 1.391968, 2.007568, 2.129364, 2.000214, 2.055817, 2.026001, 
    1.999146, 2.009308, 2.055664, 2.1026, 2.107208, 2.149078, 2.170746, 
    2.204041, 2.201965, 2.185608, 2.173767, 2.164581, 2.136108, 2.167694, 
    2.249146, 2.317749, 2.367188, 2.429932, 2.513855, 2.542145, 2.563751, 
    2.572174, 2.522339, 2.422607, 2.29657, 2.134216, 1.950592, 1.861847, 
    1.92804, 2.023834, 2.106201, 2.094208, 2.107086, 2.569, 2.937683, 
    2.691345, 2.144867, 1.77298, 1.974091, 2.258423, 2.362244, 2.467224, 
    2.575653, 2.596497, 2.506104, 2.424286, 2.33847, 2.195374, 2.016541, 
    1.923645, 1.865631, 1.843231, 1.897247, 1.97467, 2.067444, 2.141846, 
    2.644989, 4.216614, 4.178528, 4.160431, 4.277222,
  4.217712, 4.118683, 3.780457, 3.807739, 3.775024, 3.534851, 3.294525, 
    3.324921, 3.444733, 3.306335, 2.446991, 4.086304, 3.791779, 3.616516, 
    4.013672, 4.049286, 2.800323, 3.011719, 4.416016, 4.072205, 3.911682, 
    3.196686, 2.963806, 3.065094, 3.088257, 3.112823, 3.177917, 2.481903, 
    2.073608, 2.122681, 2.245148, 2.383026, 2.083984, 1.992645, 1.944855, 
    1.981903, 2.050476, 2.045563, 2.069122, 2.026276, 2.043427, 2.048828, 
    2.017853, 2.022522, 1.974609, 1.910858, 1.830078, 1.774048, 1.784882, 
    1.831238, 1.923706, 2.034363, 2.118561, 2.200958, 2.273651, 2.345825, 
    2.367462, 2.387329, 2.402985, 2.332306, 2.225464, 2.092773, 1.927795, 
    1.884888, 1.877655, 1.93692, 2.191986, 2.506927, 2.604553, 2.82077, 
    2.609589, 2.092194, 1.782227, 1.921021, 2.027802, 2.129425, 2.267761, 
    2.388672, 2.585602, 2.579559, 2.584717, 2.540619, 2.491974, 2.406189, 
    2.280029, 2.151367, 2.06427, 2.077484, 2.024292, 1.970123, 2.016144, 
    2.266907, 3.630676, 3.979248, 3.862762, 4.056244,
  3.782166, 4.015442, 3.928375, 3.795502, 3.717926, 3.398285, 3.425659, 
    3.352478, 3.304871, 3.674164, 3.79187, 3.708435, 3.827881, 3.584595, 
    3.64267, 3.750488, 3.383301, 3.734009, 4.228027, 4.055817, 4.228333, 
    4.036438, 3.797974, 4.351715, 2.633881, 3.634033, 2.901062, 2.564453, 
    2.784882, 3.387085, 2.915497, 2.829529, 2.842041, 2.131775, 1.984833, 
    1.981903, 2.042786, 2.098236, 2.142365, 2.066681, 2.018433, 2.007874, 
    1.980316, 1.962036, 1.881897, 1.833923, 1.769135, 1.67749, 1.613159, 
    1.561066, 1.604401, 1.699219, 1.819641, 1.949341, 2.06427, 2.16452, 
    2.213867, 2.221436, 2.207275, 2.221436, 2.195465, 2.121002, 2.016754, 
    1.879547, 1.846344, 2.025391, 2.795959, 2.931335, 2.876709, 3.015533, 
    2.502533, 2.342255, 2.101807, 2.241608, 1.934479, 1.967224, 2.1008, 
    2.175201, 2.332428, 2.417847, 2.493164, 2.510345, 2.474823, 2.430511, 
    2.367584, 2.346069, 2.338074, 2.297546, 2.196381, 2.076508, 1.967529, 
    1.951111, 2.420105, 3.607239, 3.784698, 3.564789,
  3.428223, 3.353485, 3.11676, 3.329742, 3.419861, 2.630585, 2.985046, 
    3.06485, 2.596863, 3.153992, 3.143585, 3.220306, 3.443054, 3.013245, 
    2.228333, 2.456482, 2.640442, 3.218292, 4.411865, 4.088837, 4.273895, 
    8.061707, 5.909653, 4.772827, 4.373322, 5.028015, 4.138824, 2.85376, 
    3.213715, 4.224182, 3.737732, 3.813171, 3.549011, 1.619324, 1.514709, 
    2.090881, 2.197418, 2.233734, 2.236481, 2.251617, 2.228241, 2.168427, 
    2.117554, 2.056519, 1.952759, 1.866333, 1.796204, 1.762238, 1.710419, 
    1.632416, 1.597565, 1.564514, 1.619995, 1.771027, 1.891724, 1.989105, 
    2.060547, 2.050385, 2.035614, 2.080017, 2.087158, 2.030792, 1.960724, 
    1.858002, 1.957092, 2.717194, 2.546112, 2.196655, 2.105743, 2.236816, 
    2.103943, 1.971008, 1.706818, 1.766357, 2.026093, 1.911316, 2.003052, 
    2.044342, 2.069458, 2.020447, 2.047211, 2.142639, 2.201691, 2.172638, 
    2.12323, 2.105804, 2.105286, 2.198242, 2.325195, 2.248566, 2.0625, 
    1.966064, 1.943512, 2.273041, 3.335175, 3.479767,
  3.07373, 2.655304, 2.72406, 2.794342, 2.70636, 2.501099, 2.234131, 
    2.248566, 2.565125, 2.688202, 2.627167, 2.756622, 3.003204, 2.885773, 
    2.176544, 2.196075, 1.963867, 2.453369, 5.517792, 5.250488, 5.501984, 
    5.482315, 5.280701, 4.460114, 4.268768, 3.848969, 3.423004, 2.683197, 
    4.771057, 4.426666, 3.2547, 3.809418, 3.380157, 2.352234, 2.420685, 
    2.219269, 2.75589, 2.81485, 2.31015, 2.265442, 2.246887, 2.214203, 
    2.195892, 2.164063, 2.117371, 2.037109, 1.938721, 1.917969, 1.914673, 
    1.864594, 1.809692, 1.752869, 1.728882, 1.761597, 1.848755, 1.971283, 
    2.045227, 2.067383, 2.087616, 2.046356, 2.001831, 2.016876, 2.016144, 
    1.929932, 2.143829, 2.016998, 1.584045, 1.498657, 1.61145, 2.030823, 
    2.007721, 2.26123, 2.277954, 2.156677, 2.323395, 2.462402, 2.252533, 
    2.164124, 2.15506, 2.186646, 2.14035, 1.898163, 1.733215, 1.804626, 
    1.81192, 1.727875, 1.626251, 1.659698, 1.973175, 2.27948, 2.28894, 
    2.131317, 1.964996, 2.08847, 2.423767, 3.219055,
  2.719238, 2.52832, 2.604553, 2.63208, 2.667511, 2.461548, 2.720459, 
    2.163879, 2.287811, 2.403076, 3.274078, 4.676453, 3.957672, 2.427917, 
    2.195435, 2.669861, 1.905823, 1.7789, 2.937927, 4.885178, 4.430038, 
    4.247559, 4.898987, 3.454269, 3.878479, 3.670776, 4.207275, 4.726471, 
    5.997742, 5.791382, 4.733185, 4.383362, 4.820984, 5.114349, 4.967651, 
    2.654053, 2.446045, 3.023163, 2.466125, 2.465363, 2.472931, 2.486053, 
    2.493561, 2.409821, 2.322784, 2.283569, 2.202606, 2.116608, 2.047394, 
    2.036194, 2.036896, 1.958771, 1.913452, 1.956329, 1.965118, 1.95163, 
    1.963806, 1.979187, 2.022064, 2.04895, 2.051697, 1.9823, 1.936005, 
    2.117218, 2.927155, 3.889099, 4.276276, 4.064148, 3.033112, 1.180054, 
    1.206848, 2.132294, 2.875641, 2.685364, 2.402649, 2.767151, 3.169128, 
    3.094299, 2.896149, 2.759766, 2.552917, 2.194092, 1.681335, 1.388123, 
    1.522186, 1.454681, 1.181824, 0.8501282, 0.9023438, 1.522736, 2.006653, 
    2.05957, 1.973877, 2.170959, 2.889832, 3.024445,
  2.686615, 2.440826, 2.598175, 3.417664, 2.741486, 3.371918, 3.598236, 
    2.719696, 2.036224, 2.198792, 2.947876, 3.877258, 3.871979, 2.298218, 
    2.538818, 3.324402, 3.674438, 2.613312, 2.908112, 4.815735, 4.337738, 
    3.972748, 3.86795, 4.10257, 4.153015, 3.961884, 3.654465, 3.37973, 
    3.936829, 3.953018, 3.602692, 3.794159, 3.665268, 3.431152, 3.663895, 
    3.60347, 2.745544, 2.485596, 3.137146, 3.344177, 3.658539, 3.041168, 
    2.585663, 2.310577, 2.159668, 2.113007, 2.119293, 2.106354, 2.018188, 
    1.946625, 1.985535, 2.032288, 2.074341, 2.138214, 2.19223, 2.183838, 
    2.145386, 2.094666, 2.062439, 2.034454, 2.022675, 1.974152, 2.008087, 
    2.30191, 3.625885, 3.737152, 2.992218, 2.473999, 2.538574, 2.465454, 
    2.92157, 3.731293, 4.273865, 3.687073, 3.280487, 4.455902, 4.813904, 
    4.586884, 4.038757, 3.691498, 2.967957, 2.290558, 2.301483, 1.993896, 
    1.734192, 1.435028, 0.8988953, 0.544281, 0.5380249, 0.9596252, 1.512512, 
    1.877808, 1.95932, 2.026886, 2.674377, 2.730072,
  2.700684, 2.909973, 4.592621, 4.766632, 3.839905, 4.088959, 4.382263, 
    3.052368, 2.284546, 2.025574, 2.094635, 2.414368, 2.623596, 2.333191, 
    2.28772, 3.980957, 4.754517, 4.804779, 4.787659, 5.166168, 5.235046, 
    4.856354, 3.672501, 3.287323, 3.895325, 3.634781, 3.390656, 3.457123, 
    3.538483, 2.915512, 2.593506, 3.183807, 3.108414, 3.000092, 3.450012, 
    3.475143, 2.814468, 2.538086, 3.129639, 2.874084, 2.666077, 2.405334, 
    2.325043, 2.145325, 2.022095, 1.957184, 1.920654, 1.993011, 2.020996, 
    1.977173, 2.052246, 2.199646, 2.285065, 2.310974, 2.378937, 2.45694, 
    2.393066, 2.275513, 2.23172, 2.193115, 2.211639, 2.150848, 2.117126, 
    2.511169, 3.824127, 3.21759, 2.771515, 2.905487, 3.648071, 4.586365, 
    4.969849, 4.494415, 5.049103, 4.841644, 5.639282, 5.926483, 5.862152, 
    5.930878, 6.273193, 6.013306, 3.544708, 2.824951, 2.290283, 1.87088, 
    1.69281, 1.604736, 1.078735, 0.3865356, 0.1334839, 0.453064, 0.8852844, 
    1.322662, 1.641693, 1.790619, 2.031097, 2.565186,
  1.996735, 2.360657, 3.585022, 3.963165, 3.782318, 4.006989, 4.077881, 
    3.457001, 3.18335, 3.169434, 3.079468, 2.912354, 2.962402, 2.970032, 
    3.008942, 3.235321, 3.659607, 3.502045, 3.044495, 3.284271, 4.206421, 
    4.623596, 3.798874, 3.165466, 3.251572, 2.953598, 3.045273, 2.990829, 
    2.987061, 2.977493, 3.301895, 3.301453, 2.872345, 2.991043, 3.4655, 
    3.04454, 2.723267, 4.159912, 8.413956, 4.793518, 2.872345, 2.572266, 
    2.53302, 2.290619, 2.205627, 2.196075, 2.155701, 2.095673, 2.114929, 
    2.164825, 2.234924, 2.395782, 2.597168, 2.736877, 2.809601, 2.861115, 
    2.840057, 2.670746, 2.51181, 2.449371, 2.446594, 2.416534, 2.989258, 
    3.479248, 3.691895, 3.802979, 4.294586, 5.551788, 6.663391, 6.813263, 
    6.079132, 6.31076, 6.655945, 6.893997, 7.441833, 8.106537, 8.188065, 
    7.372604, 6.822617, 6.518661, 4.194916, 5.879211, 3.111725, 2.358124, 
    1.873291, 1.464752, 0.7315369, -0.2174377, -0.7832336, -0.5765381, 
    0.1332703, 0.9026794, 1.396301, 1.53894, 1.642761, 1.721283,
  1.706146, 1.853027, 2.393738, 2.731659, 3.194183, 3.381104, 3.644501, 
    3.688141, 3.259796, 2.844086, 2.429138, 2.259857, 2.393768, 2.872803, 
    2.987793, 2.636993, 2.338348, 2.562408, 2.573059, 2.563583, 2.723724, 
    3.086487, 3.049652, 3.303604, 3.418121, 3.292725, 3.140305, 3.177048, 
    2.803925, 2.897079, 3.376068, 2.633743, 2.780548, 3.469604, 3.477097, 
    2.543121, 2.892273, 5.568893, 10.26085, 6.951538, 3.918671, 3.354126, 
    3.823395, 2.437897, 2.415558, 2.296875, 2.181946, 2.012115, 2.025696, 
    2.227509, 2.42514, 2.742523, 3.098236, 3.345612, 3.308777, 3.253235, 
    3.113312, 2.92807, 2.767029, 2.683044, 2.649445, 4.286652, 4.512726, 
    4.607605, 4.627777, 4.847015, 5.708893, 6.889877, 7.675095, 7.665253, 
    7.60556, 7.695328, 8.752121, 10.10895, 12.00916, 17.4639, 11.63095, 
    9.014938, 8.005371, 8.822113, 9.22496, 7.692108, 3.731506, 2.315613, 
    1.687195, 1.531738, 0.9805908, 0.05776978, -0.6775208, -0.7682495, 
    -0.1921387, 0.6628418, 1.233459, 1.382477, 1.380249, 1.601532,
  1.237671, 1.430359, 1.658173, 3.095673, 2.874512, 2.098022, 2.203766, 
    2.666321, 2.531006, 2.694946, 2.969391, 2.822021, 2.738953, 3.033966, 
    2.984802, 2.974548, 2.754639, 2.630692, 2.771057, 2.924637, 3.19696, 
    3.40686, 3.268692, 3.036087, 3.072021, 3.012115, 3.348068, 2.668961, 
    2.654572, 2.725464, 2.751251, 2.578079, 2.845917, 3.204758, 2.687515, 
    2.471558, 3.343567, 6.100418, 10.26089, 10.75653, 10.18097, 8.383148, 
    6.029831, 4.498779, 3.428375, 2.940643, 3.09201, 3.609253, 3.769012, 
    3.832611, 4.094421, 4.485931, 4.609619, 4.77832, 6.942871, 3.846497, 
    3.500946, 3.008484, 2.932983, 3.207458, 5.823029, 6.046844, 6.040787, 
    6.113434, 6.637466, 7.758896, 8.248535, 7.99025, 7.484589, 7.673981, 
    9.299301, 11.04709, 15.80458, 18.4277, 20.37163, 20.50381, 12.83519, 
    10.06551, 10.00398, 11.31625, 15.22769, 9.480957, 5.393921, 3.844116, 
    2.287323, 2.163483, 1.833405, 1.241699, 0.7218323, 0.5707397, 0.7484741, 
    1.039551, 1.25296, 1.348053, 1.345978, 1.484528,
  0.90802, 1.188904, 2.18634, 2.307587, 2.740723, 3.321777, 3.246307, 
    2.887207, 2.362854, 2.069305, 2.240936, 2.691315, 2.838638, 2.918335, 
    3.314087, 3.758804, 3.573517, 3.200348, 3.013947, 3.084, 3.254044, 
    3.94989, 4.056854, 4.147476, 3.991562, 3.227692, 3.616547, 3.65184, 
    3.513809, 3.371826, 2.99617, 2.73674, 2.909195, 3.256989, 3.758865, 
    4.060562, 4.210892, 4.352875, 5.109589, 5.223663, 5.586151, 5.044159, 
    5.261993, 5.778595, 6.13739, 7.022934, 8.80014, 13.34103, 12.59183, 
    12.63324, 13.69482, 14.71585, 11.76697, 10.62776, 9.63559, 8.885895, 
    8.518967, 7.658249, 7.363266, 7.244812, 7.205887, 7.350037, 7.606232, 
    7.843262, 7.860825, 8.591339, 8.77327, 8.668503, 8.537323, 8.966171, 
    10.62625, 13.18275, 14.94478, 16.68526, 17.07927, 15.88747, 11.9874, 
    11.00047, 12.34293, 14.32236, 16.26944, 13.68904, 9.401489, 6.543274, 
    5.855347, 2.678802, 1.944611, 1.658173, 1.454834, 1.488556, 1.403168, 
    1.089355, 0.5020447, 0.2110291, 0.6318054, 0.841095,
  0.5424805, 0.7898254, 0.6204224, 2.081421, 2.591766, 3.102722, 6.42334, 
    3.950012, 3.655884, 3.18927, 2.983795, 3.174957, 3.348923, 3.178467, 
    2.947678, 2.670715, 2.992142, 3.347549, 4.079575, 4.683151, 4.753983, 
    4.85907, 4.544083, 4.405609, 4.617203, 3.867401, 3.555359, 3.52951, 
    3.53302, 3.335312, 3.314011, 3.184647, 3.594803, 4.342072, 4.352036, 
    4.734848, 5.30809, 5.026047, 5.661285, 5.664337, 5.676315, 5.714478, 
    5.84761, 6.00444, 6.000092, 5.741165, 5.902023, 6.339859, 7.363754, 
    9.6633, 11.43999, 16.91866, 11.77267, 10.03712, 8.569489, 7.843399, 
    7.55217, 7.814209, 7.634781, 7.279587, 7.682953, 8.206924, 8.637848, 
    9.033493, 9.257385, 8.675018, 8.435043, 8.420731, 8.399612, 8.801254, 
    8.94838, 9.461609, 10.40152, 11.0941, 11.84, 11.49142, 10.60802, 
    10.06995, 9.84584, 10.17137, 10.86678, 10.97098, 8.462936, 7.03656, 
    5.911819, 5.440338, 4.62059, 1.64624, 1.894196, 2.531067, 3.328918, 
    5.470032, 2.543457, 1.265381, 0.4125366, 0.2746277,
  1.090454, 0.6763916, 0.463562, 0.2519836, -0.1156616, 2.210114, 2.726868, 
    3.07074, 3.549713, 3.967102, 4.833496, 6.897736, 8.59729, 9.33197, 
    5.549194, 4.692322, 3.922089, 3.884781, 4.373657, 4.907639, 5.235825, 
    5.411728, 5.312775, 5.06778, 4.925079, 4.840897, 4.516617, 4.151382, 
    3.792801, 3.929642, 4.337646, 4.638687, 4.87027, 4.806076, 5.310242, 
    5.245529, 5.074951, 5.426376, 5.681137, 6.120056, 6.363815, 6.284134, 
    6.185501, 6.328918, 6.637314, 6.337906, 6.437393, 6.576843, 7.219681, 
    8.204971, 9.84819, 11.03922, 11.3905, 9.711533, 9.046509, 9.002625, 
    9.020462, 9.310165, 8.623779, 9.491486, 10.08849, 9.425018, 9.554108, 
    9.164474, 8.782379, 8.116028, 7.965378, 8.345322, 8.980103, 9.008926, 
    9.070984, 8.824036, 9.139999, 9.440308, 9.864655, 10.15575, 10.39253, 
    10.27065, 10.21844, 10.04449, 9.853348, 8.094696, 8.158813, 7.473709, 
    6.529694, 6.010895, 5.576447, 5.730804, 6.883926, 8.627106, 12.71793, 
    13.59157, 13.3616, 7.987915, 3.569061, 2.067871,
  3.689789, 2.433777, 1.581757, 1.194305, 0.8101196, 1.067017, 1.880402, 
    3.018921, 4.32666, 5.702484, 7.218597, 9.440613, 11.7652, 12.30392, 
    10.09569, 8.451263, 7.291168, 7.058548, 6.844101, 6.050858, 5.864349, 
    5.818375, 5.877304, 5.700867, 5.503403, 5.27475, 5.256851, 5.070724, 
    5.084457, 5.569931, 5.435242, 5.702164, 5.707306, 5.738098, 5.699432, 
    5.26915, 5.855423, 5.976776, 6.248199, 6.348328, 6.077164, 6.319611, 
    6.324692, 6.324829, 6.50737, 6.713028, 6.827759, 6.889008, 6.902161, 
    7.133606, 7.442596, 7.820465, 8.156525, 8.385361, 8.729309, 8.847672, 
    8.968826, 9.161148, 9.215042, 9.258286, 9.106979, 8.939468, 8.70372, 
    8.66655, 8.262253, 7.954315, 7.874756, 8.052032, 8.263229, 8.514328, 
    8.557755, 8.573914, 8.138824, 8.766037, 9.216217, 9.401047, 9.706268, 
    9.13913, 9.352753, 9.630356, 8.637665, 8.523773, 8.155426, 7.033279, 
    6.273331, 5.559586, 4.410568, 4.12468, 4.947739, 6.450287, 8.483673, 
    10.3609, 11.25816, 11.53421, 11.53963, 8.033813,
  10.16762, 7.091919, 4.34964, 3.286407, 3.856934, 7.143402, 11.48877, 
    12.20152, 12.76137, 12.49443, 12.04086, 11.60056, 11.02991, 10.37495, 
    9.629761, 9.184128, 8.582047, 8.353729, 8.107758, 7.808014, 7.498199, 
    7.207504, 6.93335, 6.699692, 6.396835, 7.052353, 7.060501, 6.832901, 
    6.920792, 7.219345, 7.211792, 6.039017, 6.320404, 6.368835, 6.303543, 
    6.248718, 6.318497, 6.379318, 6.509186, 6.550659, 6.584641, 6.660889, 
    6.741028, 6.828018, 6.907959, 6.878265, 6.865067, 6.911209, 6.996826, 
    7.118896, 7.279114, 7.440964, 7.637589, 7.826904, 8.000153, 8.094482, 
    8.135956, 8.117401, 8.088623, 8.152359, 8.29039, 8.392334, 8.397018, 
    8.437775, 8.492401, 8.220917, 8.186996, 8.07547, 8.005539, 8.068176, 
    8.166885, 8.435562, 8.564209, 8.746765, 8.79155, 8.551254, 9.056061, 
    8.55484, 9.189529, 8.471695, 7.884201, 7.607834, 7.42807, 7.102097, 
    6.817001, 6.338684, 5.900604, 5.634003, 5.917526, 6.770584, 8.00679, 
    9.367081, 10.55263, 11.14331, 11.26221, 10.8031,
  10.20679, 9.760818, 9.268402, 8.77066, 9.577759, 9.734528, 9.965057, 
    10.25562, 10.43973, 10.3952, 10.23752, 9.93335, 9.577164, 9.214996, 
    8.842529, 8.613815, 8.441437, 8.329697, 8.227631, 8.142212, 7.969742, 
    7.791092, 7.524948, 7.238617, 6.991806, 7.212326, 7.181717, 6.286545, 
    6.70697, 6.81427, 6.913956, 7.015778, 7.106064, 7.035767, 6.982574, 
    6.820328, 6.649094, 6.529968, 6.476654, 6.439209, 6.451065, 6.494034, 
    6.602295, 6.756729, 6.868195, 6.97821, 7.042725, 7.117401, 7.220596, 
    7.313431, 7.396042, 7.495132, 7.617981, 7.684586, 7.649628, 7.620789, 
    7.62027, 7.613617, 7.650986, 7.737839, 7.905685, 8.070343, 8.284988, 
    8.48999, 8.696304, 8.839005, 8.963165, 8.955612, 8.970459, 8.931915, 
    9.113953, 8.293243, 8.364868, 8.512589, 8.396103, 8.224701, 8.05275, 
    7.915253, 7.68634, 7.41571, 7.197021, 6.936935, 6.723129, 6.631714, 
    6.541489, 6.520004, 6.445389, 6.579178, 7.077682, 7.836014, 8.753723, 
    9.563293, 10.76291, 10.64507, 10.72391, 10.49493,
  10.75575, 10.71219, 10.61017, 10.4875, 10.29689, 10.1424, 10.02039, 
    9.811279, 9.637314, 9.498398, 9.40654, 9.333023, 9.247147, 9.142075, 
    9.020264, 8.912064, 8.813171, 8.719482, 8.622925, 8.512115, 8.397476, 
    8.299957, 8.215652, 8.102356, 7.980484, 7.878464, 7.730881, 7.524689, 
    7.420654, 7.356003, 7.324554, 7.290894, 7.209061, 7.173584, 7.130478, 
    7.16864, 7.192535, 7.169403, 7.165573, 7.20842, 7.2491, 7.263947, 
    7.272552, 7.293243, 7.332825, 7.3685, 7.387192, 7.396881, 7.437714, 
    7.499817, 7.578201, 7.61116, 7.659134, 7.6633, 7.721237, 7.849625, 
    7.93895, 8.037842, 8.147614, 8.209717, 8.330215, 8.49617, 8.62175, 
    8.725998, 8.848907, 8.951309, 9.069931, 9.171692, 9.258224, 9.375854, 
    9.371368, 9.452225, 9.608154, 9.656723, 9.656799, 9.7034, 9.684387, 
    9.5168, 9.663696, 9.754837, 9.819733, 9.701462, 9.729309, 9.725723, 
    9.852951, 10.00159, 10.05412, 10.10809, 10.34039, 10.4648, 10.71629, 
    10.97339, 11.06264, 11.02332, 10.94891, 10.85822,
  10.30843, 10.30269, 10.19618, 10.13979, 10.08673, 10.05074, 9.972672, 
    9.893631, 9.807968, 9.753143, 9.696899, 9.649567, 9.56987, 9.462387, 
    9.370392, 9.327942, 9.300278, 9.263367, 9.228912, 9.179321, 9.115448, 
    9.026764, 8.941803, 8.797211, 8.693237, 8.636551, 8.594681, 8.488815, 
    8.425858, 8.382507, 8.361282, 8.321365, 8.303329, 8.30014, 8.254837, 
    8.230942, 8.257843, 8.306335, 8.335831, 8.353668, 8.359329, 8.386597, 
    8.425018, 8.447601, 8.466293, 8.480103, 8.486542, 8.502045, 8.508881, 
    8.50769, 8.551331, 8.569946, 8.568695, 8.549118, 8.543121, 8.569351, 
    8.574173, 8.571182, 8.606995, 8.609451, 8.629059, 8.675735, 8.716034, 
    8.775604, 8.852676, 8.896439, 8.905884, 8.986862, 9.054901, 9.094208, 
    9.161987, 9.234268, 9.312653, 9.379242, 9.429321, 9.490128, 9.55014, 
    9.605759, 9.690964, 9.773712, 9.864929, 9.955414, 10.03432, 10.10576, 
    10.17261, 10.21635, 10.25522, 10.30959, 10.33817, 10.37932, 10.43668, 
    10.46211, 10.4545, 10.42442, 10.35002, 10.32613,
  3.033844, 3.013794, 2.997513, 2.982925, 2.97258, 2.959229, 2.946991, 
    2.938858, 2.943115, 2.947739, 2.953217, 2.959717, 2.959061, 2.957901, 
    2.945068, 2.92691, 2.8974, 2.861862, 2.819611, 2.777618, 2.733353, 
    2.686539, 2.647598, 2.615067, 2.588165, 2.56662, 2.550919, 2.541351, 
    2.544479, 2.557053, 2.577881, 2.600143, 2.62735, 2.657303, 2.685944, 
    2.718246, 2.74765, 2.789429, 2.832275, 2.872574, 2.904938, 2.939957, 
    2.975113, 3.006424, 3.036499, 3.061249, 3.068085, 3.086639, 3.100708, 
    3.108246, 3.116013, 3.123474, 3.10936, 3.07785, 3.150253, 3.154541, 
    3.177002, 3.170486, 3.2341, 3.218719, 3.233643, 3.264755, 3.287216, 
    3.363266, 3.436508, 3.51268, 3.582916, 3.656052, 3.702194, 3.712418, 
    3.72641, 3.733261, 3.741196, 3.808441, 3.694778, 3.658051, 3.635986, 
    3.60083, 3.557144, 3.507797, 3.478363, 3.455261, 3.434753, 3.409607, 
    3.391052, 3.367157, 3.343277, 3.315796, 3.282928, 3.249069, 3.21463, 
    3.186508, 3.157608, 3.126022, 3.095871, 3.062363,
  2.861053, 2.875702, 2.89888, 2.92691, 2.964539, 3.020386, 3.070724, 
    3.115051, 3.147156, 3.168442, 3.187057, 3.19371, 3.207642, 3.233612, 
    3.244751, 3.270401, 3.288422, 3.275986, 3.241104, 3.182693, 3.082108, 
    2.959198, 2.824371, 2.706528, 2.600998, 2.51474, 2.464737, 2.450867, 
    2.452698, 2.458542, 2.498322, 2.563614, 2.648453, 2.733643, 2.829346, 
    2.933182, 3.045746, 3.162216, 3.287872, 3.404022, 3.512939, 3.611572, 
    3.719833, 3.823425, 3.932144, 4.070755, 4.154907, 4.269653, 4.373108, 
    4.452789, 4.470749, 4.446259, 4.434998, 4.381042, 4.319778, 4.30069, 
    4.283829, 4.249283, 4.228287, 4.190018, 4.174316, 4.158066, 4.160339, 
    4.187744, 4.199921, 4.129211, 4.050705, 4.034882, 4.079544, 4.127655, 
    4.111893, 4.085464, 4.058319, 4.018356, 3.957275, 3.862549, 3.783051, 
    3.710587, 3.699982, 3.599396, 3.486313, 3.458832, 3.330124, 3.339172, 
    3.226288, 3.161438, 3.083908, 3.010208, 2.942947, 2.89679, 2.859421, 
    2.828949, 2.8255, 2.832336, 2.838715, 2.851944,
  2.64386, 2.8078, 3.003052, 3.15419, 3.244736, 3.243317, 3.225662, 3.210693, 
    3.197861, 3.182236, 3.185745, 3.210312, 3.197403, 3.146637, 3.104767, 
    3.101837, 3.152237, 3.182892, 3.185883, 3.147278, 3.072617, 2.985504, 
    2.845978, 2.621689, 2.395264, 2.316086, 2.394547, 2.565964, 2.677872, 
    2.694809, 2.719284, 2.753006, 2.78627, 2.815125, 2.83873, 2.858261, 
    2.888657, 2.972641, 3.064041, 3.170502, 3.288589, 3.431885, 3.58873, 
    3.78331, 4.011841, 4.125244, 4.148941, 4.162872, 4.255585, 4.464645, 
    4.477509, 4.397186, 4.359222, 4.266083, 4.072968, 3.884033, 3.712494, 
    3.476349, 3.302338, 3.175781, 3.181763, 3.246399, 3.34993, 3.363724, 
    3.362686, 3.423035, 3.501022, 3.643021, 3.800049, 3.910339, 4.006622, 
    4.026611, 3.982727, 3.973938, 3.972641, 3.968994, 3.950684, 3.92836, 
    3.829285, 3.755463, 3.691589, 3.638397, 3.592819, 3.4375, 3.300232, 
    3.219193, 3.143814, 3.075424, 2.983704, 2.85817, 2.725571, 2.58371, 
    2.488464, 2.467621, 2.47493, 2.529083,
  2.696335, 2.852188, 3.03862, 3.189667, 3.231201, 3.16597, 3.067734, 
    2.940247, 2.825989, 2.751907, 2.70639, 2.70047, 2.783035, 2.87442, 
    2.962021, 3.039703, 3.07193, 3.144638, 3.23085, 3.217682, 3.074066, 
    2.817551, 2.479477, 2.128204, 1.799683, 1.654572, 1.835297, 2.133209, 
    2.301117, 2.437973, 2.478073, 2.410629, 2.285568, 2.224747, 2.250092, 
    2.247543, 2.258911, 2.31926, 2.383057, 2.489304, 2.647125, 2.792755, 
    2.957672, 3.163727, 3.387405, 3.527466, 2.212189, 2.247498, 2.737274, 
    2.677704, 2.674103, 2.623016, 2.670288, 2.673981, 2.623657, 2.608307, 
    2.444214, 2.605072, 2.620636, 2.627686, 2.689941, 2.746063, 2.849457, 
    3.083328, 3.331238, 3.402588, 3.539108, 3.628815, 3.690674, 3.74556, 
    3.786957, 3.864517, 3.877777, 3.883896, 3.876007, 3.871399, 3.804138, 
    3.742294, 3.553772, 3.424377, 3.403931, 3.520905, 3.489471, 3.469025, 
    3.469086, 3.602081, 3.47403, 3.483368, 3.316833, 2.956848, 2.815979, 
    2.600449, 2.496994, 2.467957, 2.459946, 2.532654,
  1.983307, 2.062225, 2.273163, 2.453049, 2.548233, 2.514496, 2.511902, 
    2.511307, 2.590927, 2.534683, 2.580383, 2.630066, 2.734955, 2.872314, 
    2.768997, 2.55806, 2.457535, 2.344589, 2.130325, 2.228165, 2.328445, 
    2.169769, 2.019196, 1.967239, 1.975632, 1.933838, 1.979858, 2.050446, 
    2.170486, 2.291122, 2.340027, 2.313202, 2.240021, 2.152847, 2.15213, 
    2.188065, 2.26091, 2.341904, 2.205643, 2.031754, 1.985596, 2.112488, 
    2.253113, 2.324463, 2.370499, 2.380249, 2.194031, 1.500092, 1.088165, 
    0.812561, 0.7125549, 0.6399231, 0.6745605, 0.7897949, 0.9145203, 
    1.102356, 1.392151, 1.720123, 2.01181, 2.219147, 2.358612, 2.443237, 
    2.342346, 1.996094, 1.619659, 1.248779, 1.045258, 1.117523, 1.215454, 
    1.403534, 2.91571, 3.321503, 3.155029, 2.54007, 1.973114, 1.630737, 
    2.859924, 2.790771, 2.74231, 2.68869, 2.458405, 2.594086, 2.819885, 
    3.015961, 3.175323, 3.280792, 3.425232, 3.615662, 3.741669, 3.846832, 
    3.946381, 3.183746, 2.762207, 2.509125, 2.216721, 2.014954,
  2.289917, 1.894928, 2.412323, 2.201569, 1.948578, 1.777039, 1.812408, 
    2.006256, 2.10379, 2.183167, 2.294159, 2.305786, 2.370056, 2.359146, 
    2.233444, 2.039246, 1.880325, 1.721725, 1.56604, 1.440125, 1.35379, 
    1.275543, 1.301819, 1.390137, 1.560974, 1.630844, 1.726471, 1.760254, 
    1.867035, 1.929993, 1.891403, 1.859436, 1.79393, 1.616455, 1.541077, 
    1.398346, 1.212814, 1.078308, 0.9100952, 0.9989014, 1.114319, 1.222473, 
    1.160889, 1.01355, 0.851532, 0.4378357, 0.4665527, 0.264679, 0.03411865, 
    -0.04263306, -0.08352661, -0.08639526, -0.07797241, -0.04562378, 
    0.05456543, 0.2087402, 0.3892822, 0.5774536, 0.7164917, 0.8518372, 
    0.9902954, 1.125275, 1.156769, 1.089874, 0.9586792, 0.8688354, 0.8790588, 
    0.9202271, 1.026062, 1.217926, 1.353424, 1.371368, 1.231567, 1.004211, 
    0.815979, 0.7245483, 0.682312, 0.6857605, 1.793365, 1.992279, 2.121185, 
    2.292725, 2.341187, 2.433014, 2.537781, 2.707245, 2.888153, 3.013031, 
    3.257324, 3.538025, 3.677032, 3.735962, 3.726105, 3.636536, 3.403473, 
    2.954376,
  2.929504, 3.272552, 3.566284, 3.600616, 3.539551, 3.386108, 3.205811, 
    3.158813, 3.029572, 2.924774, 2.910309, 2.887451, 2.789368, 2.824188, 
    2.811951, 2.70639, 2.532837, 2.296234, 2.049164, 1.887817, 1.71637, 
    1.473206, 1.237915, 1.138489, 0.979187, 0.8583984, 0.6214905, 0.4649963, 
    0.3977966, 0.3809509, 0.3493958, 0.3197632, 0.3922119, 1.787109, 
    1.864746, 1.78952, 2.464691, 1.047852, 0.7713928, 0.6879272, 0.6355591, 
    0.62854, 0.618866, 0.5116272, 0.2774353, 0.04202271, -0.2114868, 
    -0.405304, -0.4749756, -0.456604, -0.3643494, -0.2722168, -0.2575073, 
    -0.289032, -0.29599, -0.2118835, -0.02185059, 0.1947327, 0.3848572, 
    0.5884399, 0.8235779, 0.996582, 1.092285, 1.12262, 1.138123, 1.197876, 
    1.283569, 1.319702, 1.285278, 1.222443, 1.191833, 1.203003, 1.183777, 
    1.164429, 1.112732, 1.012787, 0.9151306, 0.9658508, 1.429352, 2.208496, 
    2.236298, 1.803375, 1.571991, 1.498535, 1.565186, 1.730499, 1.965546, 
    2.128998, 2.235779, 2.300537, 2.35672, 2.385956, 2.436798, 2.469238, 
    2.521515, 2.710388,
  1.532074, 1.510254, 1.422638, 1.333405, 1.256439, 1.20285, 1.229401, 
    1.303284, 1.326019, 1.341492, 1.404602, 1.548065, 1.670807, 1.702637, 
    1.690979, 1.673218, 1.673096, 1.663269, 1.587006, 1.443268, 1.309265, 
    1.167542, 1.048615, 0.9757996, 0.9552307, 0.864502, 0.679718, 0.5116882, 
    0.4054565, 0.3713074, 0.3330383, 0.3228149, 0.3790894, 0.480835, 
    0.6357117, 0.7924194, 0.9418335, 0.8930054, 0.8132935, 0.822876, 
    0.8719177, 0.9124756, 0.9085693, 0.860199, 0.6963806, 0.4234009, 
    -0.02093506, -0.3808289, -0.5285645, -0.6275635, -0.7234192, -0.7463989, 
    -0.6918945, -0.6231384, -0.5141602, -0.3211975, -0.07504272, 0.144165, 
    0.2835693, 0.4915161, 0.7817993, 1.017944, 1.107697, 1.195557, 1.38089, 
    1.548859, 1.688446, 1.76886, 1.778198, 1.77243, 1.830841, 1.906219, 
    1.930389, 1.930817, 1.898987, 1.772278, 1.61676, 1.513916, 1.495209, 
    1.556213, 1.664032, 1.583496, 1.266571, 1.046783, 1.128052, 1.248596, 
    1.417816, 1.551392, 1.628723, 1.675598, 1.672363, 1.644958, 1.633514, 
    1.608124, 1.575623, 1.54776,
  1.408051, 1.310516, 1.219971, 1.103302, 1.004272, 0.9474487, 0.9814148, 
    1.000214, 1.017944, 1.040131, 1.111298, 1.240021, 1.347473, 1.431335, 
    1.491028, 1.536316, 1.583099, 1.601471, 1.530182, 1.380493, 1.304596, 
    1.202759, 1.059235, 1.017029, 1.079346, 1.072998, 1.0047, 0.9263306, 
    0.8531494, 0.758606, 0.6191711, 0.4832153, 0.3860168, 0.3432617, 
    0.3357239, 0.3488159, 0.4251404, 0.6446838, 0.9092712, 1.097748, 
    1.149963, 1.173004, 1.251801, 1.170715, 0.9957886, 0.8676758, 0.6681824, 
    0.287384, -0.1815491, -0.5282288, -0.6703491, -0.7063599, -0.6428528, 
    -0.5675964, -0.4945679, -0.2956543, -0.005889893, 0.18396, 0.217804, 
    0.3378601, 0.7293396, 1.042847, 1.141479, 1.270142, 1.566833, 1.808502, 
    1.914795, 1.970795, 2.007141, 2.043701, 2.081818, 2.080902, 2.075439, 
    2.080963, 2.016449, 1.843781, 1.573853, 1.450623, 1.482269, 1.604919, 
    1.731354, 1.860657, 1.738251, 1.364868, 1.047302, 1.014679, 1.184143, 
    1.308228, 1.382263, 1.424896, 1.515594, 1.539093, 1.497437, 1.513092, 
    1.514374, 1.490479,
  1.510834, 1.567535, 1.600891, 1.594604, 1.585266, 1.598145, 1.63858, 
    1.582245, 1.518158, 1.520721, 1.552399, 1.622284, 1.66156, 1.72113, 
    1.853424, 1.967621, 2.119629, 2.253479, 2.180176, 1.836731, 1.637756, 
    1.506989, 1.263245, 1.106873, 1.145813, 1.236481, 1.264771, 1.270081, 
    1.261078, 1.196777, 1.09967, 1.002319, 0.9066772, 0.8047485, 0.7459412, 
    0.7702942, 0.8420715, 0.9840393, 1.168854, 1.251709, 1.263184, 1.329773, 
    1.403107, 1.32019, 1.199829, 1.164459, 1.08371, 0.785614, 0.2974854, 
    -0.008972168, -0.02642822, 0.05410767, 0.09811401, 0.1146545, 0.1567688, 
    0.2674561, 0.3988342, 0.4950256, 0.5299377, 0.6738892, 0.946106, 
    1.148834, 1.269867, 1.455719, 1.721313, 1.791046, 1.750977, 1.833893, 
    1.923401, 1.91922, 1.898254, 1.949097, 2.001129, 1.964111, 1.776367, 
    1.438538, 1.349854, 1.801178, 1.814453, 1.510162, 1.46994, 1.513702, 
    1.518585, 1.207672, 1.010254, 1.264099, 1.577423, 1.746826, 1.731812, 
    1.666626, 1.67691, 1.69632, 1.694031, 1.679779, 1.622375, 1.544495,
  1.990906, 2.032898, 2.104858, 2.167999, 2.217041, 2.244049, 2.266693, 
    2.275818, 2.242737, 2.271271, 2.380676, 2.457397, 2.468964, 2.498291, 
    2.54834, 2.594238, 2.749847, 2.956207, 2.936432, 2.680756, 2.53598, 
    2.49231, 2.242218, 1.900879, 1.739288, 1.787292, 1.836548, 1.780823, 
    1.666046, 1.544891, 1.453308, 1.41037, 1.350739, 1.216461, 1.118744, 
    1.081421, 1.119324, 1.191467, 1.291138, 1.430084, 1.527679, 1.550659, 
    1.516602, 1.47525, 1.484833, 1.505066, 1.390839, 1.173218, 0.836853, 
    0.6345825, 0.6621094, 0.785675, 0.8551636, 0.8718262, 0.8943176, 
    0.9503784, 0.9937439, 1.066345, 1.144989, 1.242767, 1.37558, 1.470001, 
    1.577332, 1.692627, 1.799805, 1.819855, 1.794983, 1.843109, 1.92923, 
    1.895691, 1.805725, 1.798523, 1.777557, 1.660675, 1.497742, 1.399933, 
    1.808014, 2.026825, 1.786194, 1.812164, 1.652283, 1.413025, 1.190399, 
    1.032959, 1.206726, 1.550751, 1.811798, 1.99881, 2.074951, 2.073212, 
    2.07251, 2.05484, 2.034607, 2.051483, 2.081543, 2.022797,
  2.115295, 2.172119, 2.280334, 2.3349, 2.385742, 2.473297, 2.644318, 
    2.805573, 2.847595, 2.908997, 3.062714, 3.198395, 3.29007, 3.301788, 
    3.193909, 3.079529, 3.113892, 3.260529, 3.278748, 3.299469, 3.382568, 
    3.28418, 2.898315, 2.521545, 2.346344, 2.296997, 2.253265, 2.05957, 
    1.798157, 1.611938, 1.575836, 1.608459, 1.597015, 1.523315, 1.441925, 
    1.410095, 1.442902, 1.460266, 1.437805, 1.542236, 1.814056, 1.87793, 
    1.809296, 1.829712, 1.968628, 2.130798, 2.072632, 1.864441, 1.586243, 
    1.480316, 1.650726, 1.784454, 1.794983, 1.715607, 1.590302, 1.568176, 
    1.605286, 1.6875, 1.728973, 1.74173, 1.752014, 1.791595, 1.859772, 
    1.869019, 1.894623, 1.946411, 1.946564, 1.914063, 1.900391, 1.834198, 
    1.70163, 1.636719, 1.57135, 1.479034, 1.419861, 1.418427, 1.83255, 
    2.234314, 2.684174, 2.023163, 1.716919, 1.3927, 1.182281, 1.248718, 
    1.637177, 1.98288, 2.094025, 2.135803, 2.208191, 2.214325, 2.183746, 
    2.192261, 2.18924, 2.171997, 2.166992, 2.135406,
  2.289703, 2.320618, 2.433777, 2.564514, 2.730194, 3.076874, 3.503601, 
    3.757019, 3.913696, 4.11264, 4.263611, 4.193481, 3.923431, 3.665741, 
    3.445892, 3.34021, 3.279083, 3.207794, 3.225861, 3.306763, 3.241943, 
    2.890411, 2.472534, 2.243042, 2.155212, 2.132874, 2.1362, 2.004578, 
    1.889648, 1.876556, 1.915253, 1.931427, 1.901367, 1.812317, 1.795776, 
    1.859497, 1.858063, 1.738403, 1.681, 2.006775, 2.512878, 2.517303, 
    2.384644, 2.377808, 2.449677, 2.589386, 2.789581, 2.561584, 2.486908, 
    2.505402, 2.611053, 2.524475, 2.349915, 2.167145, 2.011536, 1.996033, 
    2.025269, 2.005402, 1.980804, 1.96347, 1.929962, 1.936401, 1.95105, 
    2.002808, 2.019073, 2.018158, 2.022217, 1.926697, 1.828247, 1.783478, 
    1.723694, 1.666534, 1.615173, 1.53949, 1.463348, 1.357605, 1.662689, 
    3.365234, 4.054749, 2.266724, 1.827728, 1.69928, 1.800781, 2.02005, 
    2.222992, 2.370392, 2.368164, 2.300446, 2.267639, 2.263062, 2.254028, 
    2.277924, 2.278778, 2.269135, 2.295898, 2.294312,
  2.063019, 2.109253, 2.276062, 2.54245, 2.896393, 3.331055, 3.642059, 
    4.169647, 4.311981, 3.956299, 3.439392, 3.010559, 2.683655, 2.471161, 
    2.412567, 2.565887, 2.650452, 2.616669, 2.56778, 2.417267, 2.245117, 
    2.110565, 2.000336, 1.958923, 1.938141, 1.969086, 2.034393, 2.020874, 
    2.089203, 2.218506, 2.202209, 2.143616, 2.089142, 1.997986, 2.100525, 
    2.144867, 2.039398, 2.070435, 2.444977, 3.684448, 2.976715, 3.07962, 
    3.217316, 3.049011, 2.914703, 2.953247, 3.071167, 3.346954, 2.770264, 
    2.606781, 2.527405, 2.468231, 2.38385, 2.356781, 2.276733, 2.218353, 
    2.126221, 2.030548, 2.036987, 2.026154, 2.014313, 2.050903, 2.028442, 
    2.057404, 2.080475, 2.05014, 2.072906, 2.038605, 1.927979, 1.86554, 
    1.785614, 1.739471, 1.668091, 1.542572, 1.482269, 1.346558, 1.518036, 
    3.499725, 3.663239, 2.204956, 1.706573, 1.915955, 2.225708, 2.431305, 
    2.429108, 2.410919, 2.386658, 2.37149, 2.3909, 2.371796, 2.316132, 
    2.278961, 2.213043, 2.139862, 2.054291, 2.040222,
  1.930206, 1.914001, 2.013916, 2.168671, 2.372833, 2.585785, 2.860565, 
    3.037964, 2.844055, 2.427673, 1.841858, 1.85965, 1.87616, 1.946533, 
    1.968872, 2.062378, 2.101898, 2.013062, 1.952728, 1.858978, 1.824219, 
    1.883728, 1.864197, 1.902161, 1.882355, 1.960876, 2.089447, 2.132477, 
    2.292786, 2.322784, 2.116913, 2.162109, 2.048035, 1.917877, 1.994781, 
    2.001556, 2.093872, 3.348511, 3.961639, 4.152802, 3.297974, 2.903839, 
    3.610626, 3.377228, 3.106812, 3.118378, 2.970978, 2.704559, 2.350067, 
    2.061218, 2.092896, 2.124634, 2.139984, 2.136139, 2.107819, 2.118896, 
    2.065887, 2.066742, 2.132751, 2.142456, 2.127014, 2.164307, 2.185791, 
    2.177124, 2.164978, 2.091614, 2.054169, 1.973114, 1.853729, 1.77063, 
    1.642487, 1.595245, 1.531586, 1.327911, 1.254761, 1.180878, 1.439178, 
    3.456299, 3.605652, 1.67804, 1.189697, 1.814056, 2.185608, 2.330078, 
    2.237518, 2.184448, 2.205597, 2.259155, 2.344391, 2.279816, 2.183655, 
    2.139771, 2.065674, 2.019012, 1.95517, 1.933319,
  1.688568, 1.671295, 1.665802, 1.819855, 2.214844, 3.93924, 3.920258, 
    3.496246, 2.91275, 2.055237, 2.051575, 2.287018, 2.253632, 2.26828, 
    2.22403, 2.194092, 2.288818, 2.227081, 2.16687, 2.11673, 2.145386, 
    2.147064, 2.128326, 2.164886, 2.17865, 2.195526, 2.271362, 2.251892, 
    2.146545, 1.858978, 1.963806, 3.315094, 3.476044, 3.185669, 3.419922, 
    3.488281, 4.030334, 3.894867, 3.709595, 3.377075, 2.49472, 2.333984, 
    2.141083, 2.124207, 2.382416, 2.524292, 2.305603, 1.945129, 1.88385, 
    2.032104, 2.115692, 2.153717, 2.205322, 2.165436, 2.083771, 2.031433, 
    2.022919, 2.055725, 2.095367, 2.132294, 2.090881, 2.060333, 2.076874, 
    2.03952, 1.992188, 1.860046, 1.751495, 1.627533, 1.510071, 1.418427, 
    1.304962, 1.217712, 1.154755, 1.113403, 1.028076, 1.031067, 1.372009, 
    2.736511, 3.738861, 2.394806, 2.175842, 2.370941, 2.217255, 2.301361, 
    2.203827, 2.202148, 2.314636, 2.328064, 2.362823, 2.279022, 2.202087, 
    2.051453, 1.928314, 1.889832, 1.83548, 1.765839,
  1.522552, 1.534058, 1.750763, 2.049225, 2.59668, 3.839203, 3.818939, 
    3.082947, 2.662262, 2.077362, 1.991547, 2.180023, 2.130737, 2.243164, 
    2.42157, 2.490479, 2.53595, 2.51712, 2.436981, 2.372528, 2.288239, 
    2.241882, 2.172943, 2.08197, 2.02005, 1.941193, 1.894867, 1.91568, 
    1.99765, 2.002594, 2.446686, 3.784973, 3.913147, 3.527649, 3.471924, 
    3.701752, 4.078125, 3.548248, 2.767731, 2.455292, 2.030945, 1.988647, 
    1.512299, 1.602295, 1.927155, 2.108673, 2.147125, 2.108002, 2.145386, 
    2.230713, 2.208374, 2.164734, 2.133484, 2.040497, 2.006378, 1.982086, 
    1.953064, 1.953705, 1.878784, 1.860107, 1.817841, 1.766479, 1.735138, 
    1.619232, 1.564575, 1.417511, 1.322266, 1.200195, 1.092499, 1.086578, 
    1.021149, 1.064453, 0.9993286, 1.022858, 0.9207764, 1.212708, 1.742767, 
    2.709106, 4.240448, 2.960785, 2.237885, 2.776093, 2.615173, 2.638031, 
    2.347473, 2.272766, 2.327545, 2.282623, 2.213257, 2.117126, 2.030487, 
    1.921295, 1.858521, 1.772186, 1.661835, 1.582825,
  1.668549, 1.871735, 2.18158, 2.574615, 3.314056, 3.846558, 3.794678, 
    3.411255, 3.341339, 3.20755, 2.160828, 2.237366, 2.442078, 2.212891, 
    2.275055, 2.371094, 2.268097, 2.13385, 2.043732, 1.993744, 1.902679, 
    1.87677, 1.882813, 1.865875, 1.880219, 1.886353, 1.926819, 2.071747, 
    2.228394, 2.255096, 2.612244, 3.958069, 4.158081, 3.625824, 3.604675, 
    3.877014, 3.643555, 2.865479, 2.530212, 2.004211, 1.481567, 1.937042, 
    1.920258, 2.111542, 2.171295, 2.214447, 2.2901, 2.267303, 2.216156, 
    2.172394, 2.139404, 2.102356, 2.085144, 2.028839, 2.017853, 1.985809, 
    1.895081, 1.868103, 1.844849, 1.776581, 1.672546, 1.555603, 1.52298, 
    1.395691, 1.282166, 1.138336, 1.042511, 0.986145, 1.014648, 1.05545, 
    1.047577, 1.050964, 0.9614563, 1.038147, 1.100067, 1.638062, 2.298096, 
    3.263214, 5.366333, 3.294739, 1.750061, 2.790039, 2.969574, 2.690613, 
    2.453766, 2.322113, 2.231201, 2.169922, 2.018951, 1.846924, 1.756439, 
    1.698242, 1.674072, 1.657227, 1.633911, 1.638458,
  2.059692, 2.314178, 2.473297, 2.69693, 3.699341, 3.47052, 3.381165, 
    3.549805, 3.60144, 3.041412, 2.274261, 2.180847, 2.403107, 2.726105, 
    2.305664, 2.277466, 2.13092, 2.025055, 2.014923, 2.004608, 1.969727, 
    1.942383, 1.986572, 1.984711, 2.002289, 2.094452, 2.270325, 2.445496, 
    2.516663, 2.461975, 2.454559, 2.774872, 3.848633, 3.897919, 3.676056, 
    3.49057, 3.218384, 2.70401, 2.512238, 1.878571, 2.030975, 2.056519, 
    2.124146, 2.170258, 2.154572, 2.191925, 2.202026, 2.187653, 2.160675, 
    2.128754, 2.096985, 2.060028, 2.047058, 2.068634, 2.060883, 2.072601, 
    2.021088, 1.944153, 1.926697, 1.84317, 1.78125, 1.690247, 1.589783, 
    1.424103, 1.287048, 1.227142, 1.217896, 1.228302, 1.241791, 1.29895, 
    1.278381, 1.296814, 1.299133, 1.473907, 1.518097, 1.840637, 2.399475, 
    3.506256, 4.697601, 3.123627, 1.922974, 2.815948, 3.047516, 2.863678, 
    2.856964, 3.18808, 2.155457, 2.044189, 1.936584, 1.777069, 1.759491, 
    1.751221, 1.82077, 1.823517, 1.898438, 1.967896,
  2.520325, 2.702271, 2.776672, 2.630341, 3.277283, 3.079163, 2.947083, 
    3.147217, 3.198975, 2.531372, 2.765778, 2.408661, 2.384247, 2.480133, 
    2.358612, 2.358765, 2.240173, 2.176239, 2.191986, 2.201569, 2.185242, 
    2.191132, 2.196136, 2.201477, 2.276825, 2.390869, 2.527405, 2.612488, 
    2.594391, 2.54837, 2.446167, 2.453796, 2.632996, 3.657623, 3.335083, 
    2.655518, 2.642181, 2.418488, 2.563019, 2.044647, 2.044403, 2.150574, 
    2.195313, 2.184357, 2.164307, 2.161591, 2.107147, 2.184296, 2.236969, 
    2.224731, 2.197723, 2.154877, 2.133545, 2.123047, 2.141754, 2.12149, 
    2.106201, 2.083069, 2.072266, 1.970703, 1.9487, 1.865448, 1.772766, 
    1.693115, 1.649933, 1.641937, 1.618805, 1.680969, 1.689697, 1.722656, 
    1.70105, 1.726227, 1.758392, 1.831451, 1.804169, 2.255585, 3.714294, 
    4.735992, 3.555084, 2.864838, 2.651825, 2.779114, 2.823029, 2.858978, 
    3.181885, 3.364502, 2.105255, 2.119904, 2.030396, 2.007935, 2.044189, 
    2.098053, 2.201935, 2.260742, 2.331116, 2.452545,
  2.761505, 2.817169, 2.724609, 2.388672, 2.937439, 2.771881, 2.821594, 
    2.91568, 2.640167, 2.550262, 2.55545, 2.46048, 2.283203, 2.391205, 
    2.37207, 2.338928, 2.30957, 2.283783, 2.296814, 2.347473, 2.366547, 
    2.397339, 2.371368, 2.374786, 2.43515, 2.459564, 2.547577, 2.616302, 
    2.528442, 2.428375, 2.446991, 2.46994, 2.451904, 2.305359, 2.29068, 
    2.693359, 2.794983, 2.304565, 2.068085, 2.141998, 2.136414, 2.232422, 
    2.212372, 2.115326, 2.044159, 2.012177, 1.9505, 2.012512, 2.13855, 
    2.160156, 2.159973, 2.119354, 2.172913, 2.204163, 2.226318, 2.184113, 
    2.225861, 2.236389, 2.215302, 2.169647, 2.168396, 2.118744, 2.080597, 
    2.072784, 2.026367, 2.026154, 2.041077, 2.089233, 2.075775, 2.141754, 
    2.178375, 2.265839, 2.375916, 2.313873, 2.325653, 3.035095, 3.196869, 
    3.157227, 2.989197, 2.723297, 2.829742, 2.938995, 3.025665, 2.887634, 
    2.93573, 2.791931, 2.136261, 2.246094, 2.267761, 2.274597, 2.325043, 
    2.42981, 2.478729, 2.567841, 2.655548, 2.724304,
  2.789246, 2.757538, 2.526886, 2.31601, 2.831635, 2.889282, 2.804291, 
    2.876801, 2.868805, 2.715302, 2.536987, 2.417511, 2.374939, 2.40448, 
    2.365112, 2.26712, 2.355682, 2.437317, 2.445984, 2.506317, 2.492584, 
    2.518677, 2.51712, 2.481964, 2.468445, 2.416016, 2.399078, 2.347198, 
    2.398804, 2.399933, 2.349609, 2.411377, 2.489258, 2.433411, 2.371033, 
    2.294922, 2.146698, 2.199493, 2.528473, 2.163269, 2.047485, 2.144012, 
    2.163605, 2.052948, 1.974396, 1.926758, 1.940643, 1.994659, 2.126617, 
    2.121552, 2.205139, 2.214111, 2.249542, 2.28717, 2.276154, 2.265045, 
    2.28418, 2.282349, 2.287415, 2.334656, 2.330078, 2.347992, 2.309631, 
    2.305603, 2.274292, 2.26297, 2.29303, 2.320648, 2.382294, 2.456757, 
    2.56369, 2.602875, 2.618103, 2.552734, 2.531342, 2.750061, 3.02063, 
    3.073639, 3.09845, 3.051056, 3.017212, 2.950439, 3.043945, 3.248566, 
    2.918549, 2.592499, 3.169983, 2.320709, 2.379272, 2.402863, 2.418182, 
    2.49472, 2.529694, 2.643677, 2.735535, 2.763153,
  2.484924, 2.480988, 2.316742, 2.377228, 3.539825, 3.402802, 3.132721, 
    3.084381, 2.779877, 2.300079, 1.758087, 2.44455, 2.437683, 2.474731, 
    2.490112, 2.408905, 2.41745, 2.494263, 2.52652, 2.519104, 2.494537, 
    2.515564, 2.491211, 2.495575, 2.504028, 2.500885, 2.404572, 2.337433, 
    2.503448, 2.471222, 2.358826, 2.29129, 2.416321, 2.372345, 2.362427, 
    2.472992, 2.299347, 2.632385, 2.740234, 2.72879, 1.954102, 2.183777, 
    2.288239, 2.222717, 2.13208, 2.114441, 2.203888, 2.226288, 2.319916, 
    2.334686, 2.383911, 2.437378, 2.443939, 2.478119, 2.512238, 2.519073, 
    2.486847, 2.469025, 2.4664, 2.488983, 2.486267, 2.480377, 2.473114, 
    2.453796, 2.451569, 2.428192, 2.464142, 2.480225, 2.551025, 2.589386, 
    2.635223, 2.619781, 2.580078, 2.664063, 2.641541, 2.623047, 2.880585, 
    3.218292, 3.305084, 3.148376, 3.26236, 3.114197, 3.14798, 3.843689, 
    3.282166, 2.639069, 3.252136, 2.364014, 2.422974, 2.440887, 2.527527, 
    2.565247, 2.567902, 2.600403, 2.588806, 2.546875,
  2.359619, 2.370422, 2.354034, 2.917786, 3.521851, 3.375519, 3.170441, 
    3.097015, 2.965424, 2.119781, 1.563263, 2.872528, 2.502747, 2.52655, 
    2.566345, 2.506195, 2.492645, 2.424347, 2.445374, 2.473511, 2.478638, 
    2.501312, 2.488922, 2.470825, 2.468872, 2.467102, 2.429169, 2.717834, 
    2.655914, 2.378723, 2.650146, 2.579956, 2.491394, 2.18399, 2.263855, 
    2.844543, 2.474915, 2.122711, 1.96225, 1.992706, 2.092712, 2.167847, 
    2.161407, 2.137115, 2.161469, 2.118042, 2.116272, 2.121033, 2.168884, 
    2.204773, 2.199219, 2.230011, 2.266785, 2.305206, 2.320709, 2.338867, 
    2.384583, 2.435791, 2.46048, 2.510223, 2.56076, 2.589783, 2.643677, 
    2.694855, 2.767975, 2.822662, 2.897797, 2.955658, 2.930481, 2.954315, 
    2.931854, 2.823639, 2.689545, 2.603821, 2.644592, 2.738281, 2.514862, 
    2.807373, 3.094971, 3.02832, 3.064972, 4.010742, 3.973694, 4.369812, 
    3.59848, 2.301178, 2.325775, 2.363464, 2.448517, 2.457245, 2.509491, 
    2.458923, 2.505676, 2.49646, 2.472198, 2.410675,
  2.399811, 2.535339, 2.515106, 3.157898, 3.530151, 3.520386, 3.303833, 
    3.21991, 2.881104, 2.262451, 2.006531, 3.460815, 2.890167, 2.494598, 
    2.512756, 2.611969, 2.552673, 2.511841, 2.517059, 2.516266, 2.515686, 
    2.492462, 2.506134, 2.53595, 2.497528, 2.40332, 2.392761, 2.973053, 
    2.29895, 2.389771, 2.658997, 2.419037, 2.302216, 2.257141, 2.185608, 
    2.180542, 2.041077, 2.036591, 2.100006, 2.159485, 2.166229, 2.152802, 
    2.139343, 2.129669, 2.113495, 2.111267, 2.103882, 2.088623, 2.088867, 
    2.111084, 2.119965, 2.146027, 2.177277, 2.194, 2.208588, 2.196411, 
    2.200256, 2.20871, 2.255219, 2.260437, 2.279114, 2.343567, 2.43515, 
    2.540314, 2.655487, 2.749481, 2.856964, 2.976379, 3.064392, 3.061066, 
    2.948181, 2.788483, 2.654938, 2.514008, 2.314758, 2.429382, 2.758728, 
    2.646484, 2.521149, 3.115753, 3.689514, 3.93869, 3.464966, 2.236542, 
    2.133057, 2.138153, 2.208862, 2.293823, 2.358002, 2.415405, 2.499023, 
    2.533539, 2.551514, 2.46817, 2.482147, 2.385864,
  3.373688, 2.783325, 3.320679, 3.571686, 3.307617, 3.53833, 3.693237, 
    3.529816, 3.236176, 3.411591, 2.658478, 2.533356, 3.069244, 2.539764, 
    2.552155, 2.664856, 2.632629, 2.636017, 2.599487, 2.575195, 2.527466, 
    2.510406, 2.461731, 2.495636, 2.522125, 2.552032, 2.947388, 2.963409, 
    2.226318, 2.275726, 2.323975, 2.44101, 2.233124, 2.368744, 2.12442, 
    2.088654, 2.107605, 2.139038, 2.176819, 2.228638, 2.241669, 2.258087, 
    2.256989, 2.292053, 2.327057, 2.379761, 2.41568, 2.437164, 2.485626, 
    2.504028, 2.506195, 2.495239, 2.503845, 2.497009, 2.505402, 2.473328, 
    2.447723, 2.417664, 2.364136, 2.335083, 2.294556, 2.268494, 2.26413, 
    2.297272, 2.308777, 2.392395, 2.517365, 2.674347, 2.885834, 2.938538, 
    2.888489, 2.712616, 2.536072, 2.442047, 2.396912, 2.590485, 3.130798, 
    3.768555, 3.569397, 4.423981, 3.764862, 3.216614, 2.497406, 2.136902, 
    2.154663, 2.182098, 2.254547, 2.289185, 2.353271, 2.439789, 2.509827, 
    2.524231, 2.501373, 2.529877, 3.28186, 3.282837,
  3.193481, 2.897003, 3.376587, 3.143097, 3.199677, 3.590942, 3.313782, 
    3.331909, 3.280945, 3.666656, 3.314911, 3.04187, 3.337952, 3.194794, 
    2.51178, 2.632996, 2.823853, 2.802612, 2.795074, 2.751434, 2.763733, 
    3.146484, 2.598969, 2.51004, 2.449219, 2.370758, 2.473297, 3.120331, 
    2.315552, 2.237366, 2.261017, 2.146332, 2.184906, 2.684845, 2.240936, 
    2.19693, 2.261902, 2.269409, 2.314453, 2.334625, 2.350128, 2.376373, 
    2.378723, 2.3927, 2.418304, 2.460754, 2.485992, 2.506042, 2.54126, 
    2.587219, 2.650696, 2.69635, 2.727661, 2.788208, 2.832825, 2.795166, 
    2.764984, 2.711914, 2.61496, 2.562775, 2.505859, 2.45343, 2.460358, 
    2.451843, 2.432007, 2.435028, 2.469543, 2.611969, 2.821472, 2.874847, 
    2.765442, 2.644135, 2.833771, 2.916168, 2.886322, 3.358673, 4.065552, 
    4.389465, 3.7211, 3.356964, 2.283722, 2.260834, 2.356567, 2.263397, 
    2.210297, 2.197968, 2.243042, 2.291992, 2.339996, 2.379028, 2.460419, 
    2.535858, 2.653778, 3.319214, 3.563202, 3.313568,
  3.45871, 3.124603, 2.99649, 2.676361, 2.379303, 2.557465, 2.616211, 
    2.582031, 2.837708, 3.567444, 4.034821, 4.199738, 3.663208, 3.478119, 
    2.59726, 2.558136, 2.737946, 2.819397, 2.968597, 2.933716, 4.511932, 
    4.656372, 2.706268, 2.601624, 2.463043, 2.288818, 2.288208, 3.206177, 
    3.416412, 2.691467, 2.187378, 2.204041, 2.189453, 2.714386, 2.203064, 
    2.261841, 2.313721, 2.295959, 2.325928, 2.303131, 2.316406, 2.314789, 
    2.336639, 2.328125, 2.3638, 2.389587, 2.396393, 2.453064, 2.483551, 
    2.542572, 2.607025, 2.641724, 2.678467, 2.736206, 2.793121, 2.811462, 
    2.821411, 2.798767, 2.711121, 2.613129, 2.539063, 2.511078, 2.482147, 
    2.460541, 2.449677, 2.420258, 2.390808, 2.49231, 2.65567, 2.779236, 
    2.774933, 2.811584, 3.888489, 4.131317, 2.615021, 2.705933, 2.622772, 
    2.446716, 2.375244, 2.357056, 2.289459, 2.300781, 2.232605, 2.200897, 
    2.187897, 2.23587, 2.252472, 2.329407, 2.351166, 2.388, 2.484894, 
    2.769928, 3.433655, 3.775696, 3.659821, 3.473816,
  3.60495, 3.294678, 2.928009, 2.721771, 2.495453, 2.388977, 2.351227, 
    2.30722, 2.609039, 3.017395, 3.87793, 4.288849, 3.391144, 3.054565, 
    3.352997, 2.699219, 2.622314, 2.654358, 2.855408, 2.813416, 4.878967, 
    5.359772, 2.924652, 2.753845, 2.601379, 2.526245, 3.412506, 2.474762, 
    2.191803, 1.79599, 2.080017, 2.111023, 1.946198, 1.92395, 2.033142, 
    2.110535, 2.162506, 2.171997, 2.185455, 2.180023, 2.214905, 2.196075, 
    2.230011, 2.212433, 2.207489, 2.231964, 2.240692, 2.253448, 2.295044, 
    2.350403, 2.424866, 2.529572, 2.609497, 2.664703, 2.662537, 2.681, 
    2.687195, 2.648193, 2.529236, 2.416626, 2.282959, 2.178772, 2.179169, 
    2.244995, 2.299103, 2.253906, 2.108978, 2.090729, 2.371735, 3.988464, 
    4.149353, 4.227264, 3.146729, 2.297974, 2.440308, 2.484375, 2.456055, 
    2.45697, 2.393433, 2.324158, 2.240173, 2.159058, 2.073761, 2.017578, 
    1.994995, 2.020233, 2.052734, 2.155396, 2.22467, 2.320648, 2.434509, 
    2.911743, 4.185547, 4.205078, 4.329041, 3.992493,
  3.910583, 3.586029, 3.300659, 3.044403, 2.863403, 2.691406, 2.690216, 
    2.671722, 2.820129, 2.749237, 2.29361, 3.910675, 3.456329, 3.112396, 
    3.533539, 3.589447, 2.690643, 2.678925, 2.836975, 2.761139, 4.709839, 
    4.52713, 4.356384, 4.451813, 2.85379, 3.992523, 4.040894, 2.70813, 
    1.441925, 1.434906, 2.003845, 2.151428, 1.968689, 1.884491, 1.834198, 
    1.818726, 1.871765, 1.902222, 1.937775, 1.916992, 1.947784, 1.956757, 
    1.971344, 1.991608, 1.988983, 2.042725, 2.086334, 2.119415, 2.190613, 
    2.218353, 2.285492, 2.364319, 2.415222, 2.472351, 2.516602, 2.542328, 
    2.516663, 2.481842, 2.39386, 2.243408, 2.071442, 1.89035, 1.769257, 
    1.800446, 1.946747, 2.003845, 1.897064, 2.098053, 3.423065, 3.254364, 
    2.704163, 2.403198, 2.055542, 2.012115, 2.284637, 2.378845, 2.448364, 
    2.511719, 2.476227, 2.396698, 2.320679, 2.22995, 2.110565, 1.983185, 
    1.9328, 1.91333, 1.897003, 1.935242, 1.890686, 1.915314, 2.066589, 
    2.687439, 4.329285, 4.18576, 4.286469, 4.293304,
  4.292267, 4.0961, 3.612762, 3.389038, 3.09552, 2.649078, 2.617523, 
    2.707092, 2.872864, 3.178711, 2.13205, 3.718414, 3.290314, 3.321869, 
    3.578033, 3.483582, 2.806122, 2.980591, 4.418152, 4.432098, 4.366455, 
    3.63559, 4.081909, 3.906006, 3.728973, 3.909607, 4.119141, 3.231445, 
    1.729065, 1.414948, 1.868744, 2.354126, 2.074402, 1.952148, 1.937683, 
    1.913849, 1.957886, 1.968567, 1.963989, 1.942841, 1.944641, 1.960175, 
    1.905029, 1.888611, 1.836853, 1.787384, 1.751251, 1.763031, 1.7966, 
    1.832153, 1.940094, 2.063538, 2.168823, 2.217468, 2.245758, 2.34256, 
    2.366028, 2.366608, 2.358856, 2.304626, 2.203583, 2.06543, 1.914276, 
    1.882813, 1.991394, 1.897156, 2.150391, 3.57486, 3.458282, 2.868927, 
    2.883972, 2.226257, 1.860504, 1.903687, 1.996033, 2.106506, 2.222534, 
    2.378693, 2.602539, 2.576477, 2.516083, 2.47525, 2.420624, 2.324921, 
    2.23587, 2.107635, 2.030334, 1.99942, 1.914825, 1.922211, 2.04538, 
    2.358398, 3.865173, 4.136841, 4.168762, 4.299713,
  3.926575, 4.070038, 3.727875, 3.512939, 3.273743, 2.654541, 2.74231, 
    2.782166, 2.889832, 3.321442, 3.34201, 3.114563, 3.141479, 3.574554, 
    3.911957, 3.656494, 3.465912, 4.472473, 4.976013, 4.706635, 5.026672, 
    4.839355, 4.348145, 4.091125, 2.777893, 3.424377, 3.724121, 3.234009, 
    2.668915, 3.289886, 3.457001, 3.143311, 2.922302, 2.088989, 2.044556, 
    2.004486, 2.044006, 2.109375, 2.096741, 2.04068, 1.968231, 1.956665, 
    1.916992, 1.874084, 1.794006, 1.740662, 1.727203, 1.716431, 1.700836, 
    1.662109, 1.700073, 1.733063, 1.799561, 1.877075, 1.973969, 2.122925, 
    2.217377, 2.23053, 2.189056, 2.218658, 2.15332, 2.041595, 1.964783, 
    1.967133, 1.948242, 2.10553, 3.799683, 3.888245, 3.113922, 3.171631, 
    3.132935, 2.511353, 2.229248, 2.227661, 1.78952, 1.991669, 2.102875, 
    2.139343, 2.247406, 2.333832, 2.409058, 2.445496, 2.430389, 2.401611, 
    2.343506, 2.30899, 2.300201, 2.285156, 2.203125, 2.055939, 1.952423, 
    2.062225, 2.449219, 3.431641, 3.790894, 3.637054,
  3.325562, 3.354187, 3.215485, 3.172028, 2.957367, 2.428528, 2.843414, 
    2.720428, 2.619781, 3.085449, 3.235382, 3.125336, 3.398254, 3.129211, 
    2.876984, 3.01358, 3.209869, 3.609467, 4.083557, 4.761597, 5.403534, 
    7.971039, 5.672256, 5.329529, 4.928406, 5.47229, 4.614838, 2.798981, 
    2.331726, 4.358612, 4.316376, 4.247284, 4.341156, 1.476501, 1.70816, 
    2.18042, 2.199402, 2.238281, 2.240234, 2.198425, 2.140839, 2.055817, 
    1.989441, 1.938019, 1.882904, 1.818024, 1.742828, 1.707672, 1.678131, 
    1.609009, 1.571686, 1.562927, 1.599487, 1.70285, 1.837708, 1.957611, 
    2.024597, 2.030548, 2.030975, 2.082336, 2.049225, 1.969147, 1.955139, 
    1.969788, 2.081177, 3.320313, 3.733551, 2.876465, 2.833893, 3.216766, 
    2.979553, 2.549713, 2.261475, 2.042175, 1.87204, 1.835236, 1.950256, 
    2.042511, 2.072266, 2.010406, 1.983795, 1.990082, 2.045044, 2.074432, 
    2.062836, 2.057343, 2.076691, 2.151611, 2.278687, 2.314514, 2.159058, 
    2.000458, 2.056, 2.440094, 3.497192, 3.509979,
  3.316956, 3.158813, 2.89386, 2.707031, 2.486511, 2.287689, 2.117096, 
    2.111267, 2.434052, 2.630096, 2.537903, 3.255707, 3.282318, 3.153595, 
    3.045929, 2.812286, 2.856812, 2.874451, 5.873169, 5.963745, 5.948502, 
    5.209732, 4.963974, 4.440536, 4.352402, 4.245667, 3.979248, 2.811066, 
    3.806793, 3.488281, 2.265564, 2.575134, 2.93631, 1.725952, 2.659546, 
    2.477814, 2.874329, 2.852814, 2.336121, 2.284576, 2.22995, 2.189575, 
    2.156891, 2.098267, 2.043427, 1.996674, 1.931183, 1.897461, 1.886414, 
    1.841034, 1.774536, 1.70105, 1.660675, 1.691742, 1.768829, 1.921814, 
    2.037567, 2.029419, 2.015747, 2.026154, 1.995117, 1.917206, 1.907867, 
    2.036987, 2.780304, 2.994843, 2.522247, 1.904388, 1.806946, 2.868866, 
    2.830566, 2.765869, 2.697693, 2.646515, 2.951019, 2.714813, 2.256714, 
    2.099823, 2.084442, 2.142181, 2.146423, 1.970703, 1.729095, 1.650757, 
    1.650055, 1.625977, 1.609314, 1.642303, 1.836151, 2.198761, 2.284058, 
    2.078186, 1.913605, 2.03775, 2.33255, 2.847076,
  2.465149, 2.466522, 2.489838, 2.41861, 2.406372, 2.294922, 2.422119, 
    2.18161, 2.257721, 2.524109, 3.462921, 4.977539, 3.962067, 3.09845, 
    2.282776, 2.802826, 2.48291, 2.310455, 2.790771, 4.783966, 4.02037, 
    4.321045, 4.161224, 3.775482, 4.108276, 4.218323, 4.121368, 3.928345, 
    4.293945, 4.226013, 3.789276, 3.954468, 4.075531, 3.785309, 4.044098, 
    2.704407, 2.486359, 3.357208, 2.486877, 2.532349, 2.548553, 2.520111, 
    2.521423, 2.4711, 2.3638, 2.273621, 2.168304, 2.047729, 1.968628, 
    1.931885, 1.922333, 1.851501, 1.809814, 1.866669, 1.96701, 2.04187, 
    2.065094, 2.066223, 2.094727, 2.099915, 2.094666, 1.985046, 1.936462, 
    2.324432, 3.520538, 4.696381, 5.036346, 4.021423, 2.31723, 1.572418, 
    2.392883, 2.600403, 2.858765, 3.184875, 3.664886, 4.050812, 3.982391, 
    3.227936, 2.975922, 2.885223, 2.695953, 2.376801, 1.855133, 1.159119, 
    0.8688965, 1.006378, 0.9897156, 0.8126831, 0.8367004, 1.350311, 1.904541, 
    1.964966, 1.880402, 1.92218, 2.014923, 2.318787,
  2.717743, 2.451782, 2.552429, 3.063965, 2.623444, 3.224701, 3.865021, 
    3.211517, 2.896515, 2.750397, 3.00354, 3.735107, 4.105743, 2.386108, 
    2.474304, 2.487213, 2.468262, 1.568787, 1.866425, 3.511536, 3.820618, 
    4.305481, 4.467468, 4.505432, 4.55249, 4.60907, 4.506256, 4.163177, 
    4.102112, 4.03891, 3.952942, 4.036255, 3.967804, 3.49057, 3.180222, 
    3.122498, 2.730682, 2.610779, 3.334198, 3.38205, 3.75238, 3.25351, 
    2.482727, 2.21936, 2.088104, 2.055176, 2.041687, 2.071716, 2.094299, 
    2.036499, 1.958099, 1.919708, 1.92984, 2.007233, 2.137024, 2.229523, 
    2.231934, 2.211578, 2.184387, 2.097961, 2.057159, 1.965607, 1.949554, 
    2.40799, 3.987183, 3.86377, 3.283264, 2.85202, 2.287781, 2.168701, 
    2.685577, 3.623199, 4.407379, 4.814392, 4.897156, 5.062988, 5.512329, 
    5.337128, 4.746002, 4.443848, 3.401947, 2.289551, 1.954803, 1.495087, 
    1.116272, 0.6211548, 0.4198608, 0.4104919, 0.4300842, 0.9015503, 
    1.334106, 1.678925, 1.830872, 1.862457, 1.958374, 2.654327,
  3.027374, 3.124329, 4.670197, 4.79715, 3.861877, 4.311676, 4.796692, 
    4.310486, 3.83725, 3.407562, 2.852692, 3.288574, 3.239075, 2.618835, 
    2.296692, 3.453125, 3.66745, 3.677673, 3.673981, 3.554626, 3.63089, 
    3.653015, 3.607635, 3.642685, 3.944321, 3.692245, 3.624527, 3.651413, 
    3.766251, 3.472275, 3.142456, 3.437927, 3.61496, 3.341019, 3.27948, 
    3.399536, 3.305389, 2.6828, 2.993866, 2.829468, 2.807068, 2.492889, 
    2.411346, 2.225281, 2.078247, 1.999664, 1.962799, 1.982819, 2.015442, 
    1.981354, 2.011749, 2.063751, 2.109619, 2.135895, 2.183319, 2.238403, 
    2.245087, 2.186493, 2.200806, 2.235138, 2.237671, 2.08609, 2.052643, 
    2.42569, 3.767059, 3.192261, 3.02063, 3.063293, 2.944946, 3.097931, 
    3.615387, 3.943909, 5.073242, 8.091339, 5.896576, 5.34494, 5.098663, 
    5.425934, 5.865265, 6.337067, 3.905365, 2.997375, 2.410706, 1.864227, 
    1.463959, 1.225037, 0.6382446, 0.08972168, -0.2008362, 0.1266785, 
    0.671936, 1.199799, 1.622009, 1.762177, 2.030853, 2.541382,
  2.618652, 2.850433, 4.15802, 4.884338, 4.751831, 4.609833, 4.453552, 
    4.197144, 4.1297, 4.27533, 4.518036, 4.476257, 4.086914, 3.577759, 
    3.377747, 3.528931, 3.660828, 3.495728, 3.20575, 3.226959, 3.628204, 
    3.703156, 3.393433, 3.351364, 3.293732, 3.23587, 3.341064, 3.424728, 
    3.370163, 3.268661, 3.542038, 3.578491, 3.309677, 3.148224, 3.530838, 
    3.511322, 3.037094, 4.025436, 7.83313, 10.24014, 5.596832, 3.760895, 
    2.881104, 2.531921, 2.458618, 2.306152, 2.338196, 2.360657, 2.344879, 
    2.329987, 2.317352, 2.357056, 2.40036, 2.406403, 2.388824, 2.438629, 
    2.444366, 2.369629, 2.379456, 2.348816, 2.307526, 2.263519, 2.542358, 
    2.860321, 3.133789, 3.014038, 3.795654, 4.415771, 4.575348, 4.712067, 
    4.289337, 4.333923, 4.404083, 5.071793, 5.584427, 5.988861, 6.500046, 
    6.425613, 5.958115, 5.511841, 5.339874, 6.431976, 5.139221, 2.762146, 
    1.886169, 1.278748, 0.4602356, -0.5426941, -1.069885, -0.8245239, 
    -0.04067993, 0.8285217, 1.435883, 1.640411, 1.778961, 1.93811,
  2.315216, 2.082977, 2.892365, 3.56427, 3.893188, 4.025146, 3.811951, 
    3.92984, 3.858887, 4.048431, 4.034332, 3.730164, 3.680176, 3.847961, 
    4.098083, 3.888916, 3.618103, 3.532379, 3.651886, 3.797607, 3.72435, 
    4.043381, 3.816635, 3.775269, 3.765472, 3.519501, 3.55896, 3.635193, 
    3.446915, 3.411575, 3.951874, 3.629089, 3.37355, 3.411972, 3.802582, 
    3.508316, 2.978241, 4.338715, 7.302002, 12.22012, 8.950348, 6.255676, 
    4.490448, 2.921906, 2.940979, 2.473663, 2.295471, 2.250031, 2.297089, 
    2.339264, 2.512512, 2.841522, 3.086884, 3.098755, 2.881287, 2.986694, 
    2.806091, 2.527039, 2.452637, 2.463654, 2.3591, 3.711731, 3.651581, 
    3.72406, 3.549286, 3.592987, 4.507629, 4.823456, 5.228317, 5.153564, 
    5.219208, 4.884216, 5.227509, 6.008453, 6.987732, 11.26593, 8.487152, 
    7.412552, 5.986755, 6.095551, 7.903824, 12.02194, 8.662323, 2.985779, 
    1.481934, 1.323608, 0.8424072, -0.1554565, -0.8538513, -0.854187, 
    -0.1951599, 0.6895142, 1.333252, 1.575226, 2.039795, 2.237274,
  1.428741, 1.540527, 1.54306, 3.536346, 3.741608, 2.793335, 3.351257, 
    2.766663, 2.704376, 3.23584, 3.941254, 3.913055, 3.333954, 3.414551, 
    3.552582, 3.60997, 3.295853, 3.414017, 3.784851, 4.250015, 4.407104, 
    4.411011, 4.621811, 4.593552, 4.683777, 4.558044, 4.186829, 3.683777, 
    3.50441, 3.485077, 3.383057, 3.452972, 3.433838, 3.499847, 3.436707, 
    3.700623, 3.907211, 5.166702, 7.308762, 9.827271, 9.260925, 8.502106, 
    6.194183, 5.272186, 5.668762, 3.403534, 3.733948, 4.670563, 4.629272, 
    5.195404, 5.794434, 6.291046, 5.588196, 5.131805, 5.603119, 3.323334, 
    3.097626, 2.736511, 2.696594, 2.771454, 4.876617, 4.729309, 4.301575, 
    4.366699, 4.778198, 5.476105, 5.635666, 5.163132, 4.870758, 5.147125, 
    5.910278, 6.48761, 7.870819, 8.915344, 10.29907, 11.11137, 8.546005, 
    7.329483, 6.674728, 7.499725, 9.946976, 13.26796, 8.164368, 2.598267, 
    1.145386, 1.510254, 1.675446, 1.175446, 0.5917053, 0.4606323, 0.702179, 
    1.026917, 1.314636, 1.518066, 1.575012, 1.941711,
  0.9687195, 1.167999, 2.450592, 2.887573, 3.646179, 6.123962, 3.782562, 
    3.309143, 2.776581, 2.694244, 3.039337, 3.293564, 3.270493, 3.294266, 
    3.598633, 3.905075, 4.083405, 4.144333, 4.102615, 4.258987, 4.268875, 
    5.032211, 5.385208, 5.481949, 5.479858, 4.703033, 4.739365, 4.453308, 
    4.052124, 3.743927, 3.408447, 3.409561, 3.609238, 3.886826, 4.342834, 
    4.605087, 4.711731, 4.905228, 5.255707, 5.736176, 6.030716, 5.869385, 
    5.76619, 5.460541, 5.54393, 6.763062, 9.000702, 16.1871, 15.42993, 
    14.28252, 13.6792, 12.65009, 8.08696, 6.933777, 6.307831, 6.28598, 
    6.482605, 5.95903, 5.726669, 5.696136, 5.343353, 4.983063, 4.827255, 
    5.079483, 5.657394, 6.158844, 6.019913, 5.681885, 5.758377, 6.141464, 
    6.73085, 7.114838, 7.785843, 8.435532, 8.801819, 8.962677, 8.095047, 
    7.554474, 6.832855, 7.606049, 8.230057, 8.398621, 5.078644, 2.859863, 
    2.526062, 1.810303, 1.23468, 1.205109, 1.267548, 1.405182, 1.381348, 
    1.046692, 0.3726196, 0.1701965, 0.6714478, 0.8805542,
  0.262207, 0.4883118, 0.5400696, 2.577179, 3.389923, 4.037994, 5.87912, 
    3.696091, 3.450333, 3.363678, 3.490417, 3.782501, 3.77005, 3.9375, 
    4.128525, 4.290115, 4.785736, 5.098557, 5.30722, 5.503433, 5.379745, 
    5.574326, 5.584351, 5.592438, 5.821533, 5.247772, 5.095627, 4.966125, 
    4.813461, 4.579086, 4.586761, 4.252747, 4.306473, 4.783218, 4.855545, 
    5.261612, 5.866882, 5.716995, 6.070068, 6.009705, 5.938812, 6.3685, 
    6.383972, 5.969589, 5.730774, 5.586777, 5.681763, 5.750381, 5.923752, 
    6.102585, 6.344193, 7.638855, 6.489365, 6.300171, 6.035934, 6.164108, 
    6.30162, 6.484222, 6.312744, 6.147186, 6.202133, 6.315277, 6.157654, 
    6.490219, 6.338394, 6.162994, 6.194778, 6.061172, 6.194199, 6.465347, 
    6.481766, 6.611771, 7.126541, 7.626999, 7.991638, 7.894241, 7.858383, 
    7.406113, 7.071274, 7.099136, 6.542816, 5.807724, 4.413254, 3.454208, 
    2.532928, 2.491898, 2.21138, 1.264404, 1.049316, 2.080231, 3.920258, 
    4.211151, 2.729462, 0.9982605, 0.118866, 0.06085205,
  0.5985413, 0.2869568, 0.177887, 0.0652771, -0.5629883, 1.311279, 1.706635, 
    2.250244, 3.29686, 4.618698, 6.143753, 9.472855, 9.247803, 7.99733, 
    5.733597, 5.455704, 5.11412, 5.252914, 5.647766, 5.954147, 6.171661, 
    6.354797, 6.490662, 6.646988, 6.541321, 6.717636, 6.247314, 5.872086, 
    5.437378, 5.409912, 5.582764, 5.51741, 5.281845, 4.871033, 5.245514, 
    5.358475, 5.582962, 5.914673, 6.127228, 6.295456, 6.452744, 6.412521, 
    6.431198, 6.437836, 6.917557, 7.085785, 7.524719, 7.782806, 7.966583, 
    7.76503, 7.939774, 8.136124, 8.271606, 7.045242, 6.638535, 6.625565, 
    6.880249, 7.360275, 7.192169, 7.58345, 7.629211, 7.177521, 7.337418, 
    7.160797, 7.106506, 6.779602, 6.701752, 6.583908, 6.660339, 6.437744, 
    6.770096, 6.861923, 7.20932, 7.033783, 7.637573, 7.654999, 7.822998, 
    7.711014, 7.409836, 6.62088, 5.805328, 4.335587, 4.162231, 3.394699, 
    3.150436, 3.347336, 3.134399, 2.742752, 3.20253, 4.381683, 6.257736, 
    7.87178, 10.01796, 8.712799, 3.451904, 1.521515,
  3.107361, 1.761902, 1.059235, 0.7766113, 0.4829102, 0.7835388, 1.866364, 
    3.602417, 6.49292, 9.332428, 11.71417, 13.32486, 12.88304, 10.14809, 
    8.689316, 7.740036, 6.827194, 6.899338, 6.901749, 6.876678, 6.747711, 
    6.845032, 7.146271, 7.259689, 7.177979, 6.888626, 6.656265, 6.275787, 
    5.982697, 6.186142, 5.869476, 6.008926, 5.968307, 5.931854, 5.895386, 
    5.3797, 5.741669, 6.004196, 6.72937, 6.646378, 6.128998, 6.346176, 
    6.328598, 6.441025, 6.523071, 6.60083, 6.641586, 6.864685, 7.131363, 
    7.272049, 7.302856, 7.269958, 7.16066, 7.053757, 7.09198, 7.219254, 
    7.445175, 7.58287, 7.588333, 7.595093, 7.728821, 7.831223, 7.73703, 
    7.771271, 7.577972, 7.228317, 7.04071, 7.122406, 7.294861, 7.027649, 
    7.811737, 8.464081, 7.417953, 8.383804, 8.368637, 7.844604, 7.389664, 
    6.583374, 6.241196, 6.123291, 5.230911, 4.845306, 3.591919, 2.419708, 
    1.528076, 2.014404, 2.408676, 2.616486, 2.58989, 3.145691, 4.415146, 
    5.703049, 6.727524, 7.441864, 7.909637, 7.433472,
  7.712067, 6.253784, 3.44754, 3.080688, 5.205475, 8.917786, 10.97862, 
    11.00084, 10.95915, 10.59348, 10.04907, 9.4888, 9.050125, 8.449265, 
    7.966904, 7.983185, 7.947052, 8.008636, 8.057266, 8.056747, 7.875763, 
    7.71405, 7.668335, 7.693008, 7.549194, 8.043137, 7.830154, 7.330292, 
    7.096954, 6.966095, 6.635956, 6.038742, 5.985626, 6.088104, 6.155869, 
    6.346313, 6.628922, 6.73497, 6.836868, 6.907318, 7.011597, 7.112259, 
    7.16069, 7.22229, 7.263885, 7.308014, 7.335785, 7.453827, 7.571533, 
    7.699005, 7.79126, 7.823547, 7.861374, 7.896866, 7.872635, 7.769638, 
    7.591187, 7.374969, 7.159683, 7.093155, 7.106689, 7.285263, 7.471207, 
    7.794067, 8.00174, 7.577682, 7.635239, 7.654449, 7.684448, 7.821365, 
    7.940369, 8.213684, 8.267395, 8.133682, 7.790192, 6.902878, 7.133804, 
    6.320297, 6.918381, 5.778931, 4.782639, 4.126511, 3.456848, 2.640381, 
    2.190643, 2.479828, 2.873459, 3.324036, 3.65387, 4.244751, 5.083588, 
    6.104477, 6.96463, 7.488403, 7.724731, 7.766312,
  7.756165, 7.420227, 7.152863, 7.168091, 7.481369, 7.482742, 7.502655, 
    7.844894, 7.95343, 7.990936, 7.951019, 7.906097, 7.917816, 7.954727, 
    8.046799, 8.118225, 8.191711, 8.264511, 8.350769, 8.371078, 8.272186, 
    8.060211, 7.79158, 7.611252, 7.493607, 8.06636, 7.961533, 7.042175, 
    6.864334, 6.81395, 6.721436, 6.8508, 6.907776, 6.881851, 6.924179, 
    7.004257, 7.024246, 7.031799, 7.041092, 7.014206, 6.956787, 6.940445, 
    6.945923, 7.012253, 7.174423, 7.345596, 7.482056, 7.667313, 7.868591, 
    7.953506, 7.921997, 7.820175, 7.693008, 7.497604, 7.31929, 7.169678, 
    7.046432, 6.980225, 6.98674, 7.071243, 7.199875, 7.263168, 7.320786, 
    7.417007, 7.522339, 7.69104, 7.81395, 7.900925, 7.974228, 8.093506, 
    8.324753, 7.696304, 7.574753, 7.60112, 7.366226, 7.002228, 6.557632, 
    6.073837, 5.501907, 4.911926, 4.442734, 4.031784, 3.800156, 3.69455, 
    3.794357, 4.050476, 4.291031, 4.625534, 5.139084, 5.934906, 6.709259, 
    7.231003, 7.73793, 7.789688, 7.925186, 7.916443,
  8.238968, 8.116135, 8.058701, 7.998108, 7.83963, 7.760925, 7.75441, 7.6716, 
    7.614182, 7.626862, 7.663589, 7.703171, 7.748947, 7.825882, 7.848038, 
    7.890411, 7.888794, 7.868073, 7.828232, 7.75795, 7.644547, 7.569229, 
    7.435822, 7.316422, 7.239594, 7.113815, 7.002426, 6.975342, 6.972092, 
    6.979904, 7.044022, 7.203598, 7.356659, 7.490173, 7.588684, 7.630096, 
    7.66095, 7.691818, 7.703537, 7.702103, 7.676773, 7.626648, 7.586548, 
    7.501648, 7.442261, 7.474823, 7.515121, 7.514404, 7.522736, 7.54657, 
    7.565643, 7.577621, 7.575073, 7.575211, 7.563156, 7.565186, 7.609711, 
    7.682648, 7.725937, 7.789078, 7.900925, 7.966034, 8.006592, 8.025604, 
    8.033737, 8.035965, 7.986343, 7.91832, 7.874557, 7.824234, 7.772812, 
    7.80484, 7.961731, 8.039276, 8.084259, 8.082169, 7.965836, 7.916031, 
    8.026718, 8.179504, 8.235504, 8.161285, 8.076187, 7.914139, 7.936478, 
    8.137848, 8.237396, 8.351456, 8.487915, 8.446823, 8.517532, 8.591156, 
    8.490646, 8.455688, 8.415833, 8.325165,
  8.326584, 8.292206, 8.230682, 8.209, 8.173386, 8.121765, 8.052032, 
    7.980606, 7.934921, 7.876785, 7.823135, 7.777496, 7.746231, 7.693375, 
    7.623444, 7.563293, 7.494019, 7.456207, 7.416031, 7.367722, 7.335953, 
    7.306854, 7.286865, 7.2715, 7.247665, 7.243622, 7.274628, 7.287384, 
    7.28479, 7.339279, 7.34169, 7.37085, 7.393829, 7.488098, 7.54332, 
    7.557495, 7.585175, 7.651306, 7.703339, 7.753403, 7.795853, 7.820068, 
    7.84169, 7.8741, 7.92482, 7.964203, 7.990509, 8.013565, 8.039215, 
    8.057114, 8.062378, 8.07338, 8.097488, 8.125015, 8.091949, 8.056854, 
    8.041885, 8.022995, 8.003723, 8.007187, 8.016098, 8.001312, 7.965118, 
    7.968506, 7.969559, 7.981003, 8.003784, 8.037323, 8.042725, 8.025482, 
    8.033356, 8.042267, 8.042587, 8.070068, 8.106781, 8.146179, 8.168564, 
    8.191681, 8.228989, 8.266418, 8.312912, 8.333801, 8.349945, 8.3741, 
    8.39064, 8.41629, 8.422546, 8.421371, 8.428665, 8.427231, 8.455688, 
    8.447159, 8.442017, 8.425934, 8.384399, 8.360306,
  2.138275, 2.050201, 1.975189, 1.911392, 1.857483, 1.806305, 1.762131, 
    1.723465, 1.693436, 1.66922, 1.653793, 1.649948, 1.651382, 1.653976, 
    1.656525, 1.660751, 1.665451, 1.67157, 1.676514, 1.685165, 1.695602, 
    1.705032, 1.715378, 1.727692, 1.73941, 1.749695, 1.765381, 1.783615, 
    1.806717, 1.835434, 1.872284, 1.918365, 1.970718, 2.030289, 2.087906, 
    2.142914, 2.198883, 2.252213, 2.308975, 2.36673, 2.424026, 2.478577, 
    2.532089, 2.5858, 2.632172, 2.67598, 2.708664, 2.770905, 2.819138, 
    2.886002, 2.908066, 2.951691, 3.051956, 3.042786, 2.989777, 3.072006, 
    3.062637, 3.105469, 3.153915, 3.125198, 3.175583, 3.119858, 3.11412, 
    3.10788, 3.091537, 3.072144, 3.027008, 2.986786, 2.937042, 2.89122, 
    2.83255, 2.784836, 2.737244, 2.770447, 2.708405, 2.658478, 2.673706, 
    2.658386, 2.648697, 2.667175, 2.681717, 2.700455, 2.722916, 2.732239, 
    2.740631, 2.742905, 2.737183, 2.716202, 2.682098, 2.63887, 2.587112, 
    2.530731, 2.470764, 2.397141, 2.316788, 2.228714,
  1.364975, 1.217316, 1.096939, 1.004166, 0.9510651, 0.9558105, 1.034714, 
    1.185028, 1.380814, 1.580109, 1.749832, 1.855026, 1.884583, 1.826981, 
    1.748398, 1.669937, 1.579575, 1.471497, 1.356201, 1.250534, 1.177612, 
    1.133682, 1.13179, 1.1577, 1.210556, 1.288757, 1.380234, 1.477493, 
    1.568192, 1.649887, 1.724106, 1.792267, 1.865128, 1.938416, 2.019669, 
    2.123367, 2.243881, 2.382294, 2.538406, 2.707474, 2.876114, 3.079895, 
    3.256409, 3.370331, 3.485962, 3.627228, 3.716171, 3.817535, 3.890564, 
    3.920013, 3.929245, 3.867264, 3.818115, 3.753281, 3.707825, 3.531326, 
    3.411926, 3.314606, 3.244873, 3.208603, 3.148911, 3.109573, 3.072083, 
    3.070587, 3.036804, 3.00145, 2.917252, 2.866852, 2.720886, 2.609299, 
    2.596039, 2.614777, 2.601639, 2.58046, 2.60585, 2.595108, 2.590378, 
    2.604706, 2.640381, 2.66655, 2.681274, 2.697678, 2.743896, 2.688492, 
    2.653717, 2.611542, 2.555161, 2.536743, 2.511734, 2.453979, 2.338669, 
    2.188217, 2.031113, 1.853134, 1.678635, 1.516724,
  1.028198, 0.7617798, 0.5706329, 0.4753113, 0.5511322, 0.7867889, 1.129196, 
    1.483795, 1.73732, 1.838562, 1.898071, 2.006454, 2.165451, 2.332245, 
    2.473511, 2.533356, 2.550079, 2.537521, 2.528656, 2.514664, 2.545197, 
    2.550156, 2.442078, 2.157303, 1.797928, 1.701523, 1.819946, 1.972412, 
    2.035751, 1.953857, 1.822281, 1.704773, 1.596436, 1.573654, 1.613739, 
    1.731903, 1.909058, 2.087952, 2.277481, 2.482803, 2.695389, 2.953598, 
    3.231339, 3.550278, 3.924301, 4.141754, 4.248123, 4.17424, 4.008286, 
    3.844742, 3.680557, 3.449158, 3.201508, 2.970459, 2.846375, 2.789474, 
    2.704498, 2.548981, 2.461273, 2.416946, 2.367462, 2.377289, 2.470795, 
    2.568436, 2.65712, 2.649887, 2.462524, 2.286148, 2.215057, 2.215637, 
    2.271301, 2.34111, 2.386276, 2.401443, 2.374313, 2.337463, 2.397736, 
    2.373581, 2.399689, 2.443893, 2.498978, 2.57872, 2.693253, 2.712708, 
    2.555679, 2.366943, 2.179901, 1.953201, 1.869034, 1.883102, 1.832901, 
    1.862, 1.823898, 1.693619, 1.525467, 1.279694,
  1.518875, 1.56308, 1.575897, 1.681458, 1.795059, 1.956009, 2.093643, 
    2.025543, 1.863358, 1.623596, 1.467712, 1.556076, 1.810623, 2.069809, 
    2.298035, 2.543625, 2.748505, 2.934769, 3.158142, 3.241928, 2.87175, 
    2.348099, 1.929947, 1.612427, 1.385696, 1.29657, 1.356918, 1.479385, 
    1.482239, 1.43869, 1.465057, 1.510437, 1.489151, 1.44162, 1.443115, 
    1.451508, 1.48111, 1.576431, 1.705154, 1.81015, 1.871811, 2.003723, 
    2.252686, 2.681915, 3.20932, 3.561478, 4.088959, 3.993668, 3.761459, 
    3.546448, 3.235245, 2.95842, 2.805359, 2.695343, 2.641937, 2.612457, 
    2.687073, 2.144958, 2.245667, 2.309402, 2.36525, 2.433273, 2.464935, 
    2.503067, 2.559387, 2.579437, 2.663422, 2.691345, 2.610947, 2.583557, 
    2.596497, 2.62619, 2.675858, 2.74057, 2.854568, 3.025406, 3.121307, 
    3.229889, 3.247147, 3.292465, 3.229904, 3.322617, 3.262192, 3.306305, 
    3.361893, 3.400314, 3.383377, 3.424332, 3.673706, 1.992401, 1.665512, 
    1.514404, 1.468826, 1.420258, 1.402283, 1.460602,
  1.057053, 0.9035339, 0.8161011, 0.8568573, 0.9225464, 1.037918, 1.162659, 
    1.300415, 1.355484, 1.4711, 1.648453, 1.786392, 1.774994, 1.719208, 
    1.842834, 1.970062, 2.035019, 2.117447, 1.984894, 1.890045, 2.336807, 
    2.035629, 1.601196, 1.384583, 1.422974, 1.512558, 1.542572, 1.654556, 
    1.874817, 1.962631, 2.007874, 2.042709, 2.038284, 2.10553, 2.168304, 
    2.242767, 2.179031, 2.038223, 1.899612, 1.851166, 1.68959, 1.663818, 
    1.774628, 1.965256, 2.209518, 2.429001, 3.312637, 2.990723, 2.367249, 
    1.97345, 1.668121, 1.453796, 1.391418, 1.514862, 1.667938, 1.953339, 
    2.361237, 2.724701, 2.932129, 3.179962, 3.392273, 3.575867, 3.555878, 
    3.332611, 3.114777, 2.936005, 2.884979, 3.130402, 3.488678, 3.76532, 
    4.581635, 4.898712, 4.950745, 4.600586, 4.108765, 3.810364, 4.013351, 
    4.024368, 3.928207, 3.651306, 3.32489, 3.339584, 3.583221, 3.874619, 
    4.241882, 4.577118, 4.799866, 4.947815, 5.037323, 5.041504, 4.813751, 
    2.708771, 2.212677, 1.840759, 1.497223, 1.221436,
  5.101318, 4.256866, 2.856461, 2.131912, 1.605545, 1.263763, 1.145584, 
    1.315826, 1.310623, 1.447617, 1.588623, 1.693436, 1.780151, 1.866089, 
    1.869751, 1.821365, 1.511734, 1.369675, 1.34227, 1.427673, 1.600021, 
    1.687393, 1.469482, 1.189545, 1.083801, 1.024506, 0.9961243, 1.136215, 
    1.274887, 1.395584, 1.259201, 1.120331, 1.175674, 1.328003, 1.445724, 
    1.48732, 1.513046, 1.541626, 1.534729, 1.638367, 1.756851, 1.750992, 
    1.682175, 1.596176, 2.06369, 1.140198, 0.9090576, 0.2692871, 0.1218262, 
    0.1545715, 0.1744385, 0.1072388, -0.01196289, -0.08755493, -0.06704712, 
    0.04879761, 0.2293091, 0.4432678, 0.6386108, 0.8429871, 1.128845, 
    1.348206, 1.507782, 1.52887, 1.483917, 1.413269, 1.467499, 1.499725, 
    1.598724, 1.972076, 2.604156, 3.558868, 3.297089, 2.665253, 2.119019, 
    1.934265, 2.010559, 2.085052, 3.299316, 3.694214, 4.187164, 4.342865, 
    4.568634, 5.029266, 5.44696, 5.846893, 6.117676, 6.282898, 6.3974, 
    6.717712, 6.871033, 7.133362, 7.539154, 7.418121, 7.049377, 6.172729,
  5.341095, 5.68576, 6.036835, 5.97525, 5.746613, 5.333496, 5.082916, 
    4.891815, 4.613434, 4.399353, 4.329315, 4.506653, 4.398376, 4.261169, 
    4.068115, 3.908722, 3.824493, 3.570343, 3.46994, 3.504059, 3.427307, 
    3.385773, 3.071045, 2.733063, 2.358612, 1.756195, 1.264069, 0.7737732, 
    0.4527588, 0.386261, 0.3948669, 0.3380127, 0.521759, 1.859528, 2.191742, 
    2.449707, 3.610809, 1.463226, 1.120453, 1.053986, 1.273529, 1.177765, 
    1.020935, 0.9191589, 0.6546936, 0.2887573, -0.08514404, -0.3208313, 
    -0.3746033, -0.3074951, -0.1885376, -0.1210938, -0.1366577, -0.1826782, 
    -0.2102051, -0.1789551, -0.07369995, 0.04992676, 0.1627502, 0.2979431, 
    0.4865417, 0.6694031, 0.8058167, 0.9300842, 1.068451, 1.213806, 1.33725, 
    1.406982, 1.463867, 1.526093, 1.624023, 1.736633, 1.750671, 1.687164, 
    1.596832, 1.485687, 1.360809, 1.338165, 1.745239, 2.834198, 4.057495, 
    3.690308, 3.284576, 2.825592, 2.675049, 2.833923, 3.238281, 3.741211, 
    3.932556, 4.048645, 4.326691, 4.618195, 4.849701, 4.875641, 4.928131, 
    5.063538,
  1.803711, 1.851379, 1.839142, 1.754608, 1.641846, 1.566772, 1.571686, 
    1.625824, 1.612244, 1.558136, 1.541412, 1.613678, 1.687622, 1.698578, 
    1.717255, 1.764282, 1.84024, 1.847443, 1.747864, 1.573334, 1.422058, 
    1.29361, 1.186462, 1.111267, 1.074432, 1.009491, 0.8683472, 0.707428, 
    0.5790405, 0.518158, 0.4967651, 0.5098267, 0.5606079, 0.6554871, 
    0.8331909, 0.9874878, 1.084961, 1.058594, 0.9958496, 1.041595, 1.154419, 
    1.201843, 1.160614, 1.076569, 0.8832703, 0.5575562, 0.116333, -0.2349548, 
    -0.3742676, -0.419281, -0.4680786, -0.4885254, -0.4552612, -0.3772583, 
    -0.2705078, -0.1054077, 0.05859375, 0.1777344, 0.2363281, 0.3268127, 
    0.459259, 0.6211548, 0.730011, 0.8327942, 1.055908, 1.305603, 1.510864, 
    1.622681, 1.671753, 1.72876, 1.847717, 1.980469, 2.040771, 2.058716, 
    2.049408, 1.957733, 1.791016, 1.6138, 1.531189, 1.654755, 1.948364, 
    1.971222, 1.632111, 1.25946, 1.283447, 1.440369, 1.637909, 1.800079, 
    1.870453, 1.887573, 1.865143, 1.842316, 1.845947, 1.815521, 1.775269, 
    1.767456,
  1.472992, 1.474274, 1.407135, 1.283142, 1.152008, 1.068726, 1.051849, 
    1.06958, 1.094879, 1.109772, 1.158539, 1.269135, 1.357666, 1.392914, 
    1.417633, 1.463928, 1.530457, 1.569183, 1.528107, 1.426117, 1.332489, 
    1.212494, 1.054871, 1.004425, 1.077148, 1.137177, 1.149292, 1.121185, 
    1.055084, 0.9579468, 0.8087769, 0.6594849, 0.5491333, 0.4667358, 
    0.4367371, 0.4902954, 0.5846863, 0.717041, 0.9068909, 1.081573, 1.192139, 
    1.282349, 1.382294, 1.311401, 1.120056, 0.9771423, 0.8140564, 0.5292358, 
    0.1312256, -0.2092896, -0.3370667, -0.3686829, -0.348175, -0.2983093, 
    -0.2589111, -0.1607361, 0.04275513, 0.2431641, 0.2889404, 0.2849731, 
    0.4560547, 0.6708374, 0.7927856, 0.9051819, 1.177673, 1.47702, 1.637054, 
    1.68866, 1.728394, 1.803894, 1.907562, 1.998901, 2.049347, 2.067657, 
    2.009583, 1.85614, 1.652283, 1.569733, 1.566864, 1.632568, 1.747223, 
    1.832031, 1.720001, 1.391022, 1.213623, 1.193481, 1.300262, 1.393829, 
    1.483063, 1.515106, 1.530151, 1.515289, 1.49649, 1.515228, 1.509308, 
    1.479614,
  1.475128, 1.574677, 1.644775, 1.641602, 1.605469, 1.575897, 1.58313, 
    1.561768, 1.534882, 1.533936, 1.562561, 1.617065, 1.647919, 1.681061, 
    1.800934, 1.940033, 2.118622, 2.264435, 2.207214, 1.934967, 1.756195, 
    1.647125, 1.458679, 1.299225, 1.282104, 1.360657, 1.449738, 1.487244, 
    1.451172, 1.326172, 1.147797, 1.003052, 0.9182434, 0.8689575, 0.8215637, 
    0.8208923, 0.8839417, 1.003784, 1.142303, 1.213684, 1.274017, 1.369843, 
    1.445648, 1.374695, 1.293823, 1.266937, 1.169983, 0.9350891, 0.5198975, 
    0.1822205, 0.139801, 0.1936035, 0.2010193, 0.1896667, 0.2092896, 
    0.2703857, 0.3633423, 0.4692688, 0.504303, 0.5169983, 0.6787109, 
    0.8625793, 0.9779358, 1.115875, 1.386597, 1.56366, 1.56015, 1.570526, 
    1.639832, 1.735443, 1.781647, 1.81778, 1.871796, 1.848541, 1.709198, 
    1.445709, 1.404236, 1.902405, 1.940247, 1.503052, 1.475922, 1.569885, 
    1.656036, 1.428253, 1.169922, 1.29715, 1.533081, 1.721558, 1.775177, 
    1.738739, 1.743378, 1.752594, 1.714905, 1.636261, 1.543732, 1.466797,
  1.996552, 2.029022, 2.069214, 2.090973, 2.11499, 2.141724, 2.170258, 
    2.174438, 2.141602, 2.129761, 2.205261, 2.297607, 2.335022, 2.3862, 
    2.48761, 2.611603, 2.792603, 2.976837, 2.954285, 2.76239, 2.668335, 
    2.665833, 2.49649, 2.2034, 1.971344, 1.925323, 1.992432, 1.972931, 
    1.851868, 1.699921, 1.541412, 1.42569, 1.385223, 1.316162, 1.200989, 
    1.125275, 1.140869, 1.204773, 1.302948, 1.444061, 1.574677, 1.640686, 
    1.632538, 1.61673, 1.599091, 1.554504, 1.411407, 1.250183, 1.028961, 
    0.8269043, 0.8244324, 0.9100952, 0.9353638, 0.8900452, 0.8556824, 
    0.8465576, 0.854126, 0.8987732, 0.9765625, 1.041473, 1.132996, 1.234131, 
    1.336395, 1.452484, 1.596283, 1.647339, 1.625, 1.629181, 1.697174, 
    1.727753, 1.705261, 1.695435, 1.668732, 1.600525, 1.544189, 1.502716, 
    1.875458, 1.894531, 1.723175, 1.708649, 1.580078, 1.409546, 1.265045, 
    1.084381, 1.192139, 1.540314, 1.822662, 2.015564, 2.096619, 2.088287, 
    2.085785, 2.083405, 2.048218, 2.032501, 2.049408, 2.015045,
  2.136444, 2.118683, 2.201172, 2.288208, 2.351624, 2.427277, 2.552795, 
    2.669861, 2.705414, 2.795319, 2.983398, 3.108826, 3.174927, 3.214325, 
    3.198822, 3.13028, 3.146423, 3.312103, 3.394348, 3.517731, 3.6763, 
    3.575256, 3.153778, 2.704803, 2.44165, 2.333405, 2.291687, 2.200073, 
    2.025635, 1.82962, 1.699005, 1.680786, 1.690979, 1.656189, 1.59198, 
    1.552551, 1.556519, 1.568115, 1.59024, 1.735535, 2.01947, 2.075653, 
    1.973267, 1.984253, 2.144073, 2.335876, 2.076172, 1.843811, 1.657806, 
    1.540436, 1.666016, 1.792572, 1.782776, 1.660492, 1.510895, 1.432678, 
    1.406311, 1.418488, 1.463684, 1.510406, 1.541077, 1.594208, 1.647186, 
    1.670715, 1.695831, 1.734589, 1.775055, 1.787781, 1.802948, 1.796997, 
    1.73996, 1.723297, 1.681366, 1.6315, 1.59375, 1.505676, 1.728516, 
    1.942963, 2.32254, 1.972473, 1.686462, 1.325531, 1.055908, 1.017334, 
    1.384827, 1.839447, 2.094666, 2.178497, 2.24115, 2.264252, 2.240631, 
    2.231842, 2.222992, 2.211792, 2.24472, 2.221161,
  2.328339, 2.252869, 2.306396, 2.432343, 2.593689, 2.96994, 3.393494, 
    3.591492, 3.750702, 3.970123, 4.098694, 3.978577, 3.719513, 3.526031, 
    3.383667, 3.332306, 3.33783, 3.376251, 3.47525, 3.575073, 3.490784, 
    3.114563, 2.611511, 2.278198, 2.177155, 2.203247, 2.223969, 2.134766, 
    2.033447, 2.002869, 2.010223, 2.029968, 2.011383, 1.937897, 1.931061, 
    2.002716, 2.020172, 1.961243, 1.905334, 2.185425, 2.724213, 2.76413, 
    2.54187, 2.488983, 2.588806, 2.736115, 2.930664, 2.596527, 2.49057, 
    2.506104, 2.625763, 2.472961, 2.227142, 2.039703, 1.865814, 1.794586, 
    1.816467, 1.851959, 1.867584, 1.868225, 1.866547, 1.883667, 1.899689, 
    1.896606, 1.885559, 1.906311, 1.972595, 1.960938, 1.926697, 1.929108, 
    1.868011, 1.799622, 1.722809, 1.653107, 1.588989, 1.456451, 1.699738, 
    2.56073, 3.014374, 2.111725, 1.742706, 1.626495, 1.677032, 1.83847, 
    2.029175, 2.269257, 2.414215, 2.395569, 2.367767, 2.355988, 2.357483, 
    2.413727, 2.458649, 2.464783, 2.460419, 2.417725,
  2.202606, 2.171631, 2.242828, 2.448181, 2.788605, 3.19278, 3.424103, 
    3.885498, 3.916321, 3.525909, 2.986847, 2.548584, 2.295105, 2.173248, 
    2.219391, 2.49231, 2.721985, 2.822601, 2.783264, 2.635803, 2.474213, 
    2.305023, 2.137054, 2.080994, 2.079956, 2.146027, 2.195587, 2.194458, 
    2.266266, 2.388336, 2.317261, 2.260498, 2.174927, 2.027588, 2.162903, 
    2.259827, 2.139923, 2.203766, 2.466492, 2.926422, 2.902039, 3.156952, 
    3.262573, 3.001892, 2.875702, 2.959045, 3.070953, 3.192902, 2.679871, 
    2.495361, 2.370178, 2.330414, 2.258789, 2.193451, 2.12558, 2.070435, 
    2.051086, 2.049561, 2.066406, 2.050842, 2.042908, 2.085297, 2.080811, 
    2.090759, 2.090363, 2.110168, 2.153046, 2.121277, 2.067139, 2.007568, 
    1.921295, 1.884583, 1.765106, 1.599854, 1.494476, 1.289978, 1.368835, 
    2.993927, 3.057861, 2.1633, 1.627869, 1.841125, 2.170624, 2.362061, 
    2.31427, 2.318817, 2.39389, 2.413025, 2.449097, 2.468018, 2.480408, 
    2.479828, 2.410858, 2.333405, 2.260895, 2.235077,
  2.0849, 1.957825, 1.972382, 2.071533, 2.206696, 2.371674, 2.541779, 
    2.589722, 2.36972, 2.101624, 1.440613, 1.62265, 1.789063, 1.951996, 
    2.075012, 2.238129, 2.336731, 2.280457, 2.227936, 2.089111, 2.0737, 
    2.133789, 2.135986, 2.185028, 2.117493, 2.119263, 2.157745, 2.198181, 
    2.320251, 2.222534, 1.959503, 1.984955, 1.872131, 1.820313, 1.969574, 
    1.993042, 2.008728, 2.819275, 3.441345, 3.162109, 2.559509, 2.835083, 
    3.503387, 3.28595, 2.993805, 3.002289, 2.865082, 2.601044, 2.254059, 
    1.932098, 1.990814, 2.113403, 2.21759, 2.233643, 2.230408, 2.244904, 
    2.181, 2.108612, 2.133331, 2.137756, 2.166473, 2.220123, 2.20932, 
    2.215607, 2.209961, 2.151886, 2.13559, 2.05957, 1.957489, 1.873566, 
    1.706238, 1.585632, 1.449158, 1.264374, 1.144135, 1.009186, 1.269836, 
    3.236969, 3.454559, 1.902008, 1.580505, 2.03125, 2.248108, 2.33783, 
    2.15802, 2.081909, 2.160614, 2.279419, 2.434113, 2.436127, 2.40976, 
    2.3862, 2.281097, 2.253967, 2.229156, 2.175262,
  1.665741, 1.595123, 1.58075, 1.726318, 1.976563, 3.245636, 3.274994, 
    3.124023, 2.836639, 1.946686, 1.898651, 2.152039, 2.249084, 2.353302, 
    2.375793, 2.428375, 2.538269, 2.500854, 2.438202, 2.351898, 2.376373, 
    2.33667, 2.230988, 2.215546, 2.181, 2.140625, 2.123718, 2.072845, 
    1.951324, 1.740601, 1.86145, 2.651245, 2.327942, 2.263397, 2.680542, 
    3.194397, 3.38562, 3.508667, 3.69165, 3.039185, 2.396362, 2.442902, 
    2.210236, 2.142639, 2.29303, 2.358337, 2.158936, 1.880463, 1.84845, 
    2.036713, 2.184113, 2.3125, 2.375519, 2.318176, 2.257202, 2.173126, 
    2.088226, 2.045319, 2.096344, 2.135223, 2.105591, 2.130341, 2.132996, 
    2.113953, 2.062622, 1.952667, 1.876251, 1.714996, 1.572449, 1.443054, 
    1.280212, 1.157471, 1.053375, 1.004364, 0.8948669, 0.9748535, 1.497589, 
    2.914398, 3.997772, 2.470245, 2.124542, 2.531891, 2.484314, 2.313995, 
    2.174072, 2.164917, 2.300323, 2.38092, 2.429291, 2.370636, 2.334686, 
    2.234772, 2.097473, 2.034363, 1.942535, 1.830139,
  1.431519, 1.458832, 1.6763, 1.901947, 2.302155, 3.320251, 3.779114, 
    3.422394, 2.735748, 1.982758, 1.973236, 2.234894, 2.261353, 2.417053, 
    2.589111, 2.708984, 2.758209, 2.695313, 2.630005, 2.487366, 2.375519, 
    2.247589, 2.090302, 1.965485, 1.894012, 1.819, 1.770569, 1.792267, 
    1.917328, 1.966339, 2.28302, 3.012238, 2.508636, 2.79425, 3.220184, 
    3.717438, 3.767853, 3.685425, 3.277679, 2.830994, 2.59845, 2.110474, 
    1.671417, 1.779297, 2.054962, 2.19635, 2.19635, 2.179932, 2.226044, 
    2.320923, 2.292206, 2.272369, 2.224487, 2.116913, 2.057617, 2.027405, 
    1.986481, 1.974152, 1.925018, 1.920105, 1.851624, 1.827148, 1.790497, 
    1.672394, 1.58728, 1.429077, 1.328857, 1.192963, 1.106506, 1.060364, 
    0.9658203, 0.9912109, 0.9087219, 0.9498901, 0.8777466, 1.252991, 
    1.968903, 2.889374, 4.383148, 2.918274, 2.170898, 2.940948, 2.864624, 
    2.713745, 2.397064, 2.23822, 2.290344, 2.315552, 2.254089, 2.175781, 
    2.092102, 1.965942, 1.892395, 1.755798, 1.611267, 1.470306,
  1.594116, 1.794922, 2.10733, 2.493225, 3.612488, 4.118042, 4.2435, 
    3.911377, 3.049133, 2.853729, 2.120331, 2.256836, 2.245361, 2.405212, 
    2.54306, 2.61087, 2.478455, 2.299164, 2.250153, 2.156342, 2.017456, 
    1.913239, 1.850739, 1.800385, 1.791779, 1.812378, 1.866333, 2.043304, 
    2.215973, 2.240875, 2.447662, 2.936005, 3.292297, 3.644989, 3.69043, 
    3.399872, 3.259766, 3.001343, 2.520172, 2.17218, 2.167419, 1.989777, 
    2.052338, 2.194794, 2.22879, 2.273621, 2.294525, 2.282013, 2.239716, 
    2.205383, 2.162689, 2.141937, 2.140625, 2.084076, 2.024536, 1.995483, 
    1.944916, 1.912048, 1.846558, 1.800079, 1.713867, 1.597015, 1.524811, 
    1.379364, 1.291077, 1.116821, 1.005859, 0.9875488, 1.01712, 1.028778, 
    1.040497, 1.040619, 0.9522095, 1.042419, 1.171875, 1.709564, 2.377289, 
    3.47113, 4.90686, 3.158081, 2.115479, 3.112579, 3.365936, 2.884369, 
    2.740234, 2.255127, 2.13385, 2.165924, 2.036072, 1.891724, 1.761475, 
    1.646301, 1.616394, 1.575073, 1.530914, 1.52356,
  1.992584, 2.24057, 2.374542, 2.544922, 3.930725, 4.189972, 3.558136, 
    3.606293, 3.413147, 3.166901, 2.179291, 2.134766, 2.670837, 3.051483, 
    2.466858, 2.410217, 2.245178, 2.159088, 2.162842, 2.144806, 2.048309, 
    1.991669, 1.979797, 1.966339, 1.984833, 2.068207, 2.241089, 2.390259, 
    2.471283, 2.480255, 2.480804, 2.588928, 2.950348, 3.491425, 3.258514, 
    3.060028, 3.137512, 2.855743, 2.412018, 2.085815, 2.098846, 2.118378, 
    2.218994, 2.301819, 2.259827, 2.243469, 2.210022, 2.194244, 2.173553, 
    2.125763, 2.108398, 2.063538, 2.0383, 2.031189, 2.033661, 2.035736, 
    1.99649, 1.922058, 1.859589, 1.771606, 1.709656, 1.601715, 1.516205, 
    1.371613, 1.250977, 1.17807, 1.187408, 1.215363, 1.234955, 1.261139, 
    1.241211, 1.242859, 1.289246, 1.45874, 1.582031, 1.910797, 2.436401, 
    3.7612, 4.11557, 3.140442, 2.39682, 3.02713, 3.578003, 2.989349, 
    2.992645, 2.986908, 2.079956, 2.059509, 1.946869, 1.830658, 1.757813, 
    1.731049, 1.768463, 1.763855, 1.856049, 1.907898,
  2.469269, 2.606567, 2.61676, 2.379669, 3.497528, 4.052612, 3.568756, 
    3.323639, 3.482422, 3.009125, 2.660553, 2.387238, 2.789124, 2.860229, 
    2.485352, 2.324219, 2.167328, 2.184174, 2.27774, 2.290741, 2.245239, 
    2.208282, 2.237305, 2.253387, 2.318115, 2.38913, 2.502991, 2.570038, 
    2.560333, 2.531555, 2.469208, 2.41449, 2.435272, 3.040741, 2.84375, 
    2.260498, 2.537262, 2.3685, 2.564392, 2.093628, 2.162628, 2.258789, 
    2.27179, 2.331177, 2.288666, 2.244781, 2.180237, 2.20163, 2.1828, 
    2.156128, 2.139191, 2.094574, 2.059235, 2.058777, 2.076233, 2.058258, 
    2.062714, 2.004211, 1.955536, 1.8862, 1.837769, 1.720886, 1.68869, 
    1.612823, 1.550598, 1.567963, 1.559753, 1.633148, 1.662384, 1.695557, 
    1.682281, 1.717194, 1.782806, 1.802734, 1.896118, 2.333649, 3.756592, 
    4.488342, 3.419525, 2.975067, 2.828583, 2.74707, 2.824829, 2.762024, 
    3.1427, 2.976318, 2.051117, 2.136383, 2.093506, 2.043304, 2.051697, 
    2.100281, 2.195557, 2.231445, 2.28894, 2.384186,
  2.717133, 2.746918, 2.673248, 2.390381, 2.998108, 3.043823, 2.949921, 
    2.924622, 2.773834, 2.686066, 2.735138, 2.440887, 2.311707, 2.48111, 
    2.472076, 2.333649, 2.180267, 2.223938, 2.329163, 2.386597, 2.358185, 
    2.352936, 2.394592, 2.455139, 2.528778, 2.502228, 2.558197, 2.566071, 
    2.509552, 2.414063, 2.418274, 2.422607, 2.362091, 2.203522, 2.202942, 
    2.529572, 2.749878, 2.161713, 2.295837, 2.067596, 2.150391, 2.333862, 
    2.275848, 2.198303, 2.12558, 2.1185, 2.051117, 2.009583, 2.07962, 
    2.094147, 2.108398, 2.042297, 1.997528, 2.040833, 2.089233, 2.079895, 
    2.159851, 2.132233, 2.079376, 2.084442, 2.064514, 1.989716, 1.972839, 
    1.970825, 1.941284, 1.971039, 2.0047, 2.054688, 2.056488, 2.136383, 
    2.188385, 2.269257, 2.3172, 2.2211, 2.393677, 3.123749, 2.906372, 
    3.067108, 3.029938, 2.846405, 2.677338, 2.766754, 2.797394, 2.815491, 
    3.157227, 2.832123, 2.067322, 2.185791, 2.256256, 2.271027, 2.338684, 
    2.437958, 2.501373, 2.561768, 2.623871, 2.68631,
  2.693756, 2.691986, 2.526093, 2.380219, 3.093964, 3.068237, 2.953644, 
    2.698364, 2.543152, 2.421051, 2.372009, 2.326355, 2.344269, 2.460266, 
    2.401733, 2.308533, 2.281647, 2.37381, 2.460724, 2.498108, 2.466095, 
    2.492371, 2.551361, 2.602142, 2.600525, 2.559113, 2.508392, 2.357941, 
    2.398438, 2.438782, 2.39386, 2.376953, 2.432312, 2.452087, 2.383118, 
    2.404297, 2.22702, 2.175537, 2.24173, 2.039001, 2.145844, 2.235596, 
    2.203766, 2.164001, 2.086548, 2.00943, 1.962677, 1.994507, 2.060547, 
    2.078125, 2.132751, 2.087982, 2.064911, 2.092834, 2.141724, 2.176178, 
    2.187897, 2.173981, 2.162689, 2.200928, 2.199554, 2.187378, 2.172729, 
    2.198425, 2.176178, 2.188812, 2.223846, 2.252014, 2.323883, 2.444916, 
    2.540771, 2.557098, 2.55722, 2.573425, 2.579742, 2.488586, 2.848785, 
    3.089386, 2.954437, 2.849426, 2.677429, 2.795502, 2.650085, 2.855103, 
    3.002747, 2.914764, 3.054688, 2.266479, 2.350952, 2.362244, 2.394012, 
    2.448761, 2.518829, 2.595703, 2.662323, 2.673676,
  2.380615, 2.391479, 2.216522, 2.377472, 4.142639, 3.55896, 3.07251, 
    2.834503, 2.534607, 2.081177, 2.009949, 2.365753, 2.322266, 2.40033, 
    2.460785, 2.444275, 2.434418, 2.518555, 2.527679, 2.537811, 2.538879, 
    2.561249, 2.574554, 2.650116, 2.622986, 2.606842, 2.446991, 2.289764, 
    2.582672, 2.473877, 2.369812, 2.258514, 2.373962, 2.3479, 2.319031, 
    2.402985, 2.225922, 2.556061, 2.67337, 2.755524, 2.156525, 2.183014, 
    2.236664, 2.215942, 2.143097, 2.127838, 2.167694, 2.144928, 2.19519, 
    2.20343, 2.236145, 2.264587, 2.291595, 2.307495, 2.301239, 2.323059, 
    2.31366, 2.333344, 2.307556, 2.303131, 2.286133, 2.284821, 2.281647, 
    2.277161, 2.274536, 2.288025, 2.319061, 2.380676, 2.46875, 2.53125, 
    2.585815, 2.55014, 2.494995, 2.627136, 2.566467, 2.43045, 2.681335, 
    2.936401, 2.68335, 2.655884, 2.864594, 2.867767, 2.73645, 3.244537, 
    3.399292, 2.824829, 2.944122, 2.327209, 2.366669, 2.376312, 2.444397, 
    2.493744, 2.517853, 2.498779, 2.511658, 2.45462,
  2.294678, 2.322113, 2.371704, 3.427673, 4.335541, 3.357666, 3.102386, 
    3.164337, 2.737854, 1.790558, 1.630737, 3.094269, 2.436188, 2.474213, 
    2.518097, 2.535553, 2.512451, 2.462891, 2.487946, 2.518158, 2.499786, 
    2.484558, 2.473053, 2.48587, 2.483856, 2.421997, 2.314911, 2.707733, 
    2.828003, 2.40213, 2.685028, 2.657227, 2.913422, 2.267426, 2.325989, 
    2.841156, 2.700653, 2.371368, 2.266357, 2.059845, 2.057922, 2.036194, 
    2.008942, 2.014282, 2.005402, 2.020844, 1.995239, 1.955933, 1.976746, 
    1.990234, 1.961792, 1.985626, 1.981445, 1.991608, 2.02359, 2.08374, 
    2.160461, 2.241333, 2.298889, 2.384186, 2.464111, 2.504364, 2.560944, 
    2.58548, 2.65155, 2.686249, 2.695251, 2.754486, 2.736389, 2.700073, 
    2.687653, 2.568481, 2.447876, 2.403534, 2.421143, 2.430603, 2.427155, 
    2.536713, 2.532532, 2.077209, 2.682495, 3.015015, 3.405029, 3.885559, 
    3.504669, 2.219299, 2.23526, 2.327972, 2.432098, 2.435486, 2.466003, 
    2.449463, 2.477997, 2.450867, 2.435852, 2.348236,
  2.325928, 2.424164, 2.458862, 3.233459, 3.50943, 3.156464, 3.237305, 
    3.233032, 3.104431, 1.801971, 1.59317, 3.670654, 3.01947, 2.516479, 
    2.490967, 2.602081, 2.5513, 2.534943, 2.508148, 2.477539, 2.493866, 
    2.484497, 2.500275, 2.479492, 2.460297, 2.325531, 2.319031, 3.17981, 
    2.302216, 2.352356, 2.495636, 2.707214, 2.687836, 2.269226, 2.193298, 
    2.208466, 2.024353, 1.960693, 2.047729, 2.144257, 2.116516, 2.031921, 
    2.026825, 2.018616, 2.03064, 2.036987, 1.992554, 1.990295, 1.950928, 
    1.938232, 1.919281, 1.898834, 1.874542, 1.875336, 1.894318, 1.917236, 
    1.969727, 2.055145, 2.156036, 2.255341, 2.353119, 2.442596, 2.525787, 
    2.615875, 2.682983, 2.744263, 2.811066, 2.887909, 2.894531, 2.813934, 
    2.685364, 2.534302, 2.411255, 2.265808, 2.085236, 2.165771, 2.481567, 
    2.089447, 2.12558, 2.462006, 3.353119, 3.622009, 3.277679, 2.16452, 
    2.068878, 2.093811, 2.204163, 2.284485, 2.35318, 2.403625, 2.432556, 
    2.475067, 2.504669, 2.449158, 2.429474, 2.351563,
  3.071411, 2.574951, 3.120514, 3.639313, 3.563599, 3.234497, 3.322449, 
    3.237579, 3.239655, 2.610291, 2.229889, 3.220001, 3.530273, 2.571564, 
    2.581512, 2.680481, 2.638733, 2.63855, 2.585724, 2.592255, 2.531708, 
    2.438995, 2.485229, 2.567261, 2.54068, 2.452606, 3.173065, 3.36673, 
    2.161652, 2.279358, 2.343689, 2.784973, 2.233521, 2.33847, 2.120056, 
    2.131226, 2.124939, 2.17572, 2.234711, 2.235016, 2.2211, 2.204163, 
    2.232422, 2.229095, 2.255249, 2.285736, 2.269928, 2.290619, 2.305603, 
    2.320587, 2.329315, 2.303955, 2.288483, 2.265564, 2.232117, 2.222076, 
    2.232758, 2.230164, 2.213409, 2.217651, 2.223358, 2.271942, 2.292969, 
    2.31366, 2.326904, 2.406769, 2.527618, 2.685944, 2.789764, 2.710632, 
    2.626495, 2.562317, 2.462433, 2.321808, 2.186279, 2.57605, 2.364014, 
    2.697845, 2.706635, 3.750519, 3.60907, 3.125122, 2.506012, 2.061737, 
    2.135284, 2.178955, 2.229309, 2.243561, 2.303589, 2.362366, 2.409485, 
    2.408936, 2.356384, 2.430328, 2.869659, 2.874817,
  3.819336, 3.270294, 3.650848, 3.791199, 3.905548, 4.00351, 3.635223, 
    3.524567, 3.732819, 3.80188, 3.380859, 3.445251, 3.75, 3.275391, 2.49942, 
    2.665192, 2.86319, 2.851776, 2.841064, 2.819458, 2.61795, 2.828064, 
    2.561523, 2.481842, 2.377014, 2.274017, 2.453644, 3.159851, 2.18158, 
    2.191986, 2.172333, 2.129822, 2.171814, 2.759369, 2.232269, 2.273376, 
    2.315765, 2.330078, 2.364197, 2.360474, 2.377411, 2.409241, 2.410492, 
    2.421478, 2.448761, 2.451355, 2.509308, 2.536987, 2.576996, 2.584747, 
    2.600861, 2.609161, 2.590637, 2.616974, 2.595825, 2.562897, 2.539703, 
    2.490021, 2.418091, 2.382813, 2.317383, 2.287048, 2.283844, 2.303955, 
    2.314911, 2.354675, 2.450439, 2.646332, 2.764252, 2.711639, 2.62793, 
    2.570557, 2.684509, 2.804413, 2.712097, 3.055939, 3.544037, 2.995239, 
    3.358978, 3.257751, 2.283966, 2.358124, 2.376709, 2.21405, 2.170654, 
    2.16153, 2.190033, 2.232819, 2.265625, 2.324097, 2.402405, 2.375275, 
    2.469849, 3.788666, 3.975128, 3.871552,
  3.750183, 3.576233, 3.656647, 3.656067, 3.731262, 3.643372, 3.533783, 
    3.532227, 3.420502, 3.90033, 4.115875, 3.734955, 3.587372, 3.361084, 
    2.524597, 2.493561, 2.742493, 2.858795, 2.960297, 2.894928, 3.753784, 
    3.962952, 2.689056, 2.583862, 2.480072, 2.295715, 2.31842, 3.202545, 
    3.615692, 3.295624, 2.124298, 2.117706, 2.186218, 2.769775, 2.239441, 
    2.312958, 2.334686, 2.333527, 2.369781, 2.353241, 2.347931, 2.350433, 
    2.355133, 2.363708, 2.414246, 2.44043, 2.458252, 2.503326, 2.564972, 
    2.634247, 2.665161, 2.656128, 2.64389, 2.675629, 2.659302, 2.649933, 
    2.632416, 2.548767, 2.480103, 2.413544, 2.356384, 2.330017, 2.342316, 
    2.371674, 2.378601, 2.349152, 2.358917, 2.497589, 2.601105, 2.668365, 
    2.624634, 2.712067, 3.34433, 3.249146, 2.544739, 2.699585, 2.69809, 
    2.516693, 2.436646, 2.357422, 2.230988, 2.302856, 2.230011, 2.213013, 
    2.177551, 2.2117, 2.210754, 2.241608, 2.229279, 2.306244, 2.409515, 
    2.635406, 3.384308, 3.584442, 3.678375, 3.709106,
  3.847717, 4.112213, 4.264954, 4.265228, 4.006653, 3.650452, 3.691528, 
    3.709259, 3.782104, 3.722534, 3.881958, 4.14975, 3.549194, 3.307465, 
    3.061279, 2.638733, 2.549469, 2.62384, 2.861511, 2.804291, 4.040466, 
    4.413849, 2.808533, 2.727875, 2.646179, 2.651245, 3.603516, 3.091522, 
    2.45517, 1.798248, 1.94278, 1.987244, 1.873047, 1.922974, 2.082611, 
    2.202484, 2.23587, 2.258118, 2.275757, 2.27298, 2.268951, 2.234161, 
    2.239594, 2.211609, 2.226227, 2.29245, 2.297974, 2.32489, 2.362823, 
    2.425598, 2.467651, 2.507751, 2.53894, 2.522064, 2.523315, 2.524139, 
    2.510986, 2.448303, 2.367035, 2.273132, 2.185333, 2.136597, 2.147583, 
    2.208984, 2.288483, 2.219391, 2.042114, 2.138611, 2.549408, 4.294678, 
    3.952148, 4.580933, 4.093597, 2.212097, 2.423553, 2.455658, 2.420776, 
    2.399353, 2.286835, 2.247467, 2.213806, 2.175873, 2.140961, 2.093903, 
    2.072388, 2.07962, 2.05603, 2.074738, 2.064392, 2.151886, 2.281372, 
    2.795624, 3.804749, 3.61792, 3.630524, 3.62207,
  3.685089, 3.948425, 4.087708, 4.0784, 4.099884, 4.071991, 4.058014, 
    3.882416, 4.010223, 3.540741, 2.373505, 4.096558, 4.284119, 3.808716, 
    3.8125, 3.618866, 2.534821, 2.555084, 2.879608, 2.80188, 4.219849, 
    4.182404, 4.076691, 4.004944, 2.828186, 3.368896, 3.417816, 3.027802, 
    1.511597, 1.059326, 1.870972, 2.024139, 1.871765, 1.781372, 1.806366, 
    1.917358, 1.969421, 2.01825, 2.034637, 2.051178, 2.07077, 2.040771, 
    2.046875, 2.026886, 1.994202, 2.038727, 2.064117, 2.149628, 2.209625, 
    2.230713, 2.278137, 2.291809, 2.29245, 2.305359, 2.317383, 2.296753, 
    2.284454, 2.255524, 2.174988, 2.068604, 1.964325, 1.867126, 1.845367, 
    1.873627, 1.968353, 1.873505, 1.755402, 2.255646, 4.8078, 4.483856, 
    3.312164, 3.312317, 3.395447, 2.03183, 2.221924, 2.251892, 2.252716, 
    2.307404, 2.217194, 2.201874, 2.160797, 2.108521, 2.05307, 1.947632, 
    1.93222, 1.918243, 1.876801, 1.860809, 1.765869, 1.739471, 1.829895, 
    2.410797, 3.761841, 3.536194, 3.377167, 3.551056,
  3.334442, 3.653503, 3.949066, 4.04837, 3.993805, 3.783142, 3.816467, 
    3.630585, 3.613159, 3.582947, 2.321411, 4.251801, 4.398621, 4.600128, 
    4.723114, 4.114929, 2.858337, 2.98822, 4.37619, 4.339844, 4.440247, 
    3.95871, 3.813995, 3.949738, 4.058655, 3.963715, 4.115753, 3.345398, 
    1.687439, 0.848175, 1.048492, 1.14566, 1.782349, 1.798706, 1.806183, 
    1.865234, 1.951569, 2.013824, 2.007477, 2.0047, 2.022339, 2.034241, 
    1.972931, 1.926758, 1.850983, 1.795837, 1.744904, 1.765869, 1.806885, 
    1.876373, 2.008789, 2.061707, 2.122925, 2.164063, 2.131439, 2.152161, 
    2.166351, 2.142761, 2.147858, 2.094543, 2.02356, 1.95105, 1.91275, 
    1.93689, 2.012695, 1.830353, 2.101746, 4.162903, 4.670166, 4.138947, 
    3.141968, 2.325897, 2.085022, 1.989014, 2.03418, 2.006134, 2.021271, 
    2.155945, 2.364594, 2.388458, 2.34549, 2.353638, 2.3125, 2.238861, 
    2.203064, 2.078644, 2.004517, 1.947906, 1.783203, 1.708527, 1.728882, 
    1.921631, 3.128052, 3.436371, 3.388214, 3.323761,
  3.127075, 3.305603, 3.577454, 3.85553, 3.932037, 3.744141, 3.888214, 
    3.7547, 3.482422, 3.952332, 3.877472, 4.002625, 4.088654, 4.711578, 
    5.379242, 4.934143, 4.822784, 5.387817, 5.271301, 4.934753, 5.028503, 
    4.579498, 4.154053, 3.274506, 4.083282, 4.078552, 5.104889, 3.025909, 
    2.017914, 2.250397, 2.564514, 1.860657, 1.598633, 1.80307, 1.921661, 
    1.886536, 1.922211, 2.036133, 2.067841, 2.055206, 2.03418, 2.035309, 
    1.9823, 1.886414, 1.799225, 1.752472, 1.721558, 1.688995, 1.665497, 
    1.668701, 1.753174, 1.820648, 1.877716, 1.920746, 1.941986, 2.012451, 
    2.021881, 2.010437, 1.998749, 2.001617, 1.97345, 1.942688, 1.922516, 
    1.974487, 1.900391, 2.026184, 3.216644, 3.891418, 4.020874, 4.065308, 
    3.722931, 2.653839, 2.406708, 2.378784, 2.211243, 1.96225, 1.954224, 
    1.984039, 2.096619, 2.182343, 2.288483, 2.387634, 2.393646, 2.389771, 
    2.362823, 2.328705, 2.293304, 2.228363, 2.111877, 1.94516, 1.752686, 
    1.701935, 2.030884, 2.81662, 3.221863, 3.139008,
  3.358246, 3.365692, 3.325256, 3.480804, 3.577667, 2.759918, 3.745331, 
    3.709961, 2.852692, 4.009125, 4.035797, 3.973328, 4.288208, 4.803314, 
    4.711792, 4.282806, 4.534424, 4.911011, 4.795898, 5.962952, 5.817261, 
    7.237061, 5.429718, 4.285309, 4.349701, 5.74585, 4.192413, 2.446411, 
    2.616119, 4.447327, 5.032501, 4.279022, 2.682892, 1.181335, 1.722504, 
    1.993622, 1.905579, 2.010742, 2.044556, 2.056458, 2.071136, 2.061462, 
    2.035156, 1.999481, 1.931519, 1.855469, 1.792694, 1.757599, 1.727936, 
    1.684052, 1.707428, 1.745758, 1.765045, 1.819672, 1.865784, 1.86203, 
    1.864136, 1.874329, 1.867004, 1.881287, 1.913086, 1.855682, 1.864166, 
    1.939758, 2.009247, 2.992584, 3.808838, 3.956512, 3.952148, 3.740631, 
    3.326019, 2.502686, 2.13736, 2.022064, 2.032562, 1.846344, 1.85788, 
    1.902985, 1.971588, 1.945129, 1.944855, 1.998108, 2.0896, 2.15097, 
    2.160675, 2.185181, 2.204895, 2.216919, 2.251312, 2.202209, 2.037903, 
    1.863342, 1.845978, 2.028137, 2.669006, 2.977386,
  3.10553, 3.493286, 3.32312, 2.753113, 2.607086, 2.501892, 2.502686, 
    2.525726, 2.75351, 2.961639, 4.013794, 4.903168, 4.88562, 4.271545, 
    4.037903, 3.749268, 3.878632, 4.421539, 4.862946, 6.297089, 6.269928, 
    6.228912, 5.02298, 4.59903, 4.976013, 3.286926, 2.910065, 3.367462, 
    3.1362, 3.327026, 3.031433, 3.413666, 2.917084, 1.372406, 2.787354, 
    2.224945, 2.187592, 2.630341, 2.158417, 2.114807, 2.11615, 2.142853, 
    2.153412, 2.107697, 2.075653, 2.081055, 2.074677, 2.039276, 2.010284, 
    1.990356, 1.941132, 1.8685, 1.801514, 1.780731, 1.761047, 1.779175, 
    1.819, 1.812439, 1.769135, 1.785431, 1.813171, 1.813019, 1.860229, 
    1.945587, 2.483063, 2.81424, 3.092041, 2.922333, 3.512695, 3.585419, 
    3.047028, 2.540131, 2.333984, 2.200439, 2.286926, 2.344177, 2.165833, 
    2.02533, 2.004303, 2.074677, 2.174957, 2.120697, 1.940491, 1.836823, 
    1.758453, 1.692383, 1.672272, 1.661804, 1.752228, 2.035614, 2.174988, 
    1.993774, 1.794983, 1.799866, 2.01825, 2.748779,
  2.612762, 2.35968, 2.462952, 2.43689, 2.443237, 2.391357, 3.050323, 
    3.285522, 3.536407, 3.56311, 3.882477, 5.287109, 3.761993, 3.231964, 
    2.478516, 2.923309, 3.99472, 3.971283, 3.035156, 4.445129, 3.760773, 
    1.916077, 1.355408, 1.341949, 2.543976, 1.917542, 2.609436, 2.735046, 
    2.102478, 1.91098, 2.243103, 1.962708, 1.675873, 2.086517, 2.481445, 
    2.311615, 2.252655, 2.751831, 2.303986, 2.334686, 2.384979, 2.409729, 
    2.475861, 2.467133, 2.398315, 2.344452, 2.318451, 2.262024, 2.185089, 
    2.154114, 2.127136, 2.084961, 1.991791, 1.917786, 1.890961, 1.872467, 
    1.856384, 1.813477, 1.831573, 1.847321, 1.840424, 1.868561, 1.902008, 
    2.012939, 2.98761, 3.820313, 4.123108, 3.41922, 2.736267, 3.514374, 
    3.4422, 3.209534, 3.133148, 3.124603, 3.2211, 3.453308, 3.483398, 
    2.998291, 2.796875, 2.829834, 2.773224, 2.619812, 2.256592, 1.577606, 
    0.9057312, 0.852478, 0.9460754, 0.8582764, 0.8898621, 1.243805, 1.773315, 
    1.902924, 1.8526, 1.887939, 2.150909, 2.405914,
  2.4617, 2.302094, 2.40802, 2.690094, 2.490234, 3.114838, 3.886261, 
    3.657959, 3.707733, 3.638672, 3.624359, 5.098389, 4.490631, 2.469727, 
    2.722717, 2.908142, 2.399017, 3.102081, 3.025909, 2.2742, 2.381012, 
    1.960419, 1.829193, 1.603912, 1.96994, 1.872192, 2.288483, 2.075989, 
    1.921478, 1.86087, 1.714325, 1.707367, 1.930481, 2.208527, 2.39502, 
    2.107513, 2.348999, 2.33667, 3.267975, 3.405487, 3.623779, 3.264984, 
    2.704559, 2.425171, 2.286987, 2.223053, 2.206512, 2.295441, 2.366333, 
    2.30246, 2.20105, 2.130798, 2.116211, 2.108521, 2.077484, 2.02951, 
    1.989838, 1.951752, 1.901367, 1.869415, 1.890991, 1.853912, 1.815613, 
    2.068024, 4.14682, 5.00058, 4.416565, 3.3815, 2.356964, 1.943176, 
    2.433197, 2.678009, 3.129211, 3.533203, 3.621338, 4.167053, 4.399933, 
    4.30188, 4.718445, 4.344482, 3.506256, 2.726044, 2.320099, 1.643097, 
    1.114594, 0.7253418, 0.6300049, 0.3764343, 0.2502747, 0.6706848, 
    1.144348, 1.511932, 1.738495, 1.775848, 1.92981, 2.567963,
  2.25177, 2.629486, 3.509552, 3.776428, 2.95462, 3.291016, 3.538483, 
    3.396881, 3.284058, 3.191803, 2.937164, 3.146545, 2.961212, 2.094879, 
    2.015503, 1.456635, 1.454803, 1.68103, 1.815826, 1.653259, 1.684845, 
    1.98114, 2.101044, 1.952209, 2.028839, 1.890564, 2.410889, 2.795837, 
    2.44043, 2.426758, 2.584045, 2.859711, 3.038361, 3.195313, 2.521454, 
    2.536072, 2.529114, 2.38739, 2.751892, 3.060272, 2.95163, 2.532288, 
    2.470886, 2.332367, 2.246155, 2.142395, 2.124176, 2.205078, 2.25769, 
    2.235046, 2.214569, 2.235046, 2.273438, 2.261444, 2.146057, 2.004883, 
    1.948944, 1.968475, 1.971436, 1.983124, 2.0354, 1.962311, 1.970856, 
    2.259308, 3.993103, 3.278717, 3.516815, 3.311371, 2.494659, 2.239502, 
    2.704559, 3.274017, 4.009857, 6.252686, 4.474579, 4.159393, 3.881073, 
    3.917542, 4.266174, 5.037109, 3.723053, 2.98349, 2.67746, 1.890167, 
    1.316345, 1.10788, 0.6617737, 0.01159668, -0.4124451, -0.2012634, 
    0.4439392, 1.055725, 1.497711, 1.657104, 1.901123, 2.106964,
  2.046783, 2.311798, 2.917572, 3.336334, 3.114014, 3.271423, 3.523346, 
    3.345764, 3.834717, 4.032043, 3.784515, 3.408875, 2.75058, 2.078339, 
    2.084442, 1.973938, 1.565308, 1.60144, 1.977173, 1.848267, 2.089447, 
    2.092377, 2.618378, 2.947601, 2.524475, 2.094086, 2.721436, 2.830109, 
    2.662781, 2.762787, 3.303192, 3.108673, 2.68158, 2.520477, 2.492218, 
    2.09845, 1.614075, 2.593384, 5.245575, 8.569214, 5.888428, 3.751495, 
    2.834045, 2.590942, 2.588135, 2.350464, 2.378967, 2.466736, 2.432373, 
    2.401489, 2.418945, 2.471863, 2.516602, 2.463165, 2.383118, 2.268372, 
    2.070465, 2.013611, 2.100464, 2.106171, 2.074158, 2.071869, 2.231232, 
    2.527405, 2.884338, 2.687775, 3.641937, 3.303253, 3.329132, 3.858307, 
    3.783081, 3.503723, 3.562378, 3.895264, 4.116608, 3.983734, 4.029633, 
    4.096039, 4.067017, 3.966309, 5.858276, 5.107452, 5.179626, 2.702423, 
    1.744476, 1.125397, 0.2915955, -0.6752014, -1.299072, -1.154633, 
    -0.3695984, 0.559845, 1.228638, 1.483154, 1.606049, 1.696106,
  1.940887, 1.756989, 2.084442, 2.243744, 2.64679, 3.076172, 3.530609, 
    3.942322, 3.78009, 3.432373, 3.186615, 2.811401, 2.473083, 2.166168, 
    1.900909, 1.807373, 1.863617, 1.933472, 1.93927, 2.299286, 2.345581, 
    2.821045, 2.756989, 2.885101, 2.751862, 2.490448, 2.446289, 2.519989, 
    2.617279, 2.876709, 3.136536, 3.03511, 2.920914, 2.746368, 2.65242, 
    2.209839, 1.832047, 2.785431, 4.989227, 8.474304, 7.630798, 5.662537, 
    3.943298, 3.299561, 3.329742, 2.647095, 2.425598, 2.341217, 2.36499, 
    2.428131, 2.669189, 3.021484, 3.248627, 2.984375, 2.607422, 2.568024, 
    2.299347, 2.214508, 2.199219, 2.127014, 1.932922, 2.636871, 2.607941, 
    2.667145, 2.598053, 2.6633, 3.240601, 3.408478, 3.870789, 3.905304, 
    4.096039, 4.348663, 4.895569, 5.300659, 4.956268, 5.506317, 4.812958, 
    4.43544, 3.843246, 3.566437, 4.481995, 6.438416, 6.523438, 2.394012, 
    1.156067, 1.12381, 0.6714783, -0.2675171, -1.036072, -1.033722, 
    -0.3668823, 0.5246887, 1.143738, 1.323181, 1.382751, 1.680939,
  1.257874, 1.379333, 1.340027, 2.940094, 3.174683, 3.105743, 3.221863, 
    3.529236, 2.97464, 2.839081, 2.933136, 2.904907, 2.369812, 1.977814, 
    1.78244, 1.928833, 1.829895, 1.841766, 1.739563, 2.223053, 2.651398, 
    2.697601, 3.282501, 3.364166, 3.25061, 2.967072, 2.804291, 2.902954, 
    2.860565, 2.861481, 2.926651, 3.125854, 3.208359, 3.100006, 2.64917, 
    2.540771, 2.709137, 3.667084, 5.125427, 6.803925, 6.344482, 4.973755, 
    4.616287, 4.858154, 6.781525, 4.246185, 4.603973, 5.206207, 4.956451, 
    5.401611, 6.08905, 5.939514, 4.954285, 4.14798, 4.024689, 2.61322, 
    2.398499, 2.286011, 2.157898, 1.991272, 2.889404, 3.069031, 2.857391, 
    2.629333, 2.812256, 3.170593, 3.301971, 3.403381, 3.522339, 4.026123, 
    4.668457, 5.232697, 5.694672, 5.877747, 5.799561, 5.700073, 5.329437, 
    4.927536, 4.176132, 3.842102, 4.207581, 5.80069, 4.352875, 0.1266479, 
    -0.1167603, 1.114838, 1.572662, 1.167175, 0.5915833, 0.434906, 0.6733704, 
    0.9893494, 1.21521, 1.33255, 1.364624, 1.616211,
  0.9414063, 1.115814, 2.566437, 2.972015, 3.700073, 5.326019, 3.700989, 
    3.570007, 3.277222, 3.089722, 3.053467, 2.943878, 2.692078, 2.19635, 
    1.891754, 1.926239, 2.215302, 2.362457, 2.305084, 2.439987, 2.50769, 
    3.148407, 3.554047, 3.64624, 3.792252, 3.599823, 3.724686, 3.66127, 
    3.548782, 3.328857, 3.338043, 3.3284, 3.315109, 3.110184, 2.937836, 
    2.905624, 2.785355, 2.992981, 3.026062, 3.08432, 3.302689, 3.352219, 
    3.969162, 4.826843, 5.971436, 7.16687, 8.834061, 13.59727, 14.10046, 
    12.77222, 11.16208, 9.362457, 6.642334, 4.977356, 3.77417, 3.058472, 
    2.748505, 2.554382, 2.629456, 2.683929, 2.570007, 2.563873, 2.582031, 
    2.77002, 3.029968, 3.34668, 3.586304, 3.737534, 4.074036, 4.732117, 
    5.283813, 5.458145, 5.712875, 5.911255, 5.929337, 5.773346, 5.456467, 
    4.745529, 3.582245, 3.432312, 3.456604, 3.605209, 2.400024, 1.774963, 
    2.504913, 1.049103, 1.186981, 1.373169, 1.641541, 1.761597, 1.719391, 
    1.293488, 0.4902954, 0.3344421, 0.8104248, 0.9119873,
  0.5993958, 0.7445374, 0.8446655, 3.20993, 3.923706, 4.326538, 5.00412, 
    4.309326, 4.211151, 4.10321, 3.971313, 3.943909, 3.731079, 3.294678, 
    2.982971, 2.780075, 2.956787, 3.427887, 3.557831, 3.691086, 3.742661, 
    3.977554, 4.113831, 4.156128, 4.359268, 4.195267, 4.177689, 4.356339, 
    4.300735, 4.19194, 4.082443, 3.663696, 3.598785, 3.560165, 3.423721, 
    3.481583, 3.666107, 3.284775, 3.099106, 3.19635, 3.362686, 4.051056, 
    4.672729, 5.097015, 5.381668, 5.620071, 6.075867, 6.608612, 7.119934, 
    7.199173, 7.077957, 6.874954, 5.798126, 4.75444, 3.856018, 3.300537, 
    2.840454, 2.751907, 2.845581, 2.92009, 3.057831, 3.301651, 3.446167, 
    3.748276, 3.770828, 3.979462, 4.375504, 4.729019, 4.980118, 5.136246, 
    5.031235, 5.255417, 5.43692, 5.635376, 5.631973, 5.366104, 4.859711, 
    4.273056, 4.081131, 4.021103, 3.573898, 3.430481, 3.530289, 3.834183, 
    4.221237, 4.239136, 3.762787, 2.270721, 1.484589, 2.939789, 5.255035, 
    5.436798, 2.930145, 1.17572, 0.4580078, 0.428833,
  0.9482422, 0.6158752, 0.5211792, 0.4916077, -0.07336426, 2.973511, 
    3.675232, 4.525879, 5.254501, 5.916031, 6.189651, 6.549866, 5.876007, 
    4.865982, 4.14325, 3.969223, 3.994873, 4.165695, 4.476898, 4.581787, 
    4.56955, 4.638168, 4.800735, 4.869156, 4.886017, 5.141754, 4.694458, 
    4.425262, 4.097809, 4.115814, 4.280334, 4.197205, 4.036316, 3.784622, 
    3.930206, 3.749802, 3.349609, 3.73822, 3.641937, 3.968872, 4.149414, 
    4.371033, 4.762115, 5.16745, 5.904755, 6.172974, 6.743225, 7.34375, 
    7.578049, 7.360107, 7.801453, 7.891815, 7.701324, 6.470779, 5.844681, 
    5.232117, 4.859909, 4.751129, 4.622055, 4.3134, 4.112167, 4.004807, 
    4.269119, 4.28801, 4.372055, 4.428177, 4.690903, 4.959854, 5.29657, 
    5.037491, 5.334259, 5.258255, 5.297134, 4.983597, 5.406326, 4.97261, 
    5.242508, 5.012039, 4.827927, 4.131973, 3.516159, 3.189865, 3.857834, 
    4.924042, 5.366272, 5.004166, 4.030792, 4.03244, 4.652359, 5.710114, 
    6.790878, 7.621109, 8.741882, 8.884003, 4.160065, 1.847534,
  3.234985, 1.810425, 1.237152, 1.078125, 1.02832, 1.442322, 2.603485, 
    4.695984, 8.097931, 10.76532, 11.47188, 10.41023, 8.705551, 6.870529, 
    5.889069, 5.240845, 4.755692, 4.965698, 5.061081, 5.010422, 5.001053, 
    4.998703, 5.12175, 5.217514, 5.181183, 5.095566, 4.94928, 4.653458, 
    4.600708, 4.564774, 4.53978, 4.620056, 4.604416, 4.551559, 4.475723, 
    3.761078, 4.283981, 4.314331, 5.196152, 5.429565, 4.914703, 5.200851, 
    5.211594, 5.223953, 5.314072, 5.513412, 5.694916, 5.899612, 6.086212, 
    6.182938, 6.214142, 6.241943, 6.236542, 6.156662, 6.209839, 6.23381, 
    6.235443, 6.173508, 6.017197, 5.809265, 5.667496, 5.425125, 5.013138, 
    4.866821, 4.628204, 4.786072, 5.002075, 5.062378, 5.310226, 5.027557, 
    5.609756, 5.93782, 5.025665, 5.863205, 5.879166, 5.650726, 5.302612, 
    4.535095, 4.444427, 4.397018, 3.964005, 4.529053, 4.770004, 5.100327, 
    5.251831, 4.867188, 4.206909, 3.76973, 3.578262, 3.947739, 4.676437, 
    5.462387, 6.097763, 6.489594, 6.622345, 6.646301,
  6.231323, 5.100983, 3.798065, 4.388092, 6.607361, 10.05203, 9.937515, 
    9.69072, 9.109573, 8.31633, 7.767441, 7.069214, 6.436417, 5.942398, 
    5.672729, 5.58902, 5.581467, 5.745895, 5.867126, 5.807419, 5.70488, 
    5.675461, 5.607422, 5.709305, 5.671112, 6.074875, 5.994461, 5.570251, 
    5.570175, 5.576889, 5.363083, 4.521942, 4.387634, 4.3013, 4.247986, 
    4.492767, 4.747131, 4.908066, 5.108261, 5.231506, 5.327087, 5.409576, 
    5.342957, 5.272461, 5.191727, 5.141861, 5.149994, 5.267975, 5.399033, 
    5.553574, 5.680862, 5.814255, 5.920776, 6.006256, 6.087173, 6.072983, 
    5.990173, 5.869339, 5.787308, 5.808533, 5.869202, 5.946213, 6.055466, 
    6.140106, 6.132736, 5.812042, 5.724487, 5.67363, 5.588867, 5.620453, 
    5.695908, 5.768616, 5.839386, 6.062897, 5.986328, 5.038025, 5.291077, 
    4.856186, 5.729355, 5.083603, 4.621155, 4.249603, 4.109634, 4.061584, 
    4.211578, 4.486908, 4.501434, 4.119659, 3.694138, 3.702209, 4.067123, 
    4.545563, 4.881638, 5.237839, 5.656113, 6.268875,
  5.398117, 5.661087, 6.053986, 6.645889, 6.226364, 6.329819, 6.351959, 
    6.179428, 6.037766, 5.757935, 5.492508, 5.313538, 5.225906, 5.283981, 
    5.456573, 5.659317, 5.861526, 6.010223, 6.113678, 6.157288, 6.140686, 
    6.088928, 5.972198, 5.863998, 5.795441, 6.104233, 6.213287, 5.636002, 
    5.764053, 5.734177, 5.587097, 5.592514, 5.625259, 5.572083, 5.415359, 
    5.261978, 5.172974, 5.059891, 5.028381, 4.990433, 4.901886, 4.837112, 
    4.801102, 4.832214, 4.910873, 5.045059, 5.244781, 5.450653, 5.657089, 
    5.79921, 5.884766, 5.936844, 5.916016, 5.838028, 5.732483, 5.618103, 
    5.610229, 5.629623, 5.610031, 5.592575, 5.626892, 5.641922, 5.695969, 
    5.755722, 5.886002, 5.917572, 5.880325, 5.9142, 5.885025, 5.973969, 
    5.94986, 5.744858, 5.782883, 5.982224, 5.878189, 5.697266, 5.488159, 
    5.253769, 5.020782, 4.735092, 4.430588, 4.206177, 3.966537, 3.844986, 
    3.797455, 3.838531, 3.973892, 4.024872, 4.082428, 4.294022, 4.572861, 
    4.863541, 5.069397, 5.036575, 5.141602, 5.249924,
  5.208984, 5.124146, 5.104492, 5.046555, 4.894714, 4.861725, 4.861862, 
    4.865829, 4.884644, 4.921616, 4.989914, 5.059052, 5.13385, 5.244278, 
    5.344849, 5.382156, 5.388809, 5.413879, 5.445709, 5.481384, 5.495636, 
    5.476624, 5.452667, 5.407883, 5.39122, 5.348694, 5.303452, 5.248306, 
    5.299362, 5.351242, 5.364517, 5.35788, 5.340424, 5.298035, 5.276108, 
    5.177139, 5.095963, 5.050461, 5.011002, 4.952927, 4.931122, 4.956375, 
    5.018433, 5.0513, 5.106644, 5.21283, 5.288986, 5.372528, 5.493027, 
    5.605026, 5.719727, 5.810806, 5.886185, 5.976639, 6.018417, 6.03215, 
    6.006241, 5.954041, 5.922974, 5.9254, 5.931763, 5.972855, 5.98822, 
    6.044724, 6.121414, 6.211792, 6.249542, 6.279556, 6.311005, 6.359039, 
    6.401688, 6.42572, 6.524216, 6.633652, 6.662506, 6.649734, 6.666016, 
    6.65332, 6.733856, 6.712494, 6.760101, 6.639786, 6.64537, 6.498886, 
    6.505066, 6.576965, 6.490311, 6.42662, 6.37233, 6.143158, 5.970261, 
    5.836197, 5.692902, 5.532806, 5.39328, 5.299408,
  5.902344, 5.893173, 5.858337, 5.824738, 5.778976, 5.783386, 5.754562, 
    5.7155, 5.684891, 5.652084, 5.637955, 5.619919, 5.61647, 5.541016, 
    5.483139, 5.468353, 5.391479, 5.367188, 5.370697, 5.375, 5.385223, 
    5.38028, 5.382492, 5.347916, 5.333008, 5.357101, 5.3806, 5.405457, 
    5.437317, 5.434448, 5.462631, 5.525848, 5.560089, 5.562683, 5.580017, 
    5.626816, 5.660553, 5.723434, 5.762375, 5.815811, 5.888931, 5.981171, 
    6.051178, 6.109955, 6.153976, 6.19278, 6.23848, 6.278259, 6.317902, 
    6.347015, 6.333267, 6.31868, 6.332809, 6.330078, 6.327805, 6.32428, 
    6.310165, 6.328461, 6.32695, 6.317184, 6.319534, 6.230469, 6.171677, 
    6.205276, 6.245377, 6.301437, 6.337112, 6.367447, 6.342392, 6.379761, 
    6.386398, 6.373245, 6.377014, 6.429825, 6.458984, 6.432678, 6.450317, 
    6.465881, 6.480591, 6.482681, 6.478378, 6.478119, 6.475189, 6.460861, 
    6.442703, 6.40892, 6.387436, 6.365952, 6.320572, 6.273376, 6.251175, 
    6.195908, 6.134766, 6.062302, 5.993942, 5.939072,
  3.460251, 3.451065, 3.442551, 3.431732, 3.421387, 3.413513, 3.410507, 
    3.411423, 3.416504, 3.431808, 3.448669, 3.466446, 3.488052, 3.504074, 
    3.516953, 3.521713, 3.517349, 3.506866, 3.487976, 3.452774, 3.405182, 
    3.344238, 3.273209, 3.197174, 3.119965, 3.047562, 2.98259, 2.925491, 
    2.874847, 2.834152, 2.799438, 2.768845, 2.74826, 2.732315, 2.716431, 
    2.714615, 2.719177, 2.724258, 2.728485, 2.731277, 2.732712, 2.731155, 
    2.725418, 2.716049, 2.706604, 2.697174, 2.690277, 2.674057, 2.658112, 
    2.657715, 2.644623, 2.635834, 2.640717, 2.695618, 2.635056, 2.666504, 
    2.739548, 2.744492, 2.629196, 2.579147, 2.56221, 2.727051, 2.646591, 
    2.690781, 2.686356, 2.687012, 2.693726, 2.719498, 2.740585, 2.712204, 
    2.720551, 2.73558, 2.756866, 2.905365, 2.87114, 2.916763, 2.990005, 
    3.110382, 3.106873, 3.187332, 3.245407, 3.297623, 3.33493, 3.374115, 
    3.396912, 3.420532, 3.440201, 3.459534, 3.47406, 3.485123, 3.491302, 
    3.493454, 3.488708, 3.485382, 3.480164, 3.46994,
  2.941177, 2.883957, 2.858688, 2.861038, 2.901596, 2.99353, 3.122635, 
    3.283432, 3.471008, 3.676605, 3.880707, 4.087357, 4.257019, 4.370804, 
    4.393219, 4.361496, 4.298813, 4.198288, 4.057465, 3.889694, 3.733643, 
    3.577133, 3.447845, 3.354156, 3.310532, 3.285202, 3.266785, 3.252914, 
    3.242935, 3.22406, 3.193726, 3.147369, 3.098022, 3.047165, 2.995422, 
    2.949326, 2.900162, 2.849777, 2.795471, 2.74086, 2.698013, 2.638702, 
    2.59053, 2.537064, 2.51564, 2.526321, 2.545395, 2.593307, 2.659393, 
    2.749496, 2.841949, 2.848312, 2.973846, 2.966354, 3.356018, 3.023651, 
    3.071243, 3.10405, 3.099686, 3.058289, 2.99884, 2.910187, 2.843704, 
    2.759964, 2.718521, 2.693451, 2.690918, 2.749908, 2.844696, 2.852371, 
    2.750366, 2.549194, 2.402832, 2.324249, 2.430237, 2.490524, 2.57283, 
    2.649521, 2.757782, 2.850433, 2.961945, 3.019623, 3.136108, 3.133942, 
    3.302567, 3.357651, 3.379257, 3.409988, 3.404587, 3.391113, 3.367615, 
    3.319748, 3.245285, 3.161362, 3.072174, 2.998993,
  2.651459, 2.536285, 2.498077, 2.542999, 2.727112, 3.059158, 3.426025, 
    3.780716, 4.037292, 4.117111, 4.094376, 4.077728, 4.095032, 4.080963, 
    4.00824, 3.92601, 3.849258, 3.773926, 3.759735, 3.849197, 4.055847, 
    4.37056, 4.712097, 4.915863, 4.852188, 4.577255, 4.303833, 4.183899, 
    4.105515, 4.013397, 3.920685, 3.793594, 3.571716, 3.287003, 3.041245, 
    2.906281, 2.859406, 2.827774, 2.789627, 2.749451, 2.712021, 2.701859, 
    2.716873, 2.766937, 2.696121, 2.526138, 2.334076, 2.361694, 2.547821, 
    2.663818, 2.738098, 2.737961, 2.659653, 2.591492, 2.577499, 2.531464, 
    2.460831, 2.513748, 2.576645, 2.57431, 2.579453, 2.585892, 2.664215, 
    2.748322, 2.781067, 2.773911, 2.691513, 2.587402, 2.574051, 2.555237, 
    2.446945, 2.318237, 2.182495, 2.118042, 2.121628, 2.217407, 2.325668, 
    2.39299, 2.517731, 2.665451, 2.813828, 2.988174, 3.254837, 3.468246, 
    3.48172, 3.335312, 3.182373, 2.969666, 2.929703, 2.999695, 3.08934, 
    3.139786, 3.137085, 3.076782, 2.948013, 2.797821,
  2.763321, 2.76149, 2.99762, 3.450226, 3.95517, 4.301331, 4.364029, 
    4.058426, 3.565781, 3.195679, 3.128876, 3.401016, 3.783112, 4.116577, 
    4.312988, 4.536484, 4.733612, 5.054001, 5.341492, 4.936218, 4.173996, 
    3.564804, 3.169571, 2.97731, 3.226212, 3.712158, 3.837753, 3.730194, 
    3.671341, 3.62674, 3.569061, 3.437088, 3.317825, 3.293274, 3.31897, 
    3.353683, 3.332138, 3.268204, 3.15596, 2.955826, 2.69574, 2.475235, 
    2.356537, 2.431778, 2.673187, 2.851517, 2.346176, 2.474167, 2.638428, 
    2.746109, 2.805801, 2.811096, 2.773193, 2.742981, 2.71727, 2.705475, 
    2.820663, 2.528931, 2.614792, 2.688293, 2.843567, 2.963242, 2.916946, 
    2.838745, 2.693375, 2.674179, 2.641357, 2.66153, 2.631653, 2.528915, 
    2.457504, 2.310623, 2.178467, 2.17482, 2.315445, 2.476059, 2.733078, 
    2.96376, 3.248917, 3.403671, 3.825272, 4.144424, 4.484909, 4.6978, 
    4.798523, 4.852158, 4.914673, 4.949554, 5.134079, 3.357178, 3.06395, 
    2.918762, 2.79332, 2.654312, 2.700027, 2.771515,
  2.548004, 2.169281, 1.999054, 2.074051, 2.283035, 2.493973, 2.694962, 
    2.857391, 3.063644, 3.082916, 3.187729, 3.314865, 3.476532, 3.72998, 
    3.942673, 3.926529, 3.743073, 3.42244, 3.058044, 3.17366, 3.32132, 
    2.984344, 2.672226, 2.55864, 2.847229, 3.291046, 3.331161, 3.271835, 
    3.369186, 3.563507, 3.671585, 3.617294, 3.474518, 3.383499, 3.371902, 
    3.37236, 3.322952, 3.109863, 2.901138, 2.757126, 2.589294, 2.419556, 
    2.410583, 2.517715, 2.685501, 2.715057, 2.787323, 2.805283, 2.646698, 
    2.203659, 1.859116, 1.751373, 1.848694, 2.139832, 2.498962, 2.839325, 
    3.03183, 3.198364, 3.442841, 3.713531, 4.019226, 4.351044, 4.440887, 
    4.395691, 4.27832, 4.121216, 4.003448, 3.945709, 3.790039, 3.55838, 
    4.381332, 5.073257, 4.953262, 4.685242, 4.331451, 3.769226, 4.941422, 
    4.710037, 4.47052, 4.25769, 4.351837, 4.355362, 4.495529, 4.715775, 
    4.824829, 5.03627, 5.31395, 5.496445, 5.585434, 5.613235, 5.404327, 
    4.109009, 3.856064, 3.661407, 3.444153, 3.034714,
  10.22592, 7.40567, 6.131653, 5.026382, 4.154449, 3.568039, 3.315506, 
    3.50119, 3.526123, 3.596512, 3.816879, 3.475082, 3.129639, 3.098648, 
    3.000732, 2.867554, 2.582581, 2.171265, 1.875412, 2.019745, 2.124435, 
    2.078598, 1.967911, 1.911865, 1.860107, 1.787903, 1.731979, 1.714859, 
    1.820786, 2.029312, 2.228455, 2.428085, 2.59436, 2.823868, 3.019638, 
    3.066559, 2.89325, 2.673065, 2.599228, 2.603912, 2.690002, 2.749298, 
    2.934586, 3.020065, 3.404572, 3.512726, 2.978973, 1.912354, 0.6010437, 
    -0.2281189, -0.6670532, -0.7674561, -0.6877136, -0.5030518, -0.18927, 
    0.1684265, 0.5519104, 0.9281311, 1.38562, 2.038879, 2.710815, 3.342194, 
    3.770569, 3.981659, 3.952606, 3.837555, 3.712708, 3.584839, 3.711548, 
    4.326172, 5.294464, 6.375702, 6.41217, 6.348541, 6.10495, 5.641907, 
    5.190369, 5.010529, 5.159637, 5.243759, 5.226379, 5.300201, 5.440109, 
    5.659256, 5.8909, 6.228073, 6.633606, 6.941879, 7.20285, 7.637497, 
    8.426224, 9.516724, 10.76431, 11.7843, 12.10854, 11.71199,
  9.918823, 9.868164, 9.753448, 9.734589, 9.591644, 9.213531, 8.695038, 
    8.229797, 7.867523, 7.67984, 7.650513, 7.655121, 7.677795, 7.964478, 
    8.439514, 9.030853, 9.206879, 8.887177, 8.429962, 8.038269, 7.762543, 
    7.172394, 6.370453, 5.681946, 4.829254, 3.713989, 2.788513, 2.163544, 
    1.525848, 1.17923, 1.08316, 1.475525, 2.309326, 3.204773, 3.910248, 
    4.532043, 6.261505, 4.204681, 3.317841, 3.491394, 3.916473, 3.705017, 
    3.091339, 2.25061, 1.775391, 0.9458313, 0.3729858, 0.01022339, -0.238739, 
    -0.3516846, -0.3050232, -0.2137451, -0.1629639, -0.1559448, -0.1459656, 
    -0.1081848, -0.0003967285, 0.1498718, 0.3263245, 0.5178528, 0.7279663, 
    0.940155, 1.137573, 1.320038, 1.463745, 1.546875, 1.581421, 1.601257, 
    1.6362, 1.734497, 1.899231, 2.09433, 2.214905, 2.271362, 2.23938, 
    2.11087, 1.958557, 1.930206, 2.371796, 4.318085, 5.895111, 5.882141, 
    6.004578, 6.26828, 6.474091, 6.685272, 7.233917, 7.698242, 7.98996, 
    8.2146, 8.454224, 8.789246, 9.17746, 9.571106, 9.721619, 9.845306,
  2.421234, 2.356384, 2.308014, 2.306854, 2.275635, 2.213531, 2.181061, 
    2.160339, 2.120056, 2.064087, 2.029907, 2.021362, 2.044769, 2.11496, 
    2.247314, 2.379944, 2.4711, 2.466125, 2.370972, 2.207367, 2.049988, 
    1.870789, 1.658386, 1.445313, 1.278198, 1.143799, 0.9215088, 0.6842957, 
    0.5109253, 0.4283142, 0.4024658, 0.3965454, 0.4283142, 0.565033, 
    0.7928162, 0.9947205, 1.103638, 1.10083, 1.101898, 1.190613, 1.364441, 
    1.436829, 1.355865, 1.229309, 1.068115, 0.7727966, 0.3113098, 
    -0.08724976, -0.2617188, -0.2941589, -0.2808533, -0.2905579, -0.3424988, 
    -0.3601379, -0.3178406, -0.2103577, -0.06484985, 0.07241821, 0.1690063, 
    0.2544861, 0.3853455, 0.5687561, 0.7503967, 0.8957825, 1.077606, 
    1.270569, 1.46698, 1.627258, 1.710999, 1.745178, 1.772736, 1.841156, 
    1.907349, 1.975586, 2.04425, 2.061096, 1.965485, 1.808136, 1.703857, 
    1.819458, 2.167572, 2.328644, 2.190155, 1.823975, 1.766144, 1.922424, 
    2.179291, 2.428833, 2.654755, 2.732178, 2.713806, 2.689331, 2.697601, 
    2.647522, 2.584717, 2.518799,
  1.533966, 1.499817, 1.449432, 1.373657, 1.317749, 1.306244, 1.324432, 
    1.335999, 1.339844, 1.336456, 1.37207, 1.504364, 1.636841, 1.696045, 
    1.676819, 1.640808, 1.627472, 1.639648, 1.627075, 1.561981, 1.429443, 
    1.283203, 1.123291, 1.046295, 1.072021, 1.094604, 1.060608, 0.9909058, 
    0.924469, 0.8734436, 0.7933044, 0.6654358, 0.5419312, 0.4615173, 
    0.4230347, 0.4210815, 0.4829407, 0.6013489, 0.7591553, 0.940155, 
    1.100403, 1.239716, 1.375763, 1.395508, 1.308411, 1.202209, 0.9975891, 
    0.664917, 0.2876892, -0.01556396, -0.1434326, -0.2064514, -0.2541199, 
    -0.298645, -0.2966614, -0.2373047, -0.107605, 0.07305908, 0.2085266, 
    0.2823486, 0.3964844, 0.5423279, 0.6791687, 0.8017578, 1.008545, 
    1.296814, 1.501831, 1.593903, 1.654419, 1.73822, 1.839783, 1.9263, 
    1.959808, 2.00473, 2.021423, 1.959106, 1.807922, 1.744995, 1.731781, 
    1.736389, 1.793091, 1.868042, 1.787994, 1.448578, 1.304169, 1.254303, 
    1.312439, 1.397003, 1.469482, 1.490143, 1.532684, 1.574158, 1.599213, 
    1.621613, 1.603455, 1.562073,
  1.363403, 1.480316, 1.595825, 1.646545, 1.630524, 1.592316, 1.56308, 
    1.560028, 1.584961, 1.590118, 1.602417, 1.675903, 1.739166, 1.757355, 
    1.836517, 1.982971, 2.171417, 2.277679, 2.194916, 1.929565, 1.722839, 
    1.60965, 1.47879, 1.3685, 1.332031, 1.356323, 1.425934, 1.467896, 
    1.44577, 1.358704, 1.207825, 1.016022, 0.8884888, 0.8519287, 0.8417358, 
    0.8167725, 0.8305359, 0.9263611, 1.088409, 1.227295, 1.34491, 1.45813, 
    1.513275, 1.411713, 1.306488, 1.255005, 1.132996, 0.9438171, 0.6283264, 
    0.2982178, 0.2026062, 0.2142334, 0.1886597, 0.1558533, 0.1395264, 
    0.1769714, 0.255188, 0.3762207, 0.4845276, 0.5489502, 0.6590881, 
    0.7944031, 0.8881531, 0.9835205, 1.211182, 1.44696, 1.525024, 1.537598, 
    1.611877, 1.738831, 1.831665, 1.849823, 1.872833, 1.886749, 1.804138, 
    1.604187, 1.598663, 2.152496, 2.163483, 1.61203, 1.558228, 1.646027, 
    1.706329, 1.511963, 1.240936, 1.240479, 1.440582, 1.625519, 1.687378, 
    1.650848, 1.635742, 1.60202, 1.539246, 1.483795, 1.419006, 1.349274,
  1.802094, 1.850159, 1.900848, 1.924347, 1.956055, 2.00415, 2.079346, 
    2.145111, 2.154877, 2.153046, 2.209564, 2.29126, 2.306549, 2.277466, 
    2.273132, 2.350128, 2.524353, 2.675781, 2.629944, 2.463745, 2.434296, 
    2.49054, 2.38974, 2.172852, 2.01416, 1.961517, 1.963928, 1.942047, 
    1.870575, 1.744476, 1.580658, 1.411346, 1.322998, 1.31134, 1.281158, 
    1.215668, 1.193268, 1.237152, 1.333893, 1.503662, 1.651001, 1.689331, 
    1.65744, 1.640808, 1.672516, 1.617828, 1.447144, 1.262512, 1.031921, 
    0.8209534, 0.7734375, 0.8415527, 0.8378906, 0.7775879, 0.7741699, 
    0.8270874, 0.8622437, 0.9119568, 0.9994202, 1.072388, 1.172852, 1.289307, 
    1.346283, 1.388092, 1.521667, 1.639435, 1.657867, 1.665222, 1.748322, 
    1.841461, 1.846863, 1.811279, 1.78717, 1.737762, 1.664917, 1.572845, 
    1.845947, 2.016541, 1.75177, 1.658051, 1.508789, 1.452484, 1.441467, 
    1.259583, 1.168579, 1.438049, 1.724579, 1.867645, 1.882477, 1.875854, 
    1.918182, 1.930725, 1.900055, 1.913483, 1.924927, 1.85553,
  2.10849, 2.107788, 2.182922, 2.266602, 2.342316, 2.434296, 2.622192, 
    2.765411, 2.771271, 2.830322, 2.998596, 3.085388, 3.072571, 3.084991, 
    3.06311, 3.025818, 3.09964, 3.251373, 3.281952, 3.413513, 3.668884, 
    3.642731, 3.163147, 2.550201, 2.203339, 2.105591, 2.116974, 2.091797, 
    1.982239, 1.800568, 1.631836, 1.571289, 1.588287, 1.612579, 1.610626, 
    1.603302, 1.622528, 1.644012, 1.67572, 1.854889, 2.156708, 2.17688, 
    2.038361, 2.041138, 2.205719, 2.287628, 1.979492, 1.753998, 1.628632, 
    1.520721, 1.591919, 1.702545, 1.697632, 1.595428, 1.492981, 1.423248, 
    1.381287, 1.407043, 1.476624, 1.498962, 1.525787, 1.555145, 1.579224, 
    1.6539, 1.764496, 1.821228, 1.845428, 1.897766, 1.930298, 1.899536, 
    1.819916, 1.790497, 1.755096, 1.673615, 1.615234, 1.576813, 1.755249, 
    1.709229, 1.834412, 1.824677, 1.650116, 1.347534, 1.129761, 1.014832, 
    1.264404, 1.70755, 2.016144, 2.140106, 2.191528, 2.195892, 2.197266, 
    2.195496, 2.13736, 2.062286, 2.079926, 2.129456,
  2.508331, 2.429291, 2.405334, 2.470581, 2.646301, 3.027283, 3.503326, 
    3.700897, 3.776703, 3.953064, 4.15097, 3.993622, 3.599335, 3.342194, 
    3.224762, 3.178497, 3.207031, 3.272522, 3.367706, 3.493683, 3.4245, 
    3.010681, 2.402527, 1.944275, 1.843506, 2.040649, 2.201782, 2.167694, 
    2.065125, 2.020782, 2.01889, 2.027679, 1.999329, 1.937561, 1.933655, 
    1.954224, 1.976044, 1.983856, 1.963867, 2.249146, 2.792328, 2.856781, 
    2.605286, 2.552582, 2.712036, 2.879028, 2.88736, 2.606506, 2.559113, 
    2.576172, 2.671356, 2.555481, 2.302155, 2.080078, 1.913605, 1.81485, 
    1.797272, 1.842194, 1.899261, 1.884766, 1.851227, 1.87265, 1.896698, 
    1.945313, 1.96933, 1.980255, 2.015045, 2.030457, 1.996643, 1.959625, 
    1.923767, 1.865479, 1.773376, 1.659729, 1.600006, 1.51355, 1.552979, 
    1.37326, 1.635712, 1.858643, 1.721252, 1.651489, 1.689056, 1.835083, 
    1.955414, 2.098297, 2.253204, 2.295685, 2.334045, 2.347443, 2.326996, 
    2.365356, 2.363953, 2.36496, 2.476898, 2.559174,
  2.391998, 2.299744, 2.291931, 2.507874, 2.848572, 3.163757, 3.298828, 
    3.631897, 3.571625, 3.236908, 2.789764, 2.397125, 2.110687, 1.974945, 
    1.983582, 2.183258, 2.476715, 2.682556, 2.687439, 2.529053, 2.385223, 
    2.261963, 2.159454, 2.166016, 2.272522, 2.379303, 2.401794, 2.339966, 
    2.361786, 2.434326, 2.27356, 2.160095, 2.066925, 1.964966, 2.124664, 
    2.230804, 2.125793, 2.215302, 2.373627, 2.502655, 2.860229, 3.237823, 
    3.293427, 3.025299, 2.945831, 3.044189, 3.069214, 2.870422, 2.657166, 
    2.521759, 2.365173, 2.351379, 2.291992, 2.22168, 2.149567, 2.1138, 
    2.099152, 2.074982, 2.074219, 2.061066, 2.069122, 2.099731, 2.11203, 
    2.12558, 2.130737, 2.144012, 2.206055, 2.194214, 2.124603, 2.076233, 
    2.023834, 1.926941, 1.759949, 1.572968, 1.43692, 1.240967, 1.157959, 
    1.502014, 1.689667, 1.340088, 1.57077, 1.844482, 2.21524, 2.410736, 
    2.285614, 2.180725, 2.273285, 2.33432, 2.384308, 2.410553, 2.419159, 
    2.452484, 2.407684, 2.3508, 2.385101, 2.412384,
  2.214661, 2.054749, 2.001373, 2.059448, 2.094879, 2.203461, 2.364563, 
    2.269073, 2.149475, 2.127411, 1.478058, 1.595642, 1.705536, 1.78653, 
    1.855011, 2.004456, 2.149323, 2.203491, 2.186523, 2.109833, 2.174225, 
    2.284698, 2.321625, 2.411194, 2.409454, 2.364136, 2.339325, 2.32605, 
    2.389526, 2.184662, 1.831329, 1.820618, 1.79184, 1.793365, 1.943695, 
    1.945374, 1.883392, 2.285095, 2.867004, 2.924561, 2.676514, 2.88913, 
    3.457275, 3.268158, 3.002472, 3.018097, 2.868378, 2.566467, 2.228119, 
    1.952759, 2.032684, 2.178131, 2.257629, 2.290192, 2.29184, 2.26712, 
    2.22995, 2.150177, 2.14975, 2.155212, 2.197601, 2.266602, 2.243866, 
    2.23053, 2.22345, 2.172913, 2.142456, 2.065613, 1.973755, 1.870941, 
    1.72467, 1.54895, 1.379761, 1.2453, 1.09024, 0.910553, 0.9950562, 
    2.417664, 2.306641, 1.549225, 1.859497, 2.621826, 2.402161, 2.438202, 
    2.269318, 2.1026, 2.154358, 2.229309, 2.33313, 2.376373, 2.3927, 
    2.398315, 2.340515, 2.343567, 2.338928, 2.295898,
  1.698608, 1.628479, 1.61792, 1.679108, 1.780273, 3.355591, 3.627289, 
    3.583771, 3.311584, 2.051361, 1.97702, 2.135895, 2.183533, 2.17691, 
    2.145447, 2.256439, 2.408203, 2.427734, 2.430267, 2.444489, 2.508453, 
    2.525146, 2.463135, 2.439789, 2.364563, 2.262299, 2.203522, 2.108826, 
    1.971558, 1.746674, 1.780121, 2.602142, 2.484711, 2.423096, 2.809509, 
    2.952423, 2.916687, 3.215027, 3.518555, 3.454559, 3.03653, 2.596802, 
    2.320129, 2.24765, 2.340027, 2.354889, 2.210022, 1.959442, 1.940155, 
    2.134552, 2.319855, 2.442322, 2.456329, 2.373505, 2.317505, 2.266022, 
    2.195129, 2.090637, 2.072083, 2.10202, 2.121216, 2.17514, 2.139709, 
    2.121277, 2.079559, 1.979614, 1.906586, 1.747131, 1.618744, 1.442383, 
    1.241089, 1.115601, 0.9574585, 0.8867798, 0.7252808, 0.7691956, 1.233765, 
    2.417755, 3.134399, 2.306396, 2.436249, 3.088287, 2.955322, 2.410858, 
    2.300598, 2.226898, 2.301758, 2.403717, 2.436646, 2.389709, 2.347534, 
    2.263214, 2.161499, 2.084625, 1.992767, 1.852081,
  1.424927, 1.460602, 1.650665, 1.86142, 2.410278, 3.996246, 4.212891, 
    3.929932, 3.178009, 2.084564, 2.049408, 2.238556, 2.262451, 2.279694, 
    2.336578, 2.544861, 2.697998, 2.66626, 2.607025, 2.488495, 2.443359, 
    2.372925, 2.260437, 2.136902, 2.02359, 1.949097, 1.888397, 1.872589, 
    1.974792, 2.006714, 2.336365, 3.458679, 3.060455, 3.289124, 3.733917, 
    3.540283, 3.737305, 3.743042, 3.802032, 3.952972, 3.58963, 2.251434, 
    1.894073, 2.025787, 2.20639, 2.307159, 2.329773, 2.299042, 2.351227, 
    2.46875, 2.443695, 2.441864, 2.401886, 2.302856, 2.198608, 2.184631, 
    2.082245, 2.026123, 2.007416, 2.034973, 2.017059, 1.960327, 1.903717, 
    1.81485, 1.699341, 1.537201, 1.463531, 1.290222, 1.176575, 1.053894, 
    0.9225159, 0.910553, 0.8309937, 0.825531, 0.7302551, 1.115814, 1.889954, 
    2.895172, 4.063599, 3.049805, 3.104034, 3.571106, 3.417725, 3.229279, 
    2.418823, 2.229034, 2.243317, 2.316345, 2.275024, 2.224792, 2.166412, 
    2.054749, 1.94101, 1.773743, 1.634399, 1.463867,
  1.649689, 1.851105, 2.161072, 2.634766, 3.980316, 4.225372, 4.152161, 
    4.575989, 4.089386, 3.472015, 2.110565, 2.179749, 2.48114, 2.320496, 
    2.436188, 2.514496, 2.495575, 2.420135, 2.38736, 2.291229, 2.21582, 
    2.110229, 1.996429, 1.967896, 1.946289, 1.945496, 1.997864, 2.163544, 
    2.293884, 2.360809, 2.5961, 3.540833, 3.7789, 3.99231, 4.061279, 
    3.664856, 3.76236, 3.722595, 3.726227, 3.760559, 3.588867, 2.209839, 
    2.278534, 2.432892, 2.422607, 2.411957, 2.401306, 2.355652, 2.317596, 
    2.326904, 2.347412, 2.354889, 2.312866, 2.261383, 2.210602, 2.16333, 
    2.079559, 2.029755, 1.992523, 1.977753, 1.895966, 1.808594, 1.722076, 
    1.563751, 1.46991, 1.285675, 1.133484, 1.076477, 1.008209, 0.9555359, 
    0.9499207, 0.8963623, 0.8756409, 0.9279785, 1.050354, 1.556183, 2.228851, 
    3.606689, 4.370728, 3.405212, 3.625183, 3.924103, 4.16098, 3.214844, 
    2.931824, 2.280792, 2.119659, 2.166077, 2.061157, 1.976685, 1.848053, 
    1.715607, 1.637756, 1.542175, 1.525665, 1.519958,
  2.044403, 2.243866, 2.395966, 2.569397, 3.674988, 3.23822, 3.483002, 
    4.13678, 3.655853, 3.554352, 2.098511, 2.114777, 2.805084, 2.686066, 
    2.329285, 2.281372, 2.273102, 2.239044, 2.223572, 2.177277, 2.124542, 
    2.093903, 2.074799, 2.1026, 2.133667, 2.205994, 2.338867, 2.4664, 
    2.492706, 2.520508, 2.596344, 2.896149, 4.098114, 4.498108, 4.091003, 
    3.762238, 3.934753, 3.974274, 3.96756, 3.381897, 2.353638, 2.291321, 
    2.452026, 2.517914, 2.433258, 2.412109, 2.347473, 2.325195, 2.285339, 
    2.262451, 2.28125, 2.233734, 2.211456, 2.212128, 2.232422, 2.204803, 
    2.157806, 2.083527, 2.033661, 1.944183, 1.872131, 1.778076, 1.688202, 
    1.509216, 1.395111, 1.299011, 1.243683, 1.199554, 1.18158, 1.198822, 
    1.171875, 1.207397, 1.248657, 1.389069, 1.544006, 1.819519, 2.332092, 
    3.964905, 4.290466, 3.328918, 3.045959, 3.665405, 4.123352, 3.405334, 
    3.172272, 3.117554, 2.074738, 2.053711, 1.968689, 1.889343, 1.795074, 
    1.77066, 1.757263, 1.75592, 1.866486, 1.934753,
  2.45462, 2.570892, 2.489258, 2.396484, 4.270325, 4.512421, 4.3013, 
    4.246429, 3.778931, 3.296417, 2.720123, 2.274048, 2.597534, 2.685608, 
    2.349091, 2.1427, 2.15271, 2.22052, 2.238586, 2.246857, 2.268433, 
    2.249329, 2.228516, 2.274414, 2.362061, 2.421509, 2.493011, 2.538391, 
    2.528564, 2.46225, 2.478271, 2.556427, 2.747284, 3.57486, 3.147461, 
    3.031769, 3.436127, 2.725861, 3.03067, 2.372406, 2.313812, 2.46756, 
    2.528107, 2.501282, 2.422272, 2.371552, 2.295441, 2.280121, 2.225403, 
    2.240814, 2.237091, 2.18399, 2.125214, 2.159058, 2.189301, 2.153412, 
    2.114899, 2.027008, 1.975647, 1.91626, 1.871674, 1.778534, 1.764038, 
    1.69278, 1.63028, 1.600342, 1.595825, 1.634613, 1.636414, 1.652679, 
    1.639984, 1.691467, 1.709961, 1.783539, 1.976685, 2.2901, 3.884705, 
    4.321564, 3.45166, 3.330017, 3.22937, 3.462646, 3.558075, 3.270966, 
    3.592834, 3.010986, 2.081848, 2.095184, 2.067627, 2.022919, 2.008911, 
    2.074097, 2.14389, 2.212646, 2.300079, 2.382996,
  2.632019, 2.612427, 2.486694, 2.327332, 3.101105, 3.916687, 3.712555, 
    3.774078, 3.762115, 3.358124, 3.132751, 2.355591, 2.395905, 2.475861, 
    2.25766, 2.111084, 2.102417, 2.235229, 2.258331, 2.242706, 2.267273, 
    2.292389, 2.3461, 2.423126, 2.494659, 2.50174, 2.576691, 2.568359, 
    2.51236, 2.408417, 2.419006, 2.406952, 2.271362, 2.24176, 2.404297, 
    2.650452, 3.007263, 2.318298, 2.533417, 2.159332, 2.228241, 2.469147, 
    2.436676, 2.391541, 2.277527, 2.189301, 2.117981, 2.11676, 2.122467, 
    2.162903, 2.151245, 2.066467, 1.955261, 2.012115, 2.077454, 2.124359, 
    2.149292, 2.081421, 2.068298, 2.082092, 2.052032, 2.049866, 2.061798, 
    2.03009, 1.987213, 2.018097, 2.025635, 2.049225, 2.067902, 2.137634, 
    2.186859, 2.226837, 2.204559, 2.266724, 2.515778, 2.981628, 3.149475, 
    3.125702, 3.361145, 3.379303, 3.243042, 3.59256, 3.505066, 3.248108, 
    3.338806, 2.719849, 2.103638, 2.159546, 2.193542, 2.208801, 2.263153, 
    2.345764, 2.434052, 2.511536, 2.550842, 2.615875,
  2.567505, 2.529114, 2.437897, 2.34494, 2.90976, 3.012421, 2.928894, 
    2.537292, 2.715759, 2.815125, 2.872894, 2.282623, 2.418671, 2.446106, 
    2.273285, 2.226257, 2.237305, 2.377167, 2.467834, 2.492706, 2.478912, 
    2.508728, 2.541077, 2.552673, 2.607819, 2.635681, 2.581635, 2.415436, 
    2.339203, 2.439514, 2.431519, 2.453949, 2.508972, 2.462158, 2.378448, 
    2.402344, 2.270966, 2.242706, 2.53595, 2.107483, 2.192322, 2.292389, 
    2.292694, 2.299011, 2.141785, 1.997375, 1.938293, 1.993286, 2.054871, 
    2.060303, 2.089386, 2.050964, 2.003387, 2.005768, 2.067627, 2.119324, 
    2.115936, 2.1091, 2.124359, 2.154724, 2.10788, 2.123718, 2.1362, 
    2.141602, 2.128235, 2.174072, 2.209351, 2.240997, 2.317078, 2.426239, 
    2.477203, 2.491852, 2.533417, 2.595001, 2.525635, 2.874207, 3.292694, 
    3.574402, 3.574677, 2.98941, 3.064911, 3.326874, 3.201172, 3.156067, 
    3.224548, 2.885315, 2.948761, 2.253723, 2.275269, 2.272247, 2.315155, 
    2.364197, 2.449799, 2.52597, 2.579041, 2.592377,
  2.350189, 2.33139, 2.199738, 2.487762, 3.340942, 2.928131, 2.798309, 
    2.418884, 2.1539, 1.868408, 2.192322, 2.257202, 2.264801, 2.340912, 
    2.371613, 2.374756, 2.393158, 2.526306, 2.572632, 2.597321, 2.572144, 
    2.619568, 2.629364, 2.673462, 2.683716, 2.648254, 2.452667, 2.293732, 
    2.478577, 2.399414, 2.334076, 2.232056, 2.364075, 2.41452, 2.369354, 
    2.385742, 2.173218, 2.601349, 2.725067, 2.548126, 2.201691, 2.180359, 
    2.19754, 2.212219, 2.130981, 2.075836, 2.078247, 2.096436, 2.160767, 
    2.152466, 2.139587, 2.146027, 2.151947, 2.152863, 2.124084, 2.175537, 
    2.173645, 2.162781, 2.139648, 2.158264, 2.151306, 2.136963, 2.128571, 
    2.15567, 2.197083, 2.236481, 2.284576, 2.333405, 2.417145, 2.445374, 
    2.456512, 2.430939, 2.42337, 2.481842, 2.42688, 3.129944, 3.63208, 
    3.272339, 3.041077, 2.759338, 3.033142, 2.966095, 2.880341, 2.858459, 
    2.981812, 2.698303, 2.641388, 2.263336, 2.316467, 2.317383, 2.392242, 
    2.39917, 2.430267, 2.423004, 2.446228, 2.402069,
  2.242188, 2.296722, 2.369476, 3.657043, 3.87207, 2.939209, 2.907623, 
    2.726959, 2.3815, 1.617065, 1.724152, 2.595093, 2.401062, 2.449219, 
    2.436829, 2.487976, 2.546021, 2.549469, 2.565643, 2.588287, 2.586731, 
    2.589447, 2.542297, 2.542664, 2.441223, 2.378784, 2.267273, 2.623962, 
    2.56778, 2.368042, 2.739105, 2.416748, 2.626282, 2.248871, 2.295563, 
    2.673309, 2.58197, 2.266479, 2.379944, 2.071442, 2.03891, 2.02356, 
    2.009491, 2.035431, 2.006775, 1.930603, 1.865692, 1.892456, 1.942017, 
    1.957031, 1.929321, 1.953644, 1.996368, 2.041565, 2.085541, 2.146149, 
    2.198883, 2.249939, 2.286316, 2.335083, 2.348511, 2.358521, 2.395691, 
    2.428711, 2.488525, 2.509125, 2.527802, 2.554565, 2.519409, 2.432831, 
    2.399658, 2.326111, 2.216736, 2.179047, 2.174408, 2.826569, 3.082733, 
    2.980988, 3.03952, 2.936127, 3.106384, 3.771088, 3.248169, 2.802551, 
    2.767731, 2.197906, 2.167969, 2.297455, 2.388794, 2.407104, 2.439911, 
    2.392426, 2.423065, 2.40274, 2.376617, 2.320892,
  2.236023, 2.319061, 2.400391, 3.040955, 3.064178, 2.843872, 3.020691, 
    2.780487, 2.697327, 1.985535, 1.952728, 3.350342, 3.222534, 2.484894, 
    2.435242, 2.57312, 2.547668, 2.498627, 2.507111, 2.461121, 2.455353, 
    2.433075, 2.458527, 2.499176, 2.411591, 2.24408, 2.146088, 2.568756, 
    2.191284, 2.330872, 2.475403, 2.435272, 2.761993, 2.214996, 2.143555, 
    2.124146, 1.987732, 1.943359, 2.017456, 2.109955, 2.005859, 1.9552, 
    1.985138, 1.97702, 1.919922, 1.854889, 1.834717, 1.854645, 1.86795, 
    1.907928, 1.919464, 1.942017, 1.97641, 2.011444, 2.04425, 2.091339, 
    2.161865, 2.223694, 2.279358, 2.336853, 2.400909, 2.427582, 2.465118, 
    2.535736, 2.601501, 2.642456, 2.701447, 2.684448, 2.607758, 2.479248, 
    2.340027, 2.27179, 2.195313, 2.089844, 1.975769, 2.706848, 2.920837, 
    2.697449, 2.878754, 3.239899, 3.286316, 3.456512, 3.125458, 2.113159, 
    2.060364, 2.085266, 2.184845, 2.273224, 2.366089, 2.409637, 2.379883, 
    2.390411, 2.413879, 2.382355, 2.353363, 2.327606,
  2.957031, 2.527588, 2.715576, 3.05307, 3.076294, 2.992767, 2.956238, 
    2.916077, 2.953918, 1.99826, 2.213074, 3.161865, 3.120239, 2.589142, 
    2.630646, 2.687714, 2.683716, 2.653839, 2.611481, 2.620575, 2.607208, 
    2.547333, 2.535919, 2.585938, 2.560272, 2.281586, 2.634888, 3.129028, 
    2.057037, 2.169281, 2.182556, 2.865631, 2.193817, 2.25177, 2.133453, 
    2.147461, 2.129425, 2.192139, 2.243439, 2.222076, 2.171356, 2.143829, 
    2.138153, 2.150909, 2.152527, 2.158081, 2.172394, 2.182678, 2.204163, 
    2.203766, 2.211334, 2.205231, 2.208832, 2.203186, 2.188995, 2.179474, 
    2.173004, 2.148865, 2.131592, 2.103912, 2.137085, 2.157471, 2.189301, 
    2.23288, 2.255066, 2.3591, 2.470978, 2.533997, 2.502289, 2.396057, 
    2.338776, 2.365234, 2.308411, 2.093689, 2.017242, 2.826416, 2.904419, 
    3.180786, 3.361206, 3.7966, 3.336914, 2.881165, 2.460938, 1.998108, 
    2.059174, 2.076569, 2.1651, 2.207886, 2.31601, 2.36319, 2.38504, 
    2.390564, 2.314697, 2.373047, 2.711395, 2.982574,
  3.115814, 2.947083, 3.212738, 3.973053, 4.329376, 4.104645, 3.685669, 
    3.920166, 4.121216, 3.526367, 3.642761, 4.022339, 4.138397, 3.649414, 
    2.585358, 2.702789, 2.902954, 2.828705, 2.84494, 2.806305, 2.589783, 
    2.472412, 2.486511, 2.453247, 2.391357, 2.179291, 2.386536, 3.299286, 
    2.100922, 2.212372, 2.064911, 2.0224, 2.193604, 3.035858, 2.227264, 
    2.239563, 2.293823, 2.309448, 2.328918, 2.328644, 2.333466, 2.351685, 
    2.356903, 2.353363, 2.375244, 2.394653, 2.450439, 2.439667, 2.455231, 
    2.458801, 2.470978, 2.465759, 2.462036, 2.464264, 2.462219, 2.448761, 
    2.410034, 2.348938, 2.27951, 2.217773, 2.17804, 2.145325, 2.147125, 
    2.161469, 2.201447, 2.289063, 2.400238, 2.534241, 2.51825, 2.496826, 
    2.512299, 2.509247, 2.593628, 2.616608, 2.736237, 2.868958, 3.224274, 
    3.383881, 3.246246, 2.984833, 2.299927, 2.386292, 2.265228, 2.061188, 
    2.059479, 2.067566, 2.123505, 2.189056, 2.237457, 2.321167, 2.354828, 
    2.220367, 2.241882, 3.165955, 3.043121, 2.948975,
  3.838562, 3.797089, 3.746948, 3.913147, 4.18158, 4.586975, 4.488434, 
    4.184631, 4.178192, 4.642639, 4.714722, 4.445374, 4.652344, 3.935608, 
    2.560608, 2.499817, 2.769012, 2.844391, 2.973785, 2.902069, 3.267822, 
    3.208466, 2.611328, 2.585419, 2.437958, 2.303253, 2.392242, 2.025848, 
    2.570465, 3.365387, 2.150208, 2.054291, 2.158783, 3.030457, 2.209351, 
    2.268738, 2.272858, 2.325073, 2.364899, 2.358643, 2.372192, 2.367645, 
    2.37851, 2.384827, 2.441071, 2.446228, 2.499664, 2.503967, 2.531372, 
    2.557922, 2.57251, 2.558594, 2.566132, 2.562897, 2.541412, 2.510345, 
    2.447205, 2.366211, 2.30188, 2.222717, 2.166077, 2.16217, 2.177094, 
    2.200714, 2.210297, 2.204559, 2.257477, 2.361908, 2.443939, 2.528137, 
    2.409454, 2.581055, 3.394745, 2.934113, 2.48999, 2.639648, 2.595642, 
    2.449951, 2.34375, 2.272003, 2.183258, 2.238525, 2.14978, 2.104492, 
    2.051117, 2.088348, 2.113647, 2.200989, 2.225311, 2.348969, 2.379883, 
    2.453949, 3.881653, 4.453461, 4.343048, 3.958344,
  4.743683, 4.584045, 4.114441, 3.682556, 3.284576, 3.130554, 3.129242, 
    2.945038, 3.263733, 3.576233, 3.901825, 4.687714, 4.553955, 4.062744, 
    3.567383, 2.635895, 2.545166, 2.646423, 2.827545, 2.753571, 3.760223, 
    4.1474, 2.590759, 2.596283, 2.600586, 2.569031, 2.631042, 1.722534, 
    1.309265, 1.861389, 1.903778, 1.992126, 1.890686, 2.003967, 2.118164, 
    2.228516, 2.245239, 2.256042, 2.278076, 2.280273, 2.288483, 2.250671, 
    2.269409, 2.21756, 2.2276, 2.255157, 2.283844, 2.292511, 2.345581, 
    2.421722, 2.459503, 2.468628, 2.468109, 2.464203, 2.461273, 2.43338, 
    2.352722, 2.268036, 2.190552, 2.071411, 2.035675, 2.042847, 2.09726, 
    2.129608, 2.108917, 2.000122, 1.853638, 1.97052, 2.517578, 4.198425, 
    3.299591, 4.27066, 4.6362, 2.206146, 2.411865, 2.433136, 2.352142, 
    2.310425, 2.207092, 2.187714, 2.155731, 2.095642, 2.023102, 2.000305, 
    1.984558, 2.002472, 1.994598, 2.051544, 2.049438, 2.225342, 2.392639, 
    2.84375, 4.598907, 4.886963, 4.855865, 4.782623,
  4.604095, 4.419342, 4.098969, 3.906982, 3.433319, 3.361084, 3.176697, 
    3.16861, 3.395569, 3.18045, 2.324493, 4.515778, 4.839081, 4.479431, 
    4.692963, 4.217712, 2.667328, 2.583801, 2.936981, 2.843872, 3.791931, 
    4.283997, 3.510468, 2.891815, 2.439636, 2.237183, 2.868774, 2.209839, 
    1.017059, 1.427032, 1.82077, 2.074219, 1.888367, 1.912384, 1.918732, 
    2.012177, 2.079498, 2.082733, 2.10907, 2.124298, 2.122406, 2.061401, 
    2.083313, 2.028473, 1.99765, 1.998718, 1.994263, 2.024933, 2.078857, 
    2.12027, 2.1745, 2.21051, 2.249329, 2.286194, 2.295776, 2.251373, 
    2.172668, 2.081848, 1.959259, 1.834442, 1.763092, 1.69455, 1.72644, 
    1.811218, 1.862366, 1.651733, 1.489258, 2.107941, 4.570129, 4.418732, 
    3.38205, 4.113647, 4.097778, 2.099426, 2.226227, 2.203766, 2.196686, 
    2.190887, 2.115234, 2.122925, 2.100342, 2.025909, 1.965088, 1.890686, 
    1.801758, 1.798065, 1.807678, 1.812805, 1.763794, 1.857239, 2.038086, 
    2.692505, 4.522186, 4.854034, 4.766663, 4.764709,
  4.564636, 4.59201, 4.373627, 4.147095, 3.721497, 3.555603, 3.561859, 
    3.471222, 3.543243, 3.672729, 2.420013, 4.782684, 4.949921, 4.799591, 
    5.404968, 4.860291, 3.087677, 3.019989, 4.248962, 4.23288, 4.109619, 
    3.88678, 3.563171, 3.735687, 3.237366, 2.346954, 3.084778, 2.257172, 
    1.439392, 1.041138, 1.414825, 2.028198, 1.854156, 1.772644, 1.736572, 
    1.878326, 2.011475, 2.015503, 2.016449, 2.0354, 2.061005, 2.089905, 
    2.006104, 1.945648, 1.854767, 1.765472, 1.731201, 1.730743, 1.794128, 
    1.878387, 1.974426, 2.010345, 2.078186, 2.123169, 2.131378, 2.136047, 
    2.10434, 2.042755, 1.955414, 1.832275, 1.732666, 1.673126, 1.729156, 
    1.788879, 1.801758, 1.626709, 1.893158, 3.954346, 5.03952, 4.531586, 
    3.480133, 2.497467, 2.235291, 2.121277, 2.177826, 2.050385, 2.041656, 
    2.110413, 2.291687, 2.310181, 2.278198, 2.263031, 2.207855, 2.111115, 
    2.033203, 1.983124, 1.957428, 1.922211, 1.833588, 1.83429, 1.862946, 
    2.298615, 4.074738, 4.557617, 4.452148, 4.408539,
  3.960358, 4.158325, 4.082153, 4.031769, 3.783539, 3.503723, 3.703827, 
    3.644928, 3.646667, 4.031494, 4.139923, 4.251678, 4.631317, 5.374084, 
    5.539368, 5.346619, 5.33139, 5.6026, 5.402222, 5.063538, 4.411011, 
    4.035797, 3.735931, 5.078491, 5.968109, 3.448456, 2.914795, 1.88385, 
    1.842499, 1.700897, 1.681824, 1.811401, 1.982941, 1.85733, 1.891205, 
    1.953339, 2.002197, 2.039642, 2.119385, 2.156128, 2.1539, 2.144989, 
    2.089233, 1.968018, 1.853638, 1.760864, 1.717712, 1.65976, 1.656128, 
    1.732239, 1.798431, 1.854034, 1.950134, 1.972321, 1.989655, 2.050385, 
    1.997925, 1.943817, 1.871277, 1.816528, 1.747192, 1.679352, 1.7276, 
    1.761993, 1.726379, 1.914063, 2.714539, 3.210358, 3.950592, 3.942078, 
    3.632477, 2.568634, 2.42688, 2.540833, 2.752228, 2.074921, 1.992004, 
    2.010284, 2.11203, 2.15976, 2.234131, 2.31958, 2.340302, 2.338806, 
    2.316193, 2.300781, 2.241943, 2.19693, 2.101685, 1.999084, 1.838409, 
    1.814819, 2.429291, 4.013275, 4.419098, 4.033936,
  4.152222, 4.188538, 3.911133, 3.672241, 3.36792, 2.552673, 3.309174, 
    3.500702, 2.682343, 3.793549, 4.335815, 4.290253, 4.446838, 5.122131, 
    5.401306, 4.998962, 5.111786, 5.541534, 5.050598, 5.537994, 4.924011, 
    4.682739, 5.157867, 2.941742, 2.754211, 4.128296, 3.08847, 3.067688, 
    3.082855, 3.648621, 3.293243, 2.792084, 2.459778, 1.625397, 1.976868, 
    2.144318, 2.076416, 2.133087, 2.161194, 2.176544, 2.18811, 2.140106, 
    2.112762, 2.062561, 1.973236, 1.907288, 1.847412, 1.798584, 1.753632, 
    1.741272, 1.81311, 1.885925, 1.939392, 1.980621, 1.987305, 1.954865, 
    1.881836, 1.841278, 1.797699, 1.766205, 1.74588, 1.636597, 1.643158, 
    1.714508, 1.827148, 2.644958, 2.856903, 3.376953, 3.775635, 3.812714, 
    3.571136, 3.074829, 2.953827, 2.919922, 2.736176, 2.121552, 1.972809, 
    1.963867, 2.02005, 1.980682, 1.949036, 1.909973, 1.950867, 2.039642, 
    2.095428, 2.163483, 2.205078, 2.209961, 2.220703, 2.190948, 2.115875, 
    1.923706, 1.926239, 2.508331, 4.599609, 4.729431,
  4.596466, 4.797119, 4.401825, 2.763855, 2.46817, 2.34082, 2.35379, 
    2.392334, 2.624207, 2.912384, 4.425781, 4.869659, 5.393951, 4.866364, 
    4.653625, 4.648621, 4.704376, 4.39566, 4.312836, 6.03717, 5.643036, 
    5.630035, 4.938232, 3.135345, 3.806183, 2.354156, 2.378784, 2.168549, 
    2.537903, 3.379364, 3.965363, 3.242432, 2.682861, 1.751373, 2.733582, 
    2.414063, 2.658783, 2.838837, 2.335419, 2.289368, 2.27005, 2.215149, 
    2.180847, 2.135437, 2.086334, 2.083099, 2.078918, 2.048706, 1.992584, 
    1.928833, 1.93808, 1.966888, 1.970184, 1.962891, 1.947968, 1.915131, 
    1.892578, 1.822601, 1.705353, 1.654877, 1.652008, 1.630188, 1.668701, 
    1.659882, 1.719452, 2.233276, 2.90451, 3.842407, 4.50412, 4.095642, 
    3.572021, 3.120972, 3.117889, 3.133942, 3.074005, 2.980927, 2.375854, 
    2.069092, 1.926239, 1.930023, 2.016937, 1.98764, 1.804352, 1.651184, 
    1.512604, 1.512756, 1.618103, 1.668488, 1.724304, 1.90918, 2.094513, 
    2.017365, 1.809052, 1.849335, 2.356506, 4.307617,
  3.364777, 2.344604, 2.284302, 2.243988, 2.234619, 2.262634, 2.722137, 
    2.741394, 2.820679, 3.140961, 3.214539, 4.04837, 4.132294, 3.199768, 
    2.620056, 3.855774, 4.197449, 3.885559, 4.51944, 4.963623, 3.497131, 
    1.694122, 1.847961, 1.491058, 1.647003, 1.435913, 1.432739, 1.770447, 
    1.7789, 1.908478, 1.764954, 1.955475, 2.2052, 2.005463, 1.939453, 
    2.276947, 2.311676, 2.556244, 2.4375, 2.471344, 2.545074, 2.508209, 
    2.511932, 2.502014, 2.404694, 2.315613, 2.320251, 2.321228, 2.251709, 
    2.202087, 2.123169, 2.081848, 2.102356, 2.069855, 2.032288, 2.013153, 
    1.936523, 1.807556, 1.738586, 1.692505, 1.641663, 1.67688, 1.616058, 
    0.9051514, 1.046722, 1.809967, 1.991608, 1.548767, 2.311066, 3.846069, 
    3.855865, 3.486145, 3.649017, 3.726624, 3.528809, 3.659546, 3.693237, 
    2.946228, 2.580994, 2.547577, 2.514709, 2.372772, 1.995392, 1.337494, 
    0.5422363, 0.2342529, 0.5275879, 0.7936401, 0.9813232, 1.270447, 
    1.632599, 1.840424, 1.885681, 1.961914, 2.719788, 3.317902,
  2.546112, 2.198395, 2.205994, 2.379974, 2.352142, 2.807373, 3.302368, 
    3.612518, 3.431976, 3.399689, 3.215302, 4.375641, 3.886353, 2.599915, 
    3.134888, 3.49472, 3.649475, 3.150452, 3.276489, 2.600281, 1.938477, 
    1.339325, 1.284424, 1.566772, 2.330627, 2.20639, 1.703278, 1.898193, 
    1.863037, 1.640503, 1.516876, 1.625061, 1.8367, 2.115814, 2.013092, 
    1.991943, 2.385773, 2.413116, 3.067383, 3.667877, 3.649628, 3.196289, 
    2.735046, 2.450378, 2.273041, 2.177094, 2.13797, 2.198578, 2.27475, 
    2.326721, 2.274261, 2.16864, 2.133179, 2.155518, 2.106476, 2.015991, 
    1.864044, 1.738281, 1.687836, 1.623688, 1.610657, 1.650787, 1.546997, 
    0.7165527, 1.359833, 2.7276, 2.67981, 1.639954, 1.945709, 3.447968, 
    4.241394, 4.357117, 4.600372, 4.646454, 3.676697, 4.887573, 4.746948, 
    4.363068, 4.503815, 3.976074, 3.061584, 2.553619, 2.078186, 1.337799, 
    0.7760315, 0.5061035, 0.4348145, 0.3944702, 0.3182373, 0.6634827, 
    1.138794, 1.459839, 1.687744, 1.816742, 2.31424, 2.759186,
  2.161011, 2.605347, 2.879761, 3.065948, 3.199036, 3.494263, 3.576843, 
    3.877136, 4.038513, 3.772766, 3.522583, 3.612579, 3.513214, 3.102386, 
    2.198608, 2.296753, 1.57605, 1.55899, 1.609558, 1.543121, 1.745575, 
    1.652069, 1.631256, 1.332794, 1.251312, 0.8387451, 1.295563, 1.364777, 
    1.556396, 1.649872, 1.738983, 1.858459, 1.858612, 1.7948, 1.780151, 
    2.201965, 2.282104, 2.476898, 2.917358, 2.847351, 2.804688, 2.492584, 
    2.415588, 2.326538, 2.24234, 2.132935, 2.085754, 2.142914, 2.205444, 
    2.234375, 2.247253, 2.260101, 2.205139, 2.105286, 1.988403, 1.853943, 
    1.691925, 1.648041, 1.672943, 1.710785, 1.740417, 1.699646, 1.631287, 
    1.070129, 2.046692, 2.291748, 1.891266, 1.366882, 1.472656, 2.201263, 
    3.074463, 3.402527, 3.657501, 3.599731, 4.201996, 4.420441, 4.49173, 
    4.381317, 3.980469, 3.582703, 3.38208, 2.5672, 2.24353, 1.584778, 
    1.072388, 0.9002075, 0.6671448, 0.2417908, -0.1555176, -0.02578735, 
    0.596405, 1.186707, 1.600708, 1.778198, 1.913391, 2.134491,
  1.854584, 2.3237, 2.796295, 3.167908, 3.165771, 3.245239, 3.247711, 
    3.264404, 3.399475, 3.348053, 3.000854, 2.976685, 2.936829, 2.506653, 
    2.010498, 1.731812, 1.399078, 1.499939, 1.572327, 1.597717, 1.360809, 
    1.365753, 1.74649, 1.998566, 1.673492, 1.445007, 2.046112, 2.839142, 
    2.83783, 2.28894, 2.624146, 2.43457, 2.410614, 1.779694, 1.530914, 
    1.810791, 1.632477, 2.467834, 3.70462, 4.016541, 3.929688, 3.049011, 
    2.699219, 2.590698, 2.527344, 2.32486, 2.279572, 2.316345, 2.299347, 
    2.2323, 2.237701, 2.327789, 2.353851, 2.254425, 2.128845, 1.965881, 
    1.753845, 1.667755, 1.734192, 1.781525, 1.744751, 1.759521, 1.448029, 
    2.107025, 1.768311, 1.153961, 1.02832, 1.18399, 1.528778, 1.991333, 
    2.864197, 3.356201, 3.752686, 4.314697, 4.556976, 4.4039, 4.090942, 
    3.842377, 3.645752, 3.254944, 3.448853, 3.292755, 2.771698, 2.290619, 
    1.739197, 1.106384, 0.3314514, -0.4674988, -0.9579468, -0.7979431, 
    -0.02792358, 0.8173218, 1.436829, 1.710815, 1.744049, 1.749573,
  1.875092, 1.877655, 2.471619, 2.823059, 2.689728, 2.96405, 2.951752, 
    2.984894, 3.034576, 2.595306, 2.515106, 2.545197, 2.259583, 2.044006, 
    2.061646, 1.729675, 1.600739, 1.601898, 1.842194, 1.982422, 1.964386, 
    2.170288, 2.272858, 2.288086, 1.986572, 1.398438, 1.495789, 1.751312, 
    1.890961, 2.506317, 2.985931, 2.789764, 2.488983, 1.96524, 2.197449, 
    2.273712, 2.218628, 2.628784, 3.733002, 4.186096, 4.053131, 3.610168, 
    2.819336, 2.635864, 2.689056, 2.366486, 2.282959, 2.236267, 2.214386, 
    2.314301, 2.540619, 2.840424, 2.923645, 2.635284, 2.394531, 2.217194, 
    1.951935, 1.867828, 1.860748, 1.833832, 1.703796, 1.738342, 1.989594, 
    1.455231, 1.32724, 1.238922, 1.62558, 1.795898, 2.369385, 2.978699, 
    3.606964, 4.334961, 5.285736, 6.156952, 6.091003, 5.72049, 5.075653, 
    4.65976, 4.348877, 3.763977, 3.142365, 2.906525, 3.199951, 1.867188, 
    1.248505, 1.104156, 0.5565796, -0.3466797, -1.027222, -0.9544067, 
    -0.2460022, 0.6429443, 1.285522, 1.492035, 1.51236, 1.741211,
  1.345306, 1.503754, 1.522064, 2.465088, 2.613739, 2.670715, 2.198578, 
    3.375336, 3.212799, 3.155212, 3.285828, 2.957031, 2.750824, 2.554504, 
    2.4086, 2.590546, 2.358856, 1.932159, 1.629272, 1.740173, 2.151947, 
    2.080994, 2.614258, 2.64856, 2.46225, 2.069977, 2.126709, 2.356506, 
    2.51593, 2.664337, 2.750305, 2.640503, 2.303436, 1.946289, 1.748779, 
    2.019989, 2.338531, 3.01712, 3.977142, 3.944275, 3.038544, 2.306641, 
    2.364075, 2.410492, 2.674622, 2.826965, 3.364563, 3.926178, 4.250763, 
    4.612701, 4.86499, 4.39389, 3.457947, 3.044647, 2.66095, 2.1474, 
    2.040161, 2.018097, 1.917297, 1.781952, 2.413208, 2.1203, 1.543488, 
    1.3862, 1.505005, 1.771881, 2.008453, 2.443756, 3.099884, 3.79657, 
    4.462494, 5.409241, 5.443878, 5.95813, 6.28418, 6.291138, 6.003845, 
    5.322723, 4.65625, 3.984436, 3.171753, 2.802551, 1.666595, -0.1850891, 
    -0.1707153, 0.8041077, 1.308197, 0.873291, 0.3520813, 0.2177124, 
    0.4863281, 0.8516846, 1.134705, 1.2659, 1.340759, 1.402222,
  0.7839966, 0.9555969, 2.350128, 2.396484, 2.363342, 1.291473, 2.666595, 
    2.837067, 2.835236, 3.097473, 3.363739, 3.49707, 3.447083, 3.326965, 
    3.340485, 3.263489, 3.133209, 2.587097, 2.365479, 2.174866, 2.067993, 
    2.283447, 2.45697, 2.516449, 2.542175, 2.694733, 2.861053, 2.828705, 
    2.670776, 2.606445, 2.441223, 2.212799, 1.861206, 1.522705, 1.433411, 
    1.750183, 2.081879, 2.115967, 2.150635, 1.836304, 1.644409, 1.612671, 
    1.63855, 2.028564, 2.707397, 3.56427, 4.711975, 7.426178, 7.192108, 
    6.57663, 5.969391, 4.973511, 4.655212, 3.630157, 2.8013, 2.207092, 
    1.818024, 1.798767, 1.878754, 1.895691, 1.713928, 1.68631, 1.834625, 
    2.191162, 2.508545, 2.963409, 3.377472, 3.829437, 4.24649, 4.723907, 
    5.125519, 5.083801, 5.46994, 5.804962, 5.999084, 6.003143, 5.696564, 
    4.7323, 3.643311, 3.412506, 3.057495, 2.629883, 1.5625, 0.6989746, 
    1.06485, 0.325592, 0.5611267, 0.9093933, 1.145447, 1.221741, 1.220367, 
    0.821228, 0.09933472, 0.1554871, 0.6352844, 0.7571411,
  0.3575439, 0.4576111, 0.535614, 2.245697, 2.43457, 2.382355, 1.831238, 
    2.935364, 3.24472, 3.641144, 4.035217, 4.240936, 4.298248, 4.261322, 
    4.246674, 4.113037, 3.946106, 3.662292, 3.317322, 3.176758, 3.169128, 
    3.138458, 3.004028, 2.967834, 2.940613, 2.817627, 2.921997, 2.966095, 
    2.869385, 2.524139, 2.231628, 1.980011, 1.611725, 1.593231, 1.817108, 
    2.288635, 2.640259, 2.343903, 2.265442, 2.218048, 1.686722, 1.923706, 
    1.878922, 2.020844, 2.223587, 2.518219, 2.940491, 3.469513, 3.970306, 
    4.222473, 4.64621, 4.526123, 4.453003, 3.631073, 2.812622, 2.302979, 
    1.871613, 1.97403, 2.182373, 2.264893, 2.263611, 2.600586, 3.002228, 
    3.411591, 3.74292, 4.123505, 4.574097, 5.220245, 5.563232, 5.592468, 
    5.504181, 5.436676, 5.526169, 5.559341, 5.065521, 4.888046, 4.604889, 
    4.20575, 3.730621, 3.396255, 2.759888, 2.402527, 2.087097, 1.918823, 
    1.786011, 1.585693, 1.069672, 0.8192749, 0.604126, 1.573059, 2.508057, 
    2.732117, 1.574554, 0.3751831, -0.0001220703, 0.1077881,
  0.602417, 0.2645874, 0.1749878, -0.00793457, -0.5391541, 1.59552, 2.351563, 
    3.204895, 4.242828, 4.959503, 5.5401, 5.468933, 5.249146, 4.827942, 
    4.52359, 4.334076, 4.189606, 4.128403, 4.212967, 4.28537, 4.254959, 
    4.056778, 3.924881, 3.655426, 3.533554, 3.651184, 3.162979, 2.863174, 
    2.44931, 2.187637, 2.135818, 2.078735, 1.976181, 1.700348, 1.88205, 
    1.910828, 1.688873, 1.984665, 1.530807, 1.610367, 1.61557, 1.824356, 
    2.108871, 2.106415, 2.764084, 3.02092, 3.39592, 3.890839, 4.346298, 
    4.388092, 4.83342, 5.173431, 5.161835, 4.734711, 4.36673, 4.31134, 
    4.348114, 4.444611, 4.445709, 4.319214, 4.281921, 4.51358, 4.912689, 
    5.272125, 5.655426, 5.737564, 5.858795, 5.752487, 5.751373, 5.436005, 
    5.745132, 5.661072, 5.370987, 4.876068, 5.09436, 4.528931, 4.668243, 
    4.375992, 3.747025, 2.92775, 2.257996, 2.072601, 1.665955, 2.035294, 
    2.154434, 2.069351, 1.774628, 1.849167, 2.162628, 2.846863, 3.265106, 
    3.874695, 4.500061, 4.506378, 2.127167, 1.16095,
  2.355743, 1.428345, 0.861969, 0.6038513, 0.5992737, 1.039063, 2.129486, 
    3.801758, 6.276031, 7.696808, 7.936218, 7.441528, 6.289795, 5.272461, 
    4.652618, 4.617783, 4.00444, 4.108093, 4.128143, 4.41864, 4.412964, 
    4.237717, 4.076523, 3.896103, 3.643387, 3.443314, 3.168182, 2.66539, 
    2.581131, 2.184204, 2.236343, 2.035034, 2.02652, 1.786285, 1.418961, 
    1.25119, 1.292664, 1.219543, 1.788818, 2.122467, 1.823593, 2.006134, 
    2.255875, 2.477112, 2.720856, 2.896957, 3.068436, 3.318695, 3.661026, 
    3.990707, 4.32515, 4.644272, 4.933487, 5.184448, 5.465576, 5.673508, 
    5.85228, 5.946884, 5.921387, 5.842926, 5.690048, 5.510117, 5.277023, 
    5.613297, 5.397537, 5.34668, 5.43869, 5.308411, 5.513947, 5.04834, 
    5.647598, 5.579315, 4.685104, 4.965775, 4.83284, 4.491302, 4.030685, 
    3.397751, 2.941559, 2.607117, 2.250702, 2.305283, 2.169739, 2.250534, 
    2.011078, 1.660629, 1.119034, 0.9474792, 1.640503, 2.524246, 3.344452, 
    3.927856, 4.587311, 4.901093, 4.93222, 4.108582,
  4.90625, 4.055481, 3.345245, 3.622314, 5.01355, 6.897278, 7.756775, 
    7.087585, 6.85997, 6.43576, 6.032059, 5.5327, 4.985687, 4.418442, 
    4.01265, 3.871643, 3.783478, 3.824371, 3.930878, 3.965973, 3.877945, 
    3.799622, 3.620071, 3.467209, 3.195908, 3.658997, 3.479965, 2.997864, 
    3.002747, 2.992203, 2.641678, 2.032043, 1.795731, 1.611664, 1.529434, 
    1.579956, 1.709534, 1.84404, 2.07045, 2.207825, 2.46524, 2.720856, 
    2.995193, 3.150864, 3.260101, 3.362396, 3.514145, 3.698578, 3.916229, 
    4.195007, 4.522537, 4.881729, 5.238632, 5.599945, 5.829514, 6.054062, 
    6.214478, 6.286942, 6.345978, 6.461731, 6.483017, 6.575867, 6.583282, 
    6.569351, 6.580414, 6.143585, 6.050339, 5.889725, 5.741943, 5.826782, 
    5.596298, 5.278595, 5.045914, 4.986481, 4.720917, 3.947678, 3.63237, 
    3.381454, 3.527618, 3.228012, 2.991043, 2.903473, 2.83165, 2.777878, 
    2.564346, 2.179901, 2.031982, 2.177109, 2.51622, 3.198593, 3.820786, 
    4.231964, 4.530334, 4.768036, 4.865295, 5.147064,
  4.921371, 4.81012, 4.745987, 4.757507, 5.338043, 5.356003, 5.338562, 
    5.155746, 5.03862, 4.951904, 4.820526, 4.66832, 4.536346, 4.452621, 
    4.435699, 4.416489, 4.375275, 4.355362, 4.31662, 4.243256, 4.18335, 
    4.061417, 3.927628, 3.692657, 3.443253, 4.029572, 3.932373, 3.156921, 
    2.969406, 2.848465, 2.728271, 2.593964, 2.477097, 2.415909, 2.340439, 
    2.355804, 2.475998, 2.566025, 2.674362, 2.791824, 2.915771, 3.084259, 
    3.317719, 3.503464, 3.675217, 3.818314, 4.016495, 4.219223, 4.391098, 
    4.554764, 4.765839, 4.923584, 5.058029, 5.184921, 5.312897, 5.380081, 
    5.455673, 5.558731, 5.69812, 5.87027, 6.081131, 6.220901, 6.349106, 
    6.448914, 6.440506, 6.319748, 6.261658, 6.157761, 5.98616, 5.842331, 
    5.819092, 5.426712, 5.22612, 5.307892, 5.011353, 4.676178, 4.267654, 
    3.935379, 3.660309, 3.501648, 3.41069, 3.358154, 3.350281, 3.311401, 
    3.27417, 3.252686, 3.281723, 3.471115, 3.807053, 4.231659, 4.594421, 
    4.830353, 4.893768, 4.88739, 4.904312, 4.898575,
  4.908417, 4.722092, 4.57814, 4.441345, 4.256058, 4.129578, 4.047485, 
    3.99559, 3.928268, 3.884979, 3.873062, 3.864853, 3.874756, 3.87944, 
    3.886856, 3.885895, 3.880753, 3.852219, 3.806061, 3.73407, 3.655289, 
    3.556915, 3.485565, 3.401642, 3.367599, 3.336349, 3.250137, 3.191483, 
    3.119034, 3.072662, 3.129959, 3.13002, 3.144547, 3.179764, 3.22496, 
    3.23114, 3.236542, 3.277618, 3.318253, 3.396698, 3.47261, 3.572083, 
    3.637527, 3.721298, 3.789993, 3.878265, 3.97229, 4.094864, 4.202942, 
    4.345856, 4.495712, 4.651459, 4.799042, 4.907501, 4.996643, 5.071899, 
    5.153076, 5.258423, 5.401443, 5.530411, 5.62085, 5.736664, 5.893646, 
    6.002289, 6.072479, 6.100677, 6.12117, 6.121887, 6.045517, 5.992203, 
    5.96701, 5.872025, 5.907364, 5.972488, 5.827698, 5.737915, 5.696762, 
    5.571121, 5.537262, 5.629242, 5.623322, 5.533279, 5.656006, 5.616501, 
    5.616104, 5.593185, 5.592911, 5.616302, 5.735687, 5.720337, 5.666611, 
    5.664932, 5.48439, 5.295654, 5.142792, 5.014862,
  4.799881, 4.656525, 4.552094, 4.466873, 4.401443, 4.339478, 4.268829, 
    4.205734, 4.167587, 4.135696, 4.120453, 4.103333, 4.068695, 4.062195, 
    4.025406, 3.992004, 3.980087, 3.981201, 3.96817, 3.932632, 3.913422, 
    3.880234, 3.900024, 3.902298, 3.892853, 3.875931, 3.870453, 3.880875, 
    3.861938, 3.860748, 3.857956, 3.8517, 3.84462, 3.842529, 3.854828, 
    3.903015, 3.95314, 3.979309, 3.973846, 4.006927, 4.024628, 4.045578, 
    4.096039, 4.130035, 4.152161, 4.166824, 4.216995, 4.259262, 4.300659, 
    4.362198, 4.417847, 4.483032, 4.543442, 4.590057, 4.609131, 4.658554, 
    4.723587, 4.773376, 4.81694, 4.871231, 4.905289, 4.92392, 4.965317, 
    5.010117, 5.05275, 5.107437, 5.173309, 5.214859, 5.25502, 5.282166, 
    5.309723, 5.305557, 5.304764, 5.321625, 5.333618, 5.348785, 5.363617, 
    5.349365, 5.327545, 5.307251, 5.280807, 5.254318, 5.253922, 5.249039, 
    5.239532, 5.238892, 5.237839, 5.22612, 5.18367, 5.156982, 5.128723, 
    5.110703, 5.042328, 4.961151, 4.903656, 4.862778,
  2.324051, 2.33168, 2.34697, 2.372559, 2.40062, 2.432846, 2.468582, 
    2.511154, 2.559937, 2.613174, 2.658752, 2.704269, 2.750549, 2.79567, 
    2.841949, 2.885056, 2.921387, 2.948669, 2.966583, 2.973145, 2.97464, 
    2.975235, 2.975296, 2.979324, 2.982971, 2.990067, 2.998077, 3.009857, 
    3.018127, 3.029663, 3.037857, 3.045853, 3.055115, 3.063049, 3.058563, 
    3.059341, 3.058563, 3.049835, 3.039551, 3.029724, 3.018005, 3.007141, 
    2.995865, 2.981995, 2.965271, 2.94574, 2.93187, 2.925156, 2.913116, 
    2.912659, 2.903275, 2.909866, 2.947815, 2.990723, 2.96846, 3.000626, 
    3.038116, 3.077957, 3.076141, 2.977707, 2.991241, 3.076019, 2.947113, 
    2.924454, 2.881348, 2.844177, 2.803619, 2.781219, 2.759995, 2.730759, 
    2.725357, 2.726532, 2.730759, 2.798798, 2.745804, 2.741058, 2.731491, 
    2.836548, 2.681671, 2.678818, 2.649063, 2.624588, 2.593201, 2.566574, 
    2.536163, 2.505249, 2.47641, 2.448273, 2.423462, 2.401535, 2.381805, 
    2.363312, 2.342865, 2.331421, 2.325821, 2.324188,
  2.290527, 2.364365, 2.428619, 2.489426, 2.558624, 2.647232, 2.729523, 
    2.811874, 2.87561, 2.91658, 2.946381, 2.971909, 2.978226, 2.971069, 
    2.97171, 2.981415, 2.972031, 2.941177, 2.900681, 2.809982, 2.719177, 
    2.621841, 2.545929, 2.500549, 2.498459, 2.547165, 2.623276, 2.705429, 
    2.778412, 2.848343, 2.914093, 2.968323, 3.004532, 3.021332, 3.018585, 
    3.00354, 2.982849, 2.962143, 2.936752, 2.915649, 2.906403, 2.865997, 
    2.841507, 2.796982, 2.784286, 2.807129, 2.788574, 2.804718, 2.815918, 
    2.83168, 2.822235, 2.786285, 2.781219, 2.719238, 2.82666, 2.654861, 
    2.632324, 2.637787, 2.669037, 2.723923, 2.766037, 2.826538, 2.883942, 
    2.96019, 2.965393, 2.883301, 2.786224, 2.652191, 2.52269, 2.499252, 
    2.554382, 2.664032, 2.73201, 2.750092, 2.713898, 2.691437, 2.695541, 
    2.70668, 2.740463, 2.671387, 2.64267, 2.650421, 2.518845, 2.454132, 
    2.418976, 2.363129, 2.203613, 2.120987, 2.069565, 2.043381, 2.033051, 
    2.045273, 2.065979, 2.102371, 2.152832, 2.220734,
  2.189041, 2.193588, 2.265472, 2.378815, 2.478165, 2.643463, 2.865723, 
    3.04097, 3.103867, 3.157333, 3.225677, 3.193649, 3.045349, 2.86409, 
    2.686554, 2.574448, 2.556351, 2.60791, 2.711548, 2.867798, 3.128418, 
    3.393646, 3.512146, 3.299713, 2.853485, 2.469376, 2.424057, 2.532852, 
    2.696259, 2.863235, 2.983109, 3.062271, 3.099503, 3.073471, 3.012985, 
    2.97731, 2.993393, 3.024841, 3.051849, 3.070602, 3.101135, 3.174515, 
    3.27861, 3.492096, 3.682327, 3.785767, 3.693985, 3.538437, 3.496506, 
    3.451599, 3.368912, 3.205826, 2.988373, 2.687332, 2.438828, 2.236237, 
    2.010773, 1.813934, 1.68541, 1.624863, 1.658539, 1.835342, 2.123962, 
    2.402573, 2.599319, 2.658951, 2.743912, 2.790787, 2.795746, 2.760513, 
    2.803802, 2.86058, 2.917679, 2.986038, 3.016495, 2.972305, 2.916367, 
    2.854919, 2.715195, 2.618057, 2.569763, 2.543839, 2.414612, 2.263779, 
    2.101074, 1.986938, 1.925034, 1.87529, 1.941101, 2.095352, 2.034607, 
    2.078873, 2.080368, 2.103943, 2.159592, 2.17392,
  2.709015, 3.048859, 3.25882, 3.21637, 2.969833, 2.690918, 2.438843, 
    2.280243, 2.165726, 2.076324, 2.099319, 2.180634, 2.349442, 2.509277, 
    2.64801, 2.881287, 3.154327, 3.391953, 3.479385, 3.209213, 2.866119, 
    2.672821, 2.596985, 2.646713, 2.766174, 2.744766, 2.657776, 2.749313, 
    2.954193, 3.169571, 3.372375, 3.48317, 3.480759, 3.428741, 3.397369, 
    3.316895, 3.12204, 2.899368, 2.766052, 2.817932, 2.848785, 2.75412, 
    2.671707, 2.746445, 3.117081, 3.480698, 2.357285, 2.403091, 2.63887, 
    2.78418, 2.699539, 2.549606, 2.411911, 2.249741, 1.979813, 1.924088, 
    2.161987, 1.370438, 1.492508, 1.896545, 2.34758, 2.700653, 2.916733, 
    3.002808, 3.0401, 2.916672, 2.8004, 2.793884, 2.955338, 3.120239, 
    3.316727, 3.492905, 3.638107, 3.775803, 3.885513, 3.947617, 4.001923, 
    4.070084, 4.104202, 4.128281, 4.160995, 4.126617, 3.870773, 3.69075, 
    3.522659, 3.591202, 3.809433, 4.236786, 4.690689, 3.293655, 2.834503, 
    2.444107, 2.226593, 2.101013, 2.086487, 2.331024,
  2.184601, 2.246201, 2.284851, 2.226013, 2.213837, 2.316757, 2.458832, 
    2.612656, 2.847046, 2.957581, 2.995605, 2.943588, 2.944946, 2.921387, 
    2.892548, 2.950562, 3.146576, 3.206665, 3.029663, 2.760132, 2.595215, 
    2.529785, 2.455765, 2.672104, 3.102631, 3.38533, 3.345032, 3.261612, 
    3.288895, 3.260254, 3.309219, 3.558167, 3.780121, 3.847763, 3.740189, 
    3.667145, 3.630173, 3.567673, 3.394226, 3.209015, 3.117477, 3.14859, 
    3.111877, 3.063171, 3.004196, 3.078354, 2.526077, 2.392441, 2.16153, 
    1.907745, 1.673767, 1.462372, 1.291672, 1.300522, 1.376312, 1.419327, 
    1.597198, 1.774002, 2.121048, 2.573853, 3.001785, 3.300156, 3.393387, 
    3.496323, 3.632355, 3.811447, 4.052429, 4.198135, 4.336243, 4.304382, 
    5.682739, 5.590546, 5.624268, 5.511703, 5.295486, 4.866516, 5.898239, 
    5.796097, 5.719391, 5.593552, 5.432693, 4.971878, 4.612488, 4.362167, 
    4.291077, 4.399811, 4.725327, 5.017776, 5.234756, 5.337616, 4.839508, 
    4.075165, 3.095627, 2.605072, 2.327988, 2.154984,
  6.95575, 5.244431, 5.40097, 4.845779, 4.172195, 3.608658, 3.424728, 
    3.737228, 3.998566, 4.222458, 4.471161, 4.212494, 3.68808, 3.227829, 
    2.64769, 2.115341, 1.65596, 1.47171, 1.576721, 2.004715, 1.953156, 
    1.781021, 1.649475, 1.794235, 1.941376, 2.001144, 2.02359, 2.037476, 
    2.021057, 1.998932, 1.934143, 1.868454, 1.889877, 1.965332, 2.052765, 
    2.16951, 2.265594, 2.235916, 2.081421, 2.001266, 2.02034, 2.04509, 
    2.210907, 2.258224, 1.800262, 1.78067, 1.595108, 1.248962, 0.9138641, 
    0.5332947, 0.1375122, -0.0463562, 0.0262146, 0.301239, 0.6862488, 
    1.09903, 1.523499, 2.013428, 2.617004, 3.162689, 3.653717, 4.1026, 
    4.477539, 4.891479, 5.3237, 5.741089, 6.151947, 6.700073, 7.332428, 
    8.01828, 8.782471, 8.606873, 8.363434, 8.053802, 7.661865, 7.030701, 
    6.336792, 5.544281, 6.083237, 6.020935, 6.167511, 5.712418, 5.303833, 
    5.052414, 4.979935, 5.064163, 5.377182, 5.770554, 6.206543, 6.71376, 
    7.109619, 7.511551, 7.886749, 7.927917, 7.770142, 7.477646,
  12.52255, 12.68436, 12.82626, 12.67548, 12.47839, 12.10873, 11.59732, 
    11.056, 10.66812, 10.66678, 11.056, 11.50287, 11.79428, 11.79453, 
    11.25684, 9.746414, 8.052551, 6.862396, 6.476044, 6.548172, 6.3983, 
    5.908508, 5.323273, 4.663177, 3.92749, 3.351181, 2.931274, 2.857239, 
    2.849945, 2.854645, 2.749817, 1.961517, 1.469208, 1.50914, 2.008591, 
    2.901367, 5.520309, 5.95755, 5.814911, 5.069122, 4.09024, 3.633514, 
    3.573639, 3.155579, 2.109772, 0.7685547, -0.1946106, -0.5730286, 
    -0.486908, -0.3189697, -0.2883301, -0.3061218, -0.3365173, -0.2220764, 
    -0.0463562, 0.1487732, 0.3726807, 0.5848999, 0.8644714, 1.114319, 
    1.257233, 1.286835, 1.334198, 1.457428, 1.616425, 1.787811, 1.971283, 
    2.175659, 2.385162, 2.581329, 2.819, 3.084686, 3.364716, 3.522644, 
    3.56189, 3.59549, 3.779633, 4.603912, 6.065521, 7.998566, 7.490601, 
    6.884583, 6.461243, 6.381317, 6.984894, 7.573883, 8.176544, 8.63736, 
    8.909393, 9.162933, 9.327576, 9.704254, 10.25269, 10.8634, 11.49957, 
    12.07983,
  6.263489, 5.878906, 5.401367, 4.914978, 4.458771, 4.039734, 3.555847, 
    3.239532, 3.067963, 2.950012, 2.865173, 2.850769, 2.968567, 3.197113, 
    3.451935, 3.681885, 3.827423, 3.956299, 4.223328, 4.636627, 4.811401, 
    4.605255, 4.152222, 3.347931, 2.541199, 2.034119, 1.69397, 1.33548, 
    1.065155, 0.8879395, 0.776825, 0.6679688, 0.5508728, 0.5638733, 
    0.7171936, 0.9535217, 1.21463, 1.349396, 1.381775, 1.433716, 1.516144, 
    1.560333, 1.436707, 1.24295, 1.040619, 0.703064, 0.2259216, -0.1494141, 
    -0.2342224, -0.1991577, -0.1507874, -0.1153564, -0.09869385, -0.06497192, 
    0.002685547, 0.09887695, 0.2255249, 0.3662109, 0.5142517, 0.6243286, 
    0.6738892, 0.7309875, 0.8086548, 0.9294128, 1.087219, 1.255463, 1.422913, 
    1.604095, 1.77121, 1.890839, 1.983673, 2.098053, 2.211243, 2.318024, 
    2.3862, 2.380981, 2.321106, 2.273041, 2.29071, 2.351807, 2.517517, 
    3.239258, 3.881226, 3.595123, 3.677124, 4.263855, 5.123291, 5.973694, 
    6.532013, 6.693024, 6.604889, 6.606842, 6.672485, 6.68869, 6.600983, 
    6.47818,
  2.139374, 2.061737, 1.958282, 1.854156, 1.755341, 1.680786, 1.618164, 
    1.579041, 1.574036, 1.575867, 1.586182, 1.64212, 1.700653, 1.729187, 
    1.757416, 1.799561, 1.864807, 1.937439, 1.976807, 1.93277, 1.78302, 
    1.642151, 1.53125, 1.456573, 1.423431, 1.389557, 1.348236, 1.300903, 
    1.221039, 1.137482, 1.082153, 1.010284, 0.9082642, 0.8309937, 0.8022156, 
    0.7810974, 0.8065186, 0.870697, 0.9688721, 1.103912, 1.201813, 1.264771, 
    1.324036, 1.33313, 1.276642, 1.198242, 1.015503, 0.6772156, 0.3155518, 
    0.09341431, 0.03430176, 0.05911255, 0.08914185, 0.09747314, 0.1121826, 
    0.1634216, 0.2059326, 0.290863, 0.4223328, 0.5371704, 0.5809326, 
    0.6063843, 0.6723938, 0.7893982, 0.9478455, 1.202667, 1.465057, 1.666748, 
    1.79184, 1.883606, 1.968628, 2.066406, 2.155975, 2.240051, 2.276428, 
    2.1875, 1.946869, 1.796021, 1.751495, 1.76413, 1.852936, 2.086731, 
    2.225891, 1.892975, 1.615753, 1.590546, 1.691345, 1.88443, 2.091034, 
    2.159912, 2.16864, 2.217651, 2.265564, 2.271881, 2.227417, 2.18515,
  1.650391, 1.750458, 1.880859, 1.943024, 1.909454, 1.841736, 1.788879, 
    1.734375, 1.677002, 1.615173, 1.590363, 1.675446, 1.796997, 1.859253, 
    1.923615, 2.033722, 2.187225, 2.314606, 2.268097, 2.045837, 1.848846, 
    1.734009, 1.609833, 1.508453, 1.507233, 1.623505, 1.795837, 1.908386, 
    1.907288, 1.854828, 1.731964, 1.531769, 1.343842, 1.235291, 1.181305, 
    1.13443, 1.123352, 1.156311, 1.205078, 1.258148, 1.353455, 1.492706, 
    1.602081, 1.587097, 1.577087, 1.571533, 1.375519, 1.075317, 0.7350464, 
    0.4633484, 0.3632813, 0.3954468, 0.4145203, 0.3671265, 0.3316345, 
    0.3625183, 0.4499207, 0.5459595, 0.630127, 0.6921997, 0.7253418, 
    0.7756348, 0.8591919, 0.9524536, 1.108337, 1.342499, 1.549622, 1.653503, 
    1.703583, 1.769348, 1.863861, 1.95343, 2.04361, 2.101105, 2.023315, 
    1.742249, 1.719086, 2.651367, 2.615814, 1.849945, 1.763214, 1.792175, 
    1.820068, 1.582306, 1.387054, 1.384613, 1.548126, 1.688354, 1.733154, 
    1.719635, 1.734772, 1.772125, 1.794464, 1.78894, 1.723633, 1.643097,
  1.954346, 2.06076, 2.175018, 2.232666, 2.239777, 2.235199, 2.241852, 
    2.246613, 2.187317, 2.135803, 2.147003, 2.183533, 2.206055, 2.203308, 
    2.227722, 2.34726, 2.543762, 2.707092, 2.662048, 2.496918, 2.495972, 
    2.646423, 2.611603, 2.431458, 2.381287, 2.511597, 2.64798, 2.678894, 
    2.658386, 2.568817, 2.335358, 2.023712, 1.843292, 1.741669, 1.605011, 
    1.458344, 1.375916, 1.361664, 1.406067, 1.555328, 1.730164, 1.784119, 
    1.743225, 1.774994, 1.932007, 1.938385, 1.724945, 1.385223, 1.093475, 
    0.859375, 0.7871094, 0.8876953, 0.9724426, 0.9328613, 0.8758545, 
    0.9029846, 0.9632263, 1.023499, 1.098877, 1.145844, 1.163177, 1.221405, 
    1.267456, 1.324554, 1.403503, 1.506897, 1.591675, 1.667114, 1.757385, 
    1.895752, 1.994537, 2.009857, 2.01947, 2.005859, 1.881744, 1.763428, 
    2.400665, 2.474792, 1.941803, 1.817169, 1.652466, 1.594452, 1.5914, 
    1.4552, 1.347412, 1.543671, 1.802521, 1.922699, 1.926544, 1.913849, 
    1.944855, 1.951965, 1.95575, 1.990356, 1.992584, 1.940765,
  2.282959, 2.354797, 2.410309, 2.433136, 2.451355, 2.536438, 2.689392, 
    2.794525, 2.790558, 2.827423, 2.933197, 3.000061, 2.991791, 2.979553, 
    2.91745, 2.854614, 2.946289, 3.167389, 3.233398, 3.361847, 3.630615, 
    3.693176, 3.26651, 2.676361, 2.335663, 2.183929, 2.069092, 2.048096, 
    2.070435, 1.927216, 1.752808, 1.705078, 1.751617, 1.788757, 1.77124, 
    1.728058, 1.703186, 1.683228, 1.703979, 1.913483, 2.269226, 2.293701, 
    2.105011, 2.135956, 2.391327, 2.54892, 2.038605, 1.728241, 1.572662, 
    1.453522, 1.516785, 1.661987, 1.735291, 1.678986, 1.596375, 1.547607, 
    1.502533, 1.486206, 1.519287, 1.524139, 1.532166, 1.543091, 1.54837, 
    1.586853, 1.649933, 1.675079, 1.723053, 1.831573, 1.912415, 1.961792, 
    1.982483, 1.973572, 1.969147, 1.905731, 1.8013, 1.769012, 2.171692, 
    2.178864, 2.128265, 1.875214, 1.709442, 1.488678, 1.368561, 1.219025, 
    1.262177, 1.629303, 1.976654, 2.132141, 2.133545, 2.06308, 2.027802, 
    2.055084, 2.063995, 2.054932, 2.093811, 2.186798,
  2.555908, 2.539001, 2.504669, 2.521301, 2.648895, 2.997528, 3.442322, 
    3.678314, 3.78125, 3.913544, 4.020233, 3.839783, 3.414734, 3.111725, 
    2.94986, 2.9086, 2.963287, 3.068756, 3.19455, 3.303528, 3.262756, 
    2.821472, 2.061188, 1.406769, 1.119537, 1.206757, 1.515991, 1.798645, 
    1.888214, 1.905273, 1.966553, 2.024994, 2.03125, 1.992706, 2.004883, 
    2.000061, 1.986328, 2.031036, 1.942902, 2.269775, 2.853638, 2.896027, 
    2.620331, 2.539734, 2.686584, 2.831451, 2.509369, 2.439728, 2.441742, 
    2.509308, 2.686005, 2.685303, 2.484039, 2.271545, 2.092834, 1.931335, 
    1.827332, 1.81897, 1.843109, 1.819092, 1.7854, 1.769196, 1.761597, 
    1.793762, 1.819519, 1.806946, 1.839783, 1.917969, 1.972473, 2.015961, 
    2.044342, 2.022736, 1.968964, 1.876678, 1.791748, 1.694458, 1.56955, 
    1.511871, 1.612701, 1.859436, 1.733582, 1.689392, 1.772583, 1.852356, 
    1.896423, 1.993439, 2.113617, 2.139587, 2.144928, 2.14975, 2.155396, 
    2.247223, 2.277466, 2.249115, 2.326172, 2.467133,
  2.401886, 2.352264, 2.324219, 2.460938, 2.750854, 3.041534, 3.119659, 
    3.383331, 3.361206, 3.314392, 2.92511, 2.432617, 2.0177, 1.841156, 
    1.830383, 1.946228, 2.080414, 2.160156, 2.139343, 1.935364, 1.671692, 
    1.440613, 1.356567, 1.480377, 1.670105, 1.922852, 2.132813, 2.208374, 
    2.29538, 2.405792, 2.23407, 2.103699, 1.985352, 1.873322, 2.123169, 
    2.289886, 2.129639, 2.182922, 2.27063, 2.478607, 2.880066, 3.385864, 
    3.321991, 2.979034, 2.891724, 2.93866, 2.851501, 2.383453, 2.525055, 
    2.362823, 2.191803, 2.183136, 2.171295, 2.185364, 2.184509, 2.113129, 
    2.056061, 2.048248, 2.050598, 2.020569, 1.98465, 1.9711, 1.985107, 
    1.978516, 1.993683, 2.015625, 2.037323, 2.041687, 2.037903, 2.050568, 
    2.013397, 1.943146, 1.870056, 1.746552, 1.661133, 1.496552, 1.205139, 
    1.046875, 1.570068, 1.903656, 1.726746, 1.933411, 2.35144, 2.50473, 
    2.326599, 2.09549, 2.045258, 2.047791, 2.084045, 2.124756, 2.128754, 
    2.179504, 2.177826, 2.154938, 2.225433, 2.338013,
  2.262512, 2.162201, 2.076813, 2.108521, 2.203247, 2.364563, 2.525848, 
    2.333527, 2.249786, 2.232697, 1.465637, 1.360809, 1.417175, 1.49472, 
    1.529968, 1.672516, 1.847961, 1.899597, 1.849304, 1.753448, 1.812744, 
    2.00528, 2.144165, 2.297638, 2.390167, 2.392059, 2.381409, 2.348816, 
    2.367126, 2.187958, 1.814728, 1.807037, 1.830139, 1.873352, 2.096924, 
    2.166168, 2.088928, 2.489014, 2.601257, 2.651825, 2.71817, 3.061401, 
    3.510284, 3.266266, 2.960785, 2.917969, 2.683411, 2.369843, 2.036804, 
    1.646729, 1.681335, 1.945099, 2.152985, 2.256989, 2.292969, 2.243896, 
    2.198242, 2.14212, 2.106903, 2.122772, 2.12085, 2.104889, 2.108154, 
    2.112305, 2.101501, 2.072479, 1.992065, 1.927917, 1.90506, 1.845428, 
    1.752991, 1.659943, 1.539398, 1.394867, 1.229889, 0.9809875, 0.8779297, 
    1.965363, 2.212677, 2.011383, 2.067566, 2.478058, 2.48761, 2.519135, 
    2.323639, 2.028198, 1.985962, 2.048889, 2.096466, 2.128906, 2.13974, 
    2.16861, 2.112701, 2.128235, 2.202667, 2.237305,
  1.836517, 1.758331, 1.684235, 1.725189, 1.918884, 3.672577, 3.929565, 
    3.725342, 3.251343, 2.168762, 2.037048, 2.128174, 2.129639, 2.056458, 
    2.055817, 2.190125, 2.289917, 2.269775, 2.243042, 2.302155, 2.396301, 
    2.486115, 2.451355, 2.431976, 2.395416, 2.299927, 2.237762, 2.127533, 
    2.061066, 1.861786, 1.816772, 2.269989, 2.435547, 2.611908, 2.883148, 
    2.927979, 3.029877, 3.142883, 3.54837, 3.543549, 3.348358, 2.663788, 
    2.389984, 2.376617, 2.398621, 2.315948, 2.136047, 1.886261, 1.821808, 
    1.9646, 2.172546, 2.3237, 2.317444, 2.264252, 2.262085, 2.241852, 
    2.209961, 2.159119, 2.097443, 2.107819, 2.123383, 2.135529, 2.11438, 
    2.068939, 1.986084, 1.865234, 1.739838, 1.593292, 1.516418, 1.412018, 
    1.286377, 1.21759, 1.05722, 0.9580688, 0.8261719, 0.738739, 1.191223, 
    2.693359, 3.091858, 2.34375, 2.17807, 2.951233, 3.042114, 2.472015, 
    2.326294, 2.152466, 2.187042, 2.290039, 2.272614, 2.191132, 2.115875, 
    2.056641, 1.984039, 2.000061, 1.97168, 1.910614,
  1.487244, 1.487244, 1.671539, 1.927338, 2.520294, 4.152405, 4.173126, 
    3.691528, 3.136475, 2.159454, 1.992859, 2.164459, 2.17749, 2.095245, 
    2.202454, 2.411011, 2.565155, 2.534241, 2.49588, 2.479492, 2.439514, 
    2.359375, 2.270844, 2.155518, 2.082764, 2.001801, 1.939728, 1.929626, 
    2.034821, 2.091797, 2.313477, 3.265808, 3.289001, 3.31778, 3.344147, 
    3.293091, 3.115997, 3.304474, 3.309784, 3.686401, 3.494263, 2.258362, 
    1.949554, 2.022339, 2.200592, 2.273438, 2.228119, 2.182404, 2.222137, 
    2.296295, 2.281647, 2.266083, 2.251953, 2.238373, 2.230194, 2.238464, 
    2.192139, 2.172485, 2.128906, 2.09552, 2.061066, 2.018097, 1.969269, 
    1.868622, 1.702087, 1.513, 1.386719, 1.225922, 1.159363, 1.086578, 
    1.009827, 1.039185, 0.9532776, 0.8440247, 0.7521973, 0.9789124, 1.88504, 
    3.527161, 3.683411, 2.958588, 2.73999, 3.228638, 3.412109, 3.087677, 
    2.443817, 2.20929, 2.194244, 2.274353, 2.186005, 2.100006, 2.011871, 
    1.900787, 1.825836, 1.744598, 1.634705, 1.523621,
  1.691284, 1.882813, 2.238678, 2.741852, 4.271484, 4.105865, 4.105408, 
    3.979431, 3.428772, 3.301941, 2.048889, 2.101563, 2.959686, 2.256226, 
    2.343933, 2.40448, 2.446472, 2.449158, 2.403778, 2.358795, 2.302338, 
    2.204895, 2.123199, 2.096344, 2.069061, 2.073639, 2.113617, 2.276123, 
    2.381958, 2.542206, 2.762451, 3.722839, 4.123566, 4.130798, 3.800018, 
    3.39621, 3.496674, 3.358215, 3.542969, 3.553406, 3.306976, 2.287903, 
    2.435211, 2.581299, 2.496216, 2.386261, 2.293091, 2.254547, 2.192322, 
    2.16098, 2.171356, 2.200989, 2.25293, 2.265961, 2.267975, 2.238129, 
    2.221832, 2.200592, 2.154816, 2.109894, 2.01889, 1.915039, 1.816925, 
    1.658997, 1.497711, 1.280853, 1.111145, 1.066864, 1.017273, 0.973114, 
    1.000427, 0.9569092, 0.9214783, 0.9003906, 1.009094, 1.398743, 2.320892, 
    4.097351, 3.711212, 3.388489, 3.301636, 3.555786, 3.816986, 3.153259, 
    2.938629, 2.300507, 2.049988, 2.060089, 1.944916, 1.854645, 1.753784, 
    1.658081, 1.599854, 1.550964, 1.538879, 1.561859,
  2.107147, 2.338745, 2.498169, 2.696747, 4.134369, 3.534302, 3.807861, 
    3.974335, 3.30542, 3.17865, 2.069275, 2.080994, 3.227478, 2.97937, 
    2.260559, 2.302094, 2.298828, 2.278839, 2.293182, 2.260284, 2.250854, 
    2.239594, 2.241394, 2.275269, 2.300262, 2.382111, 2.483978, 2.567139, 
    2.597076, 2.72168, 2.843231, 2.933655, 4.075714, 4.165314, 3.962311, 
    3.681519, 3.683319, 3.758148, 3.67395, 3.077545, 2.399078, 2.446564, 
    2.581696, 2.615875, 2.499023, 2.411011, 2.337433, 2.292389, 2.22168, 
    2.194092, 2.221008, 2.24646, 2.294647, 2.330658, 2.340942, 2.323364, 
    2.316284, 2.263458, 2.190033, 2.079987, 1.981262, 1.867004, 1.724274, 
    1.538086, 1.383148, 1.277069, 1.218994, 1.16864, 1.169708, 1.177216, 
    1.217773, 1.210938, 1.223755, 1.3461, 1.432373, 1.680786, 2.386536, 
    4.244781, 3.690155, 3.301514, 3.385284, 3.739014, 3.983185, 3.173218, 
    3.065613, 3.1521, 2.045959, 1.997345, 1.875336, 1.799286, 1.712646, 
    1.727417, 1.722778, 1.79129, 1.878448, 1.951874,
  2.508728, 2.647583, 2.516235, 2.538483, 4.296021, 3.721802, 3.703857, 
    4.080597, 3.703308, 3.175201, 2.943939, 2.313477, 3.403107, 3.207703, 
    2.247253, 2.169617, 2.201172, 2.2276, 2.213867, 2.27417, 2.327087, 
    2.361206, 2.369324, 2.41095, 2.466553, 2.527924, 2.567444, 2.607117, 
    2.654816, 2.689636, 2.737427, 2.804138, 2.904816, 3.799286, 4.179016, 
    3.59726, 3.391846, 2.766663, 2.820374, 2.480103, 2.421875, 2.577606, 
    2.621887, 2.576111, 2.457703, 2.36969, 2.32782, 2.272369, 2.19986, 
    2.161652, 2.197327, 2.226349, 2.272186, 2.309753, 2.300964, 2.233459, 
    2.194, 2.138672, 2.071228, 2.001434, 1.916534, 1.821228, 1.750641, 
    1.673615, 1.631439, 1.618256, 1.603668, 1.602203, 1.597534, 1.601105, 
    1.601959, 1.636932, 1.647705, 1.808411, 1.919556, 2.252075, 4.145752, 
    4.404602, 3.378326, 3.486328, 3.891144, 3.700958, 3.613037, 3.19278, 
    3.361786, 2.866608, 1.999695, 1.983337, 1.962891, 1.922638, 1.939697, 
    2.046295, 2.123505, 2.220367, 2.308533, 2.377808,
  2.640106, 2.596039, 2.411377, 2.376373, 3.42514, 3.571014, 3.421814, 
    3.493683, 3.389832, 3.214722, 3.201111, 2.392761, 2.467438, 2.319275, 
    2.119568, 2.068359, 2.088348, 2.190674, 2.157166, 2.250977, 2.319275, 
    2.355713, 2.38092, 2.4151, 2.494141, 2.55249, 2.587067, 2.559296, 
    2.550537, 2.572693, 2.628143, 2.612854, 2.537476, 2.620667, 2.721008, 
    2.708405, 2.998047, 2.463867, 2.49707, 2.32785, 2.314606, 2.54303, 
    2.555725, 2.495575, 2.355011, 2.230591, 2.179901, 2.166351, 2.159119, 
    2.158203, 2.138672, 2.075592, 2.064972, 2.12323, 2.175934, 2.189209, 
    2.161255, 2.128967, 2.099823, 2.076508, 2.040039, 2.056366, 2.038879, 
    2.004883, 2.014282, 2.018433, 2.008331, 2.039337, 2.080597, 2.15918, 
    2.18158, 2.218292, 2.234711, 2.34317, 2.41452, 3.23111, 3.54718, 
    3.411591, 3.334381, 3.783142, 3.931702, 3.880463, 3.611176, 3.293304, 
    3.077545, 2.62616, 2.042328, 2.103577, 2.149292, 2.156677, 2.209442, 
    2.293823, 2.399994, 2.472961, 2.526093, 2.630219,
  2.556641, 2.506714, 2.3349, 2.30423, 2.959747, 3.486542, 3.222656, 
    3.212616, 3.273712, 3.221924, 3.257477, 2.394135, 2.441071, 2.255463, 
    2.133331, 2.196411, 2.194336, 2.273712, 2.291779, 2.369934, 2.427277, 
    2.487061, 2.478333, 2.433594, 2.483978, 2.542816, 2.478363, 2.343262, 
    2.306915, 2.442352, 2.478821, 2.482452, 2.514496, 2.509064, 2.461578, 
    2.443604, 2.352844, 2.3237, 2.752258, 2.318359, 2.37384, 2.469025, 
    2.421112, 2.36911, 2.219238, 2.013336, 1.963135, 2.025848, 2.075958, 
    2.066925, 2.045715, 1.983643, 1.938416, 1.991791, 2.086914, 2.100128, 
    2.07547, 2.100891, 2.097382, 2.105408, 2.069733, 2.091522, 2.107941, 
    2.12088, 2.131378, 2.156036, 2.194397, 2.273651, 2.353912, 2.433136, 
    2.476044, 2.503235, 2.525269, 2.490631, 2.399811, 3.162048, 3.547852, 
    4.176697, 4.02948, 3.758148, 3.641907, 3.731445, 3.274719, 3.175537, 
    3.145233, 2.786652, 2.684326, 2.162231, 2.169006, 2.184875, 2.209045, 
    2.229126, 2.393494, 2.480011, 2.552399, 2.577576,
  2.423889, 2.381287, 2.250305, 2.480652, 3.1203, 3.004211, 3.019257, 
    2.799561, 2.901428, 2.770172, 2.733917, 2.313721, 2.274963, 2.227692, 
    2.231842, 2.332947, 2.413971, 2.423279, 2.457642, 2.46463, 2.463287, 
    2.559631, 2.577637, 2.578735, 2.564484, 2.570801, 2.419342, 2.290405, 
    2.703735, 2.363251, 2.287201, 2.283386, 2.352173, 2.368622, 2.381866, 
    2.349701, 2.130341, 2.493317, 2.46991, 2.456329, 2.275513, 2.231842, 
    2.216492, 2.195618, 2.098022, 2.016693, 2.002838, 2.044006, 2.082642, 
    2.079651, 2.087982, 2.094147, 2.074707, 2.080231, 2.097687, 2.121429, 
    2.11087, 2.081329, 2.063812, 2.099213, 2.090363, 2.09668, 2.106049, 
    2.141144, 2.170563, 2.224731, 2.278564, 2.314606, 2.389587, 2.422333, 
    2.453766, 2.382721, 2.317963, 2.277863, 2.300446, 3.309052, 3.552643, 
    3.249664, 3.197845, 3.337128, 3.595245, 3.467255, 3.140778, 2.935089, 
    2.89447, 2.837311, 2.665558, 2.20575, 2.24707, 2.235779, 2.239258, 
    2.261261, 2.38092, 2.387299, 2.427734, 2.415833,
  2.401184, 2.398193, 2.423828, 3.309479, 3.072571, 2.76712, 2.796356, 
    2.581451, 2.810028, 2.245178, 2.527161, 4.033691, 2.381226, 2.2229, 
    2.385468, 2.475769, 2.552826, 2.562073, 2.590851, 2.595612, 2.598846, 
    2.634674, 2.644043, 2.62561, 2.534424, 2.409943, 2.323608, 3.1409, 
    2.814911, 2.379669, 3.159271, 3.192841, 2.894653, 2.245697, 2.322357, 
    3.046356, 3.046051, 2.91922, 2.541138, 2.066559, 2.134918, 2.107727, 
    2.11911, 2.139282, 2.075287, 2.002533, 1.990692, 2.026886, 2.043365, 
    2.033386, 2.02121, 2.057739, 2.091339, 2.117889, 2.150543, 2.173706, 
    2.200531, 2.200134, 2.19162, 2.216095, 2.222778, 2.248688, 2.268951, 
    2.272583, 2.305481, 2.309875, 2.32135, 2.329498, 2.297333, 2.249756, 
    2.195374, 2.104309, 2.019806, 1.952667, 2.076538, 3.058594, 3.25769, 
    2.96405, 2.803131, 2.863342, 2.890625, 3.529175, 3.669708, 2.780731, 
    2.712372, 2.238586, 2.131836, 2.31131, 2.363739, 2.364624, 2.357513, 
    2.375061, 2.456635, 2.456512, 2.447327, 2.407684,
  2.293365, 2.361481, 2.443359, 3.215576, 3.119659, 2.919922, 3.053528, 
    2.781372, 2.807892, 2.416748, 2.146545, 4.019562, 4.292999, 2.370636, 
    2.432892, 2.5896, 2.590149, 2.470917, 2.419037, 2.41272, 2.437988, 
    2.472412, 2.503937, 2.603546, 2.58902, 2.299316, 2.243774, 2.84552, 
    2.213257, 2.280487, 2.722443, 2.738922, 2.758972, 2.178925, 2.136719, 
    2.095978, 1.993164, 1.981262, 2.087982, 2.143188, 2.060883, 2.073181, 
    2.116974, 2.129303, 2.004669, 1.98111, 1.992401, 2.025574, 2.050568, 
    2.070374, 2.074219, 2.075043, 2.100067, 2.10318, 2.133209, 2.165222, 
    2.18927, 2.207764, 2.223907, 2.264191, 2.288544, 2.315125, 2.371368, 
    2.411072, 2.437653, 2.455475, 2.472534, 2.424103, 2.33783, 2.259094, 
    2.143494, 2.082794, 1.996613, 1.891937, 1.8685, 2.757263, 2.999603, 
    2.796021, 2.743896, 2.769989, 2.813477, 3.353424, 3.506226, 2.196869, 
    2.155212, 2.184052, 2.19043, 2.301453, 2.348572, 2.369141, 2.31366, 
    2.321747, 2.392517, 2.413208, 2.363129, 2.353516,
  2.757751, 2.495667, 2.760742, 2.9711, 3.090485, 2.983582, 3.033264, 
    3.159698, 3.098694, 2.743286, 2.808411, 3.727478, 4.262604, 2.524414, 
    2.508392, 2.667542, 2.598145, 2.520477, 2.517761, 2.552582, 2.54953, 
    2.597076, 2.652557, 2.684662, 2.615601, 2.33252, 2.834839, 2.432495, 
    2.126312, 2.220032, 2.183228, 2.613129, 2.126801, 2.208008, 2.131531, 
    2.091431, 2.072601, 2.151123, 2.248718, 2.206543, 2.161682, 2.137329, 
    2.102386, 2.131104, 2.146423, 2.169464, 2.154755, 2.184174, 2.203247, 
    2.20285, 2.217163, 2.191071, 2.191284, 2.155731, 2.119385, 2.101898, 
    2.068207, 2.040802, 2.033783, 2.030731, 2.046539, 2.074341, 2.124725, 
    2.155457, 2.181183, 2.291748, 2.366943, 2.397797, 2.349213, 2.284698, 
    2.300323, 2.317047, 2.157166, 1.982941, 1.991089, 2.903259, 2.957733, 
    3.19223, 3.408936, 3.541809, 3.295349, 3.042725, 2.444977, 2.033722, 
    2.123718, 2.150909, 2.259888, 2.322327, 2.377258, 2.385681, 2.312042, 
    2.324402, 2.287018, 2.368622, 2.868347, 2.941528,
  2.762634, 2.821472, 2.93515, 3.32605, 3.386383, 3.383026, 3.382019, 
    3.713226, 3.7742, 3.440948, 3.722137, 4.415436, 4.704712, 3.001007, 
    2.44754, 2.671997, 2.730255, 2.707977, 2.754395, 2.728088, 2.594971, 
    1.793854, 2.424011, 2.489075, 2.463959, 2.369629, 2.312866, 1.919678, 
    2.272736, 2.368805, 2.164215, 1.97998, 2.148804, 2.89975, 2.179749, 
    2.150421, 2.170654, 2.190582, 2.225983, 2.226868, 2.235077, 2.208466, 
    2.1586, 2.165161, 2.231201, 2.2677, 2.281158, 2.288025, 2.317841, 
    2.327209, 2.325134, 2.318085, 2.304016, 2.282562, 2.260468, 2.21875, 
    2.188934, 2.129639, 2.108856, 2.084045, 2.102539, 2.097443, 2.1026, 
    2.129822, 2.160522, 2.24472, 2.306122, 2.397827, 2.425354, 2.435364, 
    2.47348, 2.574738, 2.518311, 2.370758, 2.972717, 3.360687, 4.002014, 
    4.454224, 3.835236, 2.667542, 2.291779, 2.399658, 2.229095, 2.101501, 
    2.113159, 2.148102, 2.232147, 2.307312, 2.355469, 2.381317, 2.387695, 
    2.23761, 2.225891, 3.169464, 3.289124, 2.947723,
  2.709839, 2.911865, 2.983154, 3.779907, 4.368378, 4.797424, 4.493896, 
    4.718201, 5.032013, 5.549103, 5.336273, 4.350739, 5.118927, 3.993469, 
    2.67041, 2.583649, 2.772461, 2.831512, 2.88089, 2.889221, 3.060333, 
    2.17334, 2.257721, 2.565735, 2.445282, 2.362854, 2.424744, 2.447571, 
    2.174072, 2.407227, 2.277649, 2.129456, 2.102325, 3.05011, 2.145355, 
    2.162872, 2.126068, 2.185272, 2.257996, 2.259918, 2.291351, 2.260406, 
    2.283844, 2.306702, 2.353394, 2.396606, 2.425446, 2.410614, 2.403717, 
    2.402527, 2.393097, 2.385986, 2.375854, 2.342834, 2.326782, 2.305939, 
    2.274719, 2.203217, 2.169342, 2.176361, 2.184387, 2.181305, 2.201508, 
    2.21756, 2.20462, 2.20871, 2.210602, 2.289459, 2.447693, 2.523804, 
    2.441895, 2.583557, 3.510345, 3.169678, 2.285156, 2.248779, 2.256287, 
    2.16217, 2.153015, 2.216614, 2.16098, 2.153381, 2.072601, 2.065338, 
    2.067108, 2.11264, 2.125702, 2.203705, 2.235413, 2.355469, 2.38385, 
    2.405212, 3.799622, 4.610565, 3.900116, 2.940704,
  4.205109, 4.361969, 4.200806, 4.246582, 3.907471, 3.814728, 3.940765, 
    4.11911, 4.031982, 4.123352, 4.082703, 4.883301, 5.23407, 4.541138, 
    3.911163, 2.61438, 2.587646, 2.650696, 2.775848, 2.762299, 3.579987, 
    3.048126, 2.091766, 2.456421, 2.474823, 2.413025, 2.901855, 2.301727, 
    1.511169, 1.987305, 2.081116, 2.192017, 2.039642, 2.070526, 2.168884, 
    2.211853, 2.186005, 2.197723, 2.230255, 2.206329, 2.190948, 2.162781, 
    2.173431, 2.165192, 2.204834, 2.249939, 2.297638, 2.351379, 2.405273, 
    2.394867, 2.402588, 2.396729, 2.355804, 2.314331, 2.288544, 2.240387, 
    2.167053, 2.111969, 2.037292, 2.017761, 2.067261, 2.147583, 2.206055, 
    2.209839, 2.097412, 1.923248, 1.756592, 1.973053, 2.556061, 3.185425, 
    2.914063, 3.411591, 3.755981, 2.159637, 2.339661, 2.264832, 2.15799, 
    2.160492, 2.111328, 2.079224, 2.050049, 2.028381, 2.015625, 2.024292, 
    2.02713, 2.035095, 2.015167, 2.03952, 2.023834, 2.174347, 2.311584, 
    2.559631, 4.553741, 4.920166, 4.182129, 3.926025,
  4.821564, 4.93454, 4.913116, 4.823273, 4.571625, 4.187164, 3.854187, 
    3.800354, 3.725861, 3.234985, 2.339233, 4.613525, 5.06424, 4.829926, 
    4.429993, 3.682861, 2.71167, 2.625122, 2.805817, 2.696625, 3.926056, 
    3.695557, 1.899506, 1.742279, 2.440765, 2.89856, 3.196899, 2.351837, 
    1.874542, 2.450684, 2.080597, 2.254028, 2.131439, 2.144653, 2.15625, 
    2.144958, 2.15744, 2.13559, 2.179169, 2.193573, 2.140533, 2.071686, 
    2.079437, 2.055267, 1.990967, 2.049744, 2.076294, 2.095367, 2.147736, 
    2.145782, 2.1745, 2.145782, 2.124664, 2.106995, 2.08609, 1.999664, 
    1.933441, 1.872711, 1.761475, 1.697601, 1.675995, 1.706268, 1.766876, 
    1.846558, 1.749207, 1.489807, 1.285553, 1.983124, 4.376221, 3.638672, 
    3.109253, 4.134247, 3.718323, 2.158325, 2.310272, 2.247253, 2.13562, 
    2.053772, 2.013733, 1.981293, 1.966949, 1.963867, 1.964691, 1.944275, 
    1.886322, 1.88269, 1.849792, 1.816132, 1.748138, 1.781128, 1.933472, 
    2.354126, 4.110321, 4.801208, 4.630646, 4.781555,
  4.854004, 5.059723, 4.685242, 4.465424, 3.956787, 3.540619, 3.424347, 
    3.368439, 3.436951, 3.399261, 2.333466, 4.564331, 4.975098, 4.870087, 
    5.076202, 4.341705, 2.966156, 2.83963, 3.802002, 4.253082, 4.304352, 
    3.856476, 2.990204, 2.892151, 2.192291, 2.22644, 2.799896, 2.754486, 
    2.482666, 2.526031, 2.707184, 3.420654, 2.291656, 2.134674, 2.082611, 
    2.114899, 2.213013, 2.150299, 2.119415, 2.144257, 2.165253, 2.141327, 
    2.046539, 2.006378, 1.915558, 1.86322, 1.889008, 1.894135, 1.937195, 
    1.988495, 2.035339, 2.033783, 2.000061, 1.9487, 1.926636, 1.898102, 
    1.856659, 1.853851, 1.763672, 1.655457, 1.56842, 1.56723, 1.650726, 
    1.745911, 1.623657, 1.444397, 1.661926, 2.771118, 4.876099, 3.948029, 
    3.054626, 2.558594, 2.253906, 2.196594, 2.250793, 2.040436, 1.977081, 
    2.020905, 2.230713, 2.246826, 2.162811, 2.14212, 2.114502, 2.106049, 
    2.103516, 2.075989, 2.014832, 1.955139, 1.862, 1.802734, 1.745697, 
    1.923462, 3.127869, 4.165131, 4.602112, 4.752075,
  4.721954, 4.653503, 4.224976, 3.914215, 3.246155, 2.936127, 3.401947, 
    3.273865, 2.938934, 3.492188, 3.88739, 4.203247, 4.646515, 4.980316, 
    5.206604, 5.223297, 4.976593, 4.801666, 4.852173, 4.951904, 4.409485, 
    3.80838, 3.442047, 3.90332, 3.343048, 2.737885, 2.565887, 2.564056, 
    2.454498, 2.549072, 2.730804, 2.813416, 2.730743, 2.262238, 2.215118, 
    2.161316, 2.164001, 2.203369, 2.289764, 2.273041, 2.275787, 2.276215, 
    2.233673, 2.14679, 2.070068, 1.997864, 1.937958, 1.887299, 1.846741, 
    1.847839, 1.896637, 1.925659, 1.938995, 1.879211, 1.882294, 1.897797, 
    1.832275, 1.799744, 1.732574, 1.705353, 1.654022, 1.613617, 1.622528, 
    1.604492, 1.510376, 1.792633, 2.786285, 3.147919, 3.691132, 3.351746, 
    2.450623, 2.575806, 2.590759, 2.707275, 3.16861, 2.101898, 2.024017, 
    2.088654, 2.165436, 2.141022, 2.129822, 2.187347, 2.23645, 2.264862, 
    2.296356, 2.295319, 2.260742, 2.202545, 2.066864, 1.969208, 1.773773, 
    1.676208, 2.029358, 3.346344, 4.602814, 4.792114,
  4.936188, 4.744202, 4.193237, 3.339844, 2.676941, 2.25528, 2.828125, 
    2.864502, 2.253723, 3.200256, 4.068207, 4.027496, 4.178833, 4.719482, 
    5.228912, 5.340363, 5.588043, 5.941345, 5.234833, 4.833221, 4.492798, 
    5.778961, 5.464508, 2.00473, 2.46347, 2.3797, 2.394135, 3.032288, 
    2.88269, 3.293671, 3.235809, 2.892517, 2.756195, 2.045959, 2.272461, 
    2.268036, 2.222595, 2.214233, 2.19635, 2.206573, 2.217957, 2.188171, 
    2.216431, 2.184235, 2.156067, 2.178314, 2.125854, 2.107361, 2.028412, 
    1.959442, 1.973572, 1.953705, 1.961487, 1.953186, 1.930145, 1.929565, 
    1.882629, 1.822876, 1.732758, 1.699921, 1.688629, 1.615295, 1.528839, 
    1.508911, 1.78186, 2.822174, 3.37851, 3.953857, 3.882874, 2.897705, 
    2.480591, 3.100586, 3.276764, 3.329651, 3.242737, 2.316803, 2.067566, 
    2.019287, 2.042755, 2.038879, 1.988617, 1.906952, 1.864899, 1.918091, 
    2.040619, 2.154877, 2.218506, 2.226501, 2.208984, 2.184387, 2.082855, 
    1.870392, 1.800323, 2.2995, 4.433594, 5.167847,
  5.297577, 5.055023, 4.308197, 2.532074, 2.10672, 2.083679, 2.254303, 
    2.348175, 2.445953, 2.624268, 3.906708, 4.179291, 4.927277, 5.193878, 
    5.66095, 5.133026, 5.332031, 5.706879, 5.362091, 5.95047, 5.501221, 
    5.014587, 3.644318, 1.745636, 2.729614, 1.356323, 1.945709, 2.856049, 
    3.608643, 4.296539, 4.029236, 3.16864, 2.859985, 2.227234, 2.937225, 
    2.697449, 3.015961, 3.19519, 2.500793, 2.323395, 2.324738, 2.284515, 
    2.32135, 2.328125, 2.300781, 2.298248, 2.305939, 2.34668, 2.304871, 
    2.230164, 2.182404, 2.070892, 1.983124, 1.925446, 1.91217, 1.941345, 
    1.920319, 1.812103, 1.671875, 1.584442, 1.5578, 1.554291, 1.525269, 
    1.73172, 3.173767, 3.780151, 3.961243, 4.515045, 4.717529, 3.963806, 
    3.18866, 3.103455, 3.148956, 3.417053, 3.413788, 3.300995, 2.609955, 
    2.266724, 1.989563, 1.918365, 1.92804, 1.914886, 1.79657, 1.603973, 
    1.434052, 1.393677, 1.596497, 1.749298, 1.821411, 1.963806, 2.098938, 
    2.032623, 1.869324, 1.963867, 2.688629, 5.265411,
  4.178772, 2.352417, 2.225586, 2.203827, 2.103973, 2.169342, 2.873444, 
    3.297058, 2.51944, 2.55188, 2.888947, 3.375, 3.810425, 3.509247, 
    2.717896, 4.550598, 5.02597, 4.509247, 4.839905, 5.438477, 4.950134, 
    3.61145, 3.14212, 3.038727, 2.898376, 2.533905, 2.44751, 3.080444, 
    3.729675, 3.878082, 3.839172, 3.801758, 3.577087, 3.601288, 3.656525, 
    2.727539, 2.611176, 3.070007, 2.75351, 2.684235, 2.710938, 2.656189, 
    2.675323, 2.723755, 2.68222, 2.580414, 2.511841, 2.548065, 2.530609, 
    2.466614, 2.408783, 2.308716, 2.188599, 2.074219, 1.992645, 1.963806, 
    1.933594, 1.83667, 1.688019, 1.571167, 1.518799, 1.511475, 1.531982, 
    2.157928, 2.952148, 3.467438, 3.604431, 4.484497, 4.921234, 4.254486, 
    3.753845, 3.324921, 3.371735, 3.644135, 3.712494, 3.755463, 3.730469, 
    3.109772, 2.587158, 2.340363, 2.28418, 2.145508, 1.867767, 1.37915, 
    0.7700806, 0.3293152, 0.5402527, 0.9640503, 1.201904, 1.441559, 1.729828, 
    1.891663, 1.988098, 2.26767, 3.875854, 4.477478,
  2.708923, 2.095886, 2.210785, 2.802734, 2.320435, 2.19223, 2.481964, 
    2.564453, 2.389862, 2.283386, 2.530334, 2.942474, 2.922668, 2.537811, 
    3.095032, 3.594788, 3.887817, 3.537445, 3.707275, 4.068817, 3.755798, 
    3.243866, 3.278137, 3.451965, 3.202606, 3.358398, 3.475464, 3.211548, 
    3.32901, 3.362915, 3.270203, 3.291931, 3.265472, 3.49585, 3.579895, 
    3.240234, 2.630341, 2.614594, 3.122772, 3.613281, 3.578522, 3.152161, 
    2.853973, 2.743286, 2.601624, 2.475922, 2.444153, 2.419312, 2.413483, 
    2.436188, 2.412689, 2.323181, 2.222137, 2.123688, 2.02356, 1.932892, 
    1.811462, 1.68335, 1.58905, 1.513153, 1.490997, 1.528442, 1.552917, 
    1.815491, 2.035278, 2.387939, 2.85553, 3.439575, 4.014008, 4.239197, 
    4.316284, 3.864929, 3.869934, 4.127014, 3.738403, 4.096985, 4.247223, 
    4.138672, 4.206177, 3.684357, 2.752014, 2.364197, 2.047546, 1.510284, 
    1.004517, 0.7933655, 0.7317505, 0.7012634, 0.5831604, 0.8701172, 
    1.296661, 1.5401, 1.748383, 2.038086, 3.038757, 3.429291,
  2.274994, 2.10025, 2.601746, 2.868164, 2.269592, 2.40274, 2.449554, 
    2.617706, 2.424011, 2.295258, 1.876831, 2.143036, 2.498962, 2.472717, 
    2.272522, 2.641418, 2.930847, 2.843384, 3.237427, 3.641724, 3.581909, 
    3.402679, 2.95639, 2.8349, 2.75824, 2.361542, 2.070068, 2.421143, 
    2.906464, 3.017578, 2.919739, 2.530396, 2.761444, 2.901611, 2.990753, 
    2.602875, 2.557434, 2.531342, 2.926056, 2.51712, 2.596741, 2.417206, 
    2.348755, 2.357666, 2.303375, 2.23465, 2.232147, 2.267334, 2.284485, 
    2.293701, 2.291534, 2.287964, 2.243408, 2.121613, 2.002533, 1.895508, 
    1.7724, 1.661652, 1.651733, 1.702606, 1.709625, 1.636841, 1.607544, 
    1.578125, 1.847076, 2.508942, 3.08667, 3.650269, 3.818634, 4.001251, 
    4.058777, 4.217041, 4.30838, 3.470978, 4.305786, 4.671021, 4.830933, 
    4.606567, 4.228638, 3.932678, 3.231171, 2.309753, 1.975586, 1.601501, 
    1.202942, 1.020844, 0.8374329, 0.5549011, 0.1708984, 0.2122498, 
    0.8414001, 1.362701, 1.680878, 1.859375, 2.07251, 2.537781,
  1.948914, 1.858521, 1.835052, 2.009369, 2.253601, 2.253784, 2.295898, 
    2.420837, 2.604156, 2.772736, 2.801025, 2.5737, 2.941345, 3.16687, 
    3.007233, 3.309692, 3.459839, 3.383209, 3.535614, 3.825745, 3.438934, 
    3.424072, 3.034882, 2.232422, 1.900299, 1.735413, 1.641327, 1.735107, 
    2.032349, 2.072906, 1.809753, 1.750305, 1.885437, 2.050049, 1.995117, 
    1.899078, 2.065704, 2.059509, 1.93985, 2.311462, 2.908783, 2.699615, 
    2.469788, 2.384399, 2.373322, 2.289124, 2.254517, 2.257874, 2.235504, 
    2.170654, 2.160004, 2.204041, 2.229614, 2.193665, 2.135498, 2.036255, 
    1.892639, 1.796692, 1.741211, 1.709747, 1.674866, 1.757416, 1.723633, 
    2.490112, 3.104858, 2.540039, 2.892639, 2.801758, 2.996094, 3.461609, 
    3.846008, 3.908661, 4.020508, 4.123779, 4.294861, 4.160553, 3.707855, 
    3.29538, 3.159271, 2.835297, 2.68576, 2.343689, 1.985535, 2.111176, 
    1.72168, 1.067505, 0.3016968, -0.3977051, -0.7251587, -0.5596313, 
    0.1753845, 0.961792, 1.48999, 1.699402, 1.733002, 1.795685,
  1.891022, 1.7323, 1.850311, 2.242004, 2.387482, 2.434814, 2.234924, 
    2.557739, 3.153717, 3.278839, 3.280334, 3.194, 3.269287, 3.15033, 
    2.895905, 2.539642, 2.365784, 2.040558, 2.044769, 2.245636, 2.357758, 
    2.538544, 2.4599, 2.308136, 2.179474, 1.904907, 1.857971, 1.726379, 
    1.71402, 1.918945, 2.606445, 2.486664, 2.026581, 1.651489, 1.834442, 
    1.856567, 1.74173, 1.95575, 1.994141, 2.145172, 2.859955, 2.817902, 
    2.547058, 2.138336, 2.360229, 2.301971, 2.241547, 2.159698, 2.127808, 
    2.194733, 2.361023, 2.575775, 2.642426, 2.505157, 2.400116, 2.280914, 
    2.131958, 2.028778, 1.965942, 1.898621, 1.774323, 1.902527, 2.770813, 
    2.795959, 2.560181, 2.152405, 2.270508, 2.341095, 2.57312, 2.776123, 
    2.999146, 3.060486, 3.245361, 3.058197, 3.015503, 2.370636, 3.291382, 
    3.073578, 2.741669, 2.402069, 2.227539, 1.468994, 1.567169, 1.417389, 
    1.07251, 1.005737, 0.4856873, -0.3548279, -0.9366455, -0.7978516, 
    -0.03573608, 0.8084717, 1.34552, 1.527985, 1.639709, 1.734161,
  1.323242, 1.474792, 1.480255, 2.034576, 2.226044, 2.345886, 1.885559, 
    2.508392, 2.858582, 3.197388, 2.921814, 2.505402, 2.396881, 2.381256, 
    2.089203, 1.776611, 1.532623, 1.668213, 1.745422, 1.73172, 1.850525, 
    1.930939, 2.122864, 2.069214, 1.894897, 1.814301, 1.753296, 1.788025, 
    1.639191, 1.745178, 2.05423, 2.370483, 2.03125, 1.91452, 1.952454, 
    1.949371, 1.929688, 2.130554, 2.084106, 1.570435, 1.489563, 1.324341, 
    1.812439, 2.013092, 1.865631, 2.288544, 2.593933, 2.905396, 3.238281, 
    3.447906, 3.593872, 3.290375, 2.781006, 2.543945, 1.986237, 2.100128, 
    2.10202, 2.085999, 2.005005, 1.91095, 2.531891, 3.715546, 2.327148, 
    2.174347, 2.070496, 2.224945, 2.175262, 2.195068, 2.416687, 2.744141, 
    2.645508, 2.961578, 2.718689, 2.888092, 2.785858, 2.780731, 3.757294, 
    3.772858, 3.310852, 2.775513, 1.680511, 1.471497, 0.7423096, -0.1021423, 
    -0.1689453, 0.6904907, 1.031006, 0.6725769, 0.2465515, 0.2412109, 
    0.5283203, 0.8944702, 1.185303, 1.317841, 1.364258, 1.50116,
  0.7744141, 0.8408203, 1.636841, 2.12439, 1.780853, 1.155975, 1.849487, 
    1.846588, 2.116394, 2.390869, 2.480988, 2.294128, 2.000305, 1.746613, 
    1.681702, 1.766418, 1.996552, 2.280792, 2.30722, 2.416595, 2.186646, 
    2.212494, 2.300507, 2.252228, 1.951813, 1.875092, 1.775635, 1.779083, 
    1.571808, 1.294067, 1.101624, 0.9819641, 1.102081, 1.071045, 1.04245, 
    1.216339, 1.533905, 2.011963, 1.807922, 1.216522, 0.9392395, 1.386536, 
    1.55011, 1.317688, 1.481445, 1.612885, 2.03302, 2.617828, 2.57785, 
    2.573425, 2.473785, 2.175781, 1.992493, 1.708191, 1.572205, 1.895142, 
    2.229828, 1.981842, 2.062805, 1.960938, 1.933929, 2.010468, 2.244751, 
    2.129608, 2.214905, 2.260193, 2.225891, 2.407867, 2.822266, 3.019012, 
    3.159485, 2.574646, 2.972839, 3.047211, 3.019287, 2.974854, 3.68927, 
    3.3078, 2.510529, 2.212677, 1.637817, 1.201569, 0.6065979, 0.1448059, 
    0.1952515, 0.1580505, 0.366272, 0.7109985, 0.9625549, 1.13028, 1.181396, 
    0.7828064, 0.1383972, 0.190094, 0.6260376, 0.7960815,
  0.3725281, 0.4692688, 0.5335388, 1.440063, 1.731049, 1.86441, 0.8770142, 
    2.065887, 2.143219, 2.320587, 2.428986, 2.486206, 2.348969, 2.307098, 
    2.540039, 2.73764, 3.228912, 3.4505, 3.661591, 3.543365, 3.478699, 
    3.279602, 2.804565, 2.589844, 2.502686, 2.308136, 2.197632, 2.128326, 
    2.029083, 1.384125, 1.348328, 1.180023, 0.9821472, 1.100922, 1.120514, 
    1.275909, 2.206116, 1.922333, 1.842499, 1.496613, 0.8390198, 1.269775, 
    1.365875, 1.425842, 1.340942, 1.362488, 1.282867, 1.345642, 1.322998, 
    1.134888, 1.387299, 1.029877, 1.536652, 1.357422, 1.304352, 1.279755, 
    1.370178, 1.622437, 1.913666, 2.198242, 2.18335, 2.178986, 1.86792, 
    2.055725, 2.160614, 2.465729, 3.043945, 3.523834, 3.819061, 4.041351, 
    4.037048, 3.624878, 3.383942, 3.26004, 2.915161, 2.788452, 2.643768, 
    3.118591, 2.908142, 2.523163, 1.776245, 1.183014, 0.9584656, 1.320435, 
    1.349945, 1.346802, 1.096161, 0.4152527, 0.5882263, 1.306854, 1.677063, 
    1.805939, 1.14856, 0.1846924, -0.1242065, 0.02584839,
  0.5375671, 0.3875122, 0.3937378, 0.115448, -0.2626343, 1.809052, 2.262482, 
    2.421997, 2.62265, 2.614441, 3.009186, 2.773834, 2.74942, 2.599487, 
    3.281586, 3.435364, 3.663086, 3.838684, 3.876495, 3.728333, 3.516266, 
    3.193817, 2.938873, 2.669006, 2.489349, 2.573883, 2.46048, 2.294708, 
    2.159973, 2.051483, 1.948517, 1.602478, 1.410675, 1.313812, 1.818024, 
    1.687958, 1.148895, 1.404114, 0.6616516, 0.7895813, 0.4679565, 0.6096191, 
    0.6869812, 0.6767578, 1.406067, 1.544189, 1.634888, 1.715485, 1.584534, 
    1.259827, 1.38266, 1.494598, 1.503113, 1.834839, 1.933807, 2.119141, 
    2.190033, 2.452606, 3.012634, 2.816132, 3.034241, 3.168884, 3.359222, 
    3.628845, 4.24649, 4.269867, 4.329803, 4.13269, 4.040558, 3.258514, 
    3.840637, 3.851624, 3.761902, 3.105591, 3.777863, 3.07663, 3.362183, 
    3.078339, 2.977753, 2.419128, 2.034576, 1.68866, 2.15213, 2.505737, 
    2.676895, 2.413132, 2.308105, 2.383789, 2.685547, 2.971741, 2.465179, 
    2.343018, 2.297607, 1.5961, 1.24588, 0.8505859,
  1.906708, 1.356445, 0.8496704, 0.6033325, 0.4563904, 0.9065857, 1.760895, 
    2.457428, 2.805725, 3.203278, 3.496307, 3.782623, 3.634644, 3.446564, 
    3.174438, 3.837616, 3.358582, 3.332672, 3.198547, 3.635223, 3.639465, 
    3.553314, 3.439789, 3.188629, 2.927032, 2.858276, 2.883453, 2.712555, 
    2.714783, 2.287018, 2.133636, 2.074677, 2.075317, 1.938995, 1.473175, 
    1.376221, 1.415283, 1.394531, 1.693237, 1.649689, 1.327271, 1.296082, 
    1.263672, 1.216736, 1.173889, 1.092712, 1.063873, 1.145813, 1.3078, 
    1.556854, 1.82254, 2.098114, 2.312866, 2.517181, 2.705536, 2.806335, 
    2.914459, 3.002411, 3.079956, 3.054169, 3.029633, 2.962158, 2.789886, 
    4.062286, 3.920502, 4.163666, 4.308716, 3.823242, 3.71225, 2.873047, 
    3.332703, 3.468872, 3.036987, 3.867188, 3.992889, 3.915436, 3.589508, 
    3.010345, 2.820923, 2.732117, 2.575928, 3.25415, 3.053314, 3.33876, 
    3.379349, 3.187119, 2.771881, 2.742569, 3.1745, 3.555328, 3.588989, 
    3.097534, 3.187164, 2.933533, 2.673767, 2.196564,
  3.038147, 2.66217, 2.348053, 2.514069, 2.816986, 3.178894, 3.774017, 
    3.835358, 3.872589, 3.711334, 3.658478, 3.544189, 3.424164, 3.258179, 
    3.127075, 3.108978, 3.097412, 3.060608, 3.024597, 3.054504, 3.078217, 
    3.020874, 2.928558, 2.746613, 2.479156, 3.340942, 3.249786, 2.940643, 
    3.00235, 2.949615, 2.754028, 2.474731, 2.359375, 2.252869, 2.124939, 
    2.019135, 1.995331, 1.965485, 1.941467, 1.841339, 1.754486, 1.626709, 
    1.496399, 1.390289, 1.357513, 1.379425, 1.435242, 1.595642, 1.831665, 
    2.089142, 2.355072, 2.601318, 2.817719, 2.987244, 3.12973, 3.278442, 
    3.431305, 3.574341, 3.707031, 3.837311, 3.963562, 4.124207, 4.2435, 
    4.294464, 4.219788, 4.216675, 4.043884, 3.855927, 3.750458, 3.899658, 
    3.766327, 3.668335, 3.639923, 3.923889, 4.0177, 3.377533, 3.326172, 
    3.338074, 3.919983, 3.809906, 3.705383, 3.666519, 3.749435, 3.848373, 
    3.898956, 3.914383, 3.808136, 3.70108, 3.844254, 4.071243, 4.284241, 
    4.260345, 3.976715, 3.989838, 3.889313, 3.739044,
  4.058807, 3.955322, 3.91571, 3.810547, 4.236267, 4.338806, 4.426697, 
    4.110413, 4.019714, 3.922729, 3.811523, 3.67395, 3.576019, 3.479736, 
    3.439789, 3.410492, 3.438293, 3.46875, 3.527496, 3.609436, 3.641663, 
    3.673889, 3.652924, 3.476624, 3.207489, 3.966461, 3.908478, 3.258118, 
    3.164001, 3.044281, 2.837036, 2.635345, 2.511841, 2.400513, 2.251495, 
    2.159576, 2.047852, 1.980347, 1.916931, 1.895813, 1.849091, 1.840607, 
    1.848175, 1.845245, 1.849213, 1.896149, 1.983856, 2.099945, 2.156494, 
    2.222382, 2.306976, 2.407837, 2.469818, 2.493835, 2.568573, 2.687622, 
    2.808197, 2.975433, 3.127472, 3.304688, 3.415771, 3.537628, 3.602081, 
    3.591461, 3.608398, 3.563293, 3.517914, 3.494324, 3.482513, 3.513672, 
    3.548187, 3.908539, 3.81427, 4.274536, 4.331192, 4.310913, 4.229797, 
    4.14592, 4.012192, 3.908173, 3.875427, 3.861832, 3.918274, 4.035721, 
    4.111832, 4.2061, 4.195877, 4.176651, 4.251129, 4.39978, 4.52536, 
    4.547089, 4.123108, 4.064789, 4.010529, 4.036255,
  3.834839, 3.717194, 3.656982, 3.570251, 3.438293, 3.329376, 3.232483, 
    3.1427, 3.068298, 2.996735, 2.932281, 2.888611, 2.85202, 2.840942, 
    2.908997, 2.974457, 3.023895, 3.096619, 3.130005, 3.151245, 3.184448, 
    3.188538, 3.152679, 3.122009, 3.082947, 3.012329, 2.998291, 2.941345, 
    2.848572, 2.805725, 2.708008, 2.606903, 2.53299, 2.439972, 2.343231, 
    2.277588, 2.252472, 2.248444, 2.22879, 2.228973, 2.237457, 2.256256, 
    2.270447, 2.306885, 2.362305, 2.429352, 2.480225, 2.569244, 2.626282, 
    2.684113, 2.763275, 2.846161, 2.955475, 3.072205, 3.177856, 3.268494, 
    3.362183, 3.440247, 3.51535, 3.577667, 3.626617, 3.68399, 3.745758, 
    3.783203, 3.763977, 3.746094, 3.731384, 3.730225, 3.736267, 3.735077, 
    3.77533, 3.800018, 3.84845, 3.870483, 3.892853, 3.916534, 3.944855, 
    3.928009, 3.942413, 3.944611, 3.939758, 3.956421, 4.030579, 4.034668, 
    4.058258, 4.096588, 4.11441, 4.091034, 4.072876, 4.099213, 4.054108, 
    4.062836, 4.08432, 3.987579, 3.935547, 3.910858,
  3.682159, 3.683289, 3.673248, 3.637024, 3.621552, 3.611481, 3.596283, 
    3.569855, 3.557892, 3.545563, 3.535492, 3.528107, 3.527679, 3.524017, 
    3.509705, 3.480408, 3.479279, 3.452454, 3.433868, 3.423706, 3.413208, 
    3.401886, 3.381897, 3.33374, 3.312897, 3.300262, 3.306641, 3.284088, 
    3.27655, 3.25293, 3.233398, 3.210419, 3.183777, 3.136261, 3.098999, 
    3.07309, 3.007477, 2.974335, 2.955414, 2.913208, 2.884644, 2.857422, 
    2.827728, 2.814514, 2.788666, 2.753326, 2.736389, 2.716156, 2.701172, 
    2.691132, 2.69812, 2.696014, 2.732208, 2.759186, 2.801971, 2.832367, 
    2.869812, 2.903503, 2.950134, 2.96701, 2.995056, 3.021851, 3.020508, 
    3.032928, 3.05188, 3.066986, 3.073181, 3.080414, 3.097046, 3.118561, 
    3.158569, 3.1875, 3.198425, 3.208252, 3.220581, 3.238861, 3.24527, 
    3.249817, 3.268036, 3.282959, 3.318115, 3.348511, 3.393097, 3.444977, 
    3.499725, 3.540497, 3.566986, 3.585785, 3.619812, 3.66626, 3.70047, 
    3.710999, 3.717499, 3.712952, 3.70816, 3.686859,
  2.725204, 2.763428, 2.805161, 2.850479, 2.895981, 2.944611, 2.997604, 
    3.047348, 3.100723, 3.155228, 3.210831, 3.261673, 3.306259, 3.342911, 
    3.369156, 3.38028, 3.374832, 3.348785, 3.305557, 3.25145, 3.185425, 
    3.111145, 3.036407, 2.959259, 2.877487, 2.798523, 2.719543, 2.641495, 
    2.564529, 2.491623, 2.428802, 2.374435, 2.328857, 2.29454, 2.270065, 
    2.250153, 2.237183, 2.229843, 2.228729, 2.235428, 2.248657, 2.265442, 
    2.286865, 2.309982, 2.333801, 2.353729, 2.382111, 2.40126, 2.42984, 
    2.452103, 2.4758, 2.493698, 2.47345, 2.450211, 2.487396, 2.445923, 
    2.403854, 2.418839, 2.436676, 2.373962, 2.322601, 2.390656, 2.386414, 
    2.438965, 2.485321, 2.526459, 2.573334, 2.605682, 2.639267, 2.686676, 
    2.711304, 2.718658, 2.710831, 2.945007, 2.807373, 2.801056, 2.850922, 
    2.948441, 2.804565, 2.832306, 2.834778, 2.827225, 2.807571, 2.796234, 
    2.786682, 2.765259, 2.738815, 2.710495, 2.682434, 2.658615, 2.641357, 
    2.631592, 2.632965, 2.642853, 2.666107, 2.693192,
  3.781586, 3.886597, 3.936996, 3.958206, 3.942535, 3.889084, 3.808807, 
    3.720337, 3.644287, 3.594543, 3.576981, 3.588882, 3.64032, 3.733871, 
    3.835037, 3.933487, 3.985825, 3.993896, 3.914658, 3.776123, 3.582687, 
    3.374756, 3.164993, 2.989471, 2.848465, 2.744873, 2.675018, 2.624298, 
    2.586594, 2.54657, 2.500076, 2.451126, 2.398712, 2.349564, 2.306396, 
    2.273911, 2.265961, 2.286728, 2.333206, 2.398392, 2.47789, 2.607437, 
    2.745529, 2.865189, 3.008987, 3.185242, 3.289474, 3.434982, 3.59201, 
    3.761154, 3.881912, 3.961731, 4.037704, 4.076065, 4.131271, 4.109528, 
    4.112656, 4.128006, 4.081848, 4.031982, 3.93869, 3.805618, 3.671768, 
    3.536346, 3.434784, 3.361679, 3.383224, 3.509659, 3.672226, 3.915955, 
    4.030823, 4.114075, 4.164017, 4.165955, 4.015182, 3.909912, 3.877625, 
    3.896622, 4.004242, 3.844604, 3.863159, 3.92749, 3.701263, 3.681976, 
    3.606598, 3.564926, 3.362717, 3.269867, 3.209457, 3.182373, 3.177933, 
    3.212006, 3.286606, 3.391495, 3.509262, 3.64241,
  4.123978, 4.180023, 4.24762, 4.314728, 4.33316, 4.34343, 4.408936, 
    4.527634, 4.549042, 4.44519, 4.306396, 4.081589, 3.832245, 3.581268, 
    3.373978, 3.268707, 3.261795, 3.268967, 3.240631, 3.182236, 3.202042, 
    3.391937, 3.655151, 3.905685, 3.935699, 3.858215, 3.697159, 3.469864, 
    3.258881, 3.084641, 2.940842, 2.82338, 2.692917, 2.573914, 2.424042, 
    2.282562, 2.242264, 2.279846, 2.39122, 2.554642, 2.741486, 3.013428, 
    3.273514, 3.720978, 4.304565, 4.729889, 4.863235, 4.851913, 4.860703, 
    4.814667, 4.77626, 4.760315, 4.831268, 4.918518, 4.980423, 5.066483, 
    5.032959, 4.879898, 4.608353, 4.366425, 4.134644, 3.905685, 3.709198, 
    3.526505, 3.347549, 3.296967, 3.322998, 3.461212, 3.61615, 3.743835, 
    3.845001, 3.845139, 3.779373, 3.706528, 3.668823, 3.665771, 3.767258, 
    3.910492, 3.941162, 4.019485, 4.143112, 4.336548, 4.261871, 4.261856, 
    4.268768, 4.391541, 4.443375, 4.274048, 4.130737, 4.078003, 3.873779, 
    3.840897, 3.841614, 3.883087, 3.930878, 4.021622,
  4.229965, 4.309387, 4.185745, 4.004181, 3.82254, 3.680954, 3.602493, 
    3.452026, 3.302765, 3.175354, 3.120453, 3.106064, 3.112, 3.054581, 
    2.878723, 2.683029, 2.457764, 2.381393, 2.465897, 2.425659, 2.22319, 
    2.402222, 2.749817, 3.059448, 3.255432, 3.337585, 3.252625, 3.084717, 
    3.061081, 3.151199, 3.34494, 3.593445, 3.836929, 3.953857, 3.865051, 
    3.598328, 3.338882, 3.152802, 2.955933, 2.862198, 2.931656, 3.076843, 
    3.18602, 3.353073, 3.805878, 4.686539, 3.538498, 3.862656, 4.056, 
    4.264282, 4.479691, 4.624237, 4.798965, 4.925858, 4.831726, 4.759781, 
    4.391876, 4.41539, 4.220795, 4.068573, 4.039276, 4.075806, 4.052948, 
    3.850601, 3.556335, 3.246384, 3.178864, 3.213043, 3.305161, 3.387909, 
    3.439606, 3.525803, 3.590775, 3.72821, 3.927353, 4.205154, 4.425995, 
    4.616486, 4.685165, 4.691345, 4.812973, 4.91037, 4.873199, 4.84729, 
    4.860626, 4.845642, 4.998718, 5.332245, 5.385178, 4.712906, 4.170715, 
    3.796173, 3.638565, 3.645523, 3.810425, 4.071304,
  3.903534, 3.842133, 3.790955, 3.807632, 3.851456, 3.928009, 3.981918, 
    3.955154, 3.885498, 3.612518, 3.421494, 3.280548, 3.032303, 2.872604, 
    3.289139, 3.37027, 2.966095, 2.671432, 2.488831, 2.130173, 1.811737, 
    2.070068, 2.237457, 2.515259, 2.974045, 3.099884, 2.878143, 2.884262, 
    3.073578, 3.327759, 3.718307, 4.01088, 4.102493, 4.06955, 4.015701, 
    4.087189, 4.197342, 4.163025, 4.017212, 3.898788, 3.718384, 3.537323, 
    3.536087, 3.658401, 3.896881, 4.431656, 4.059448, 4.188751, 4.11174, 
    4.145523, 4.101379, 4.028412, 3.922745, 3.762115, 3.535492, 3.318054, 
    3.010941, 2.807114, 2.809326, 2.929047, 3.12085, 3.325211, 3.410248, 
    3.512772, 3.534637, 3.533157, 3.514008, 3.548187, 3.72818, 3.588608, 
    4.153458, 4.171936, 4.131897, 4.091736, 4.105667, 3.827026, 4.7491, 
    4.958618, 5.155487, 5.315704, 5.450333, 5.468811, 5.411133, 5.299744, 
    5.334396, 5.489914, 5.488174, 5.511551, 5.661606, 5.738556, 5.424637, 
    4.742844, 4.283096, 4.056015, 3.94931, 3.917191,
  7.14917, 5.934067, 6.030212, 5.453995, 4.934586, 4.531799, 4.431076, 
    4.653915, 4.974823, 5.17189, 5.347549, 5.000473, 4.469742, 3.962646, 
    3.379913, 2.934845, 2.371246, 2.094681, 2.056015, 2.147293, 1.880096, 
    1.695648, 1.734985, 1.85907, 1.97261, 2.170517, 2.412308, 2.681198, 
    2.86908, 2.898254, 2.824631, 2.773712, 2.862381, 3.034195, 3.19754, 
    3.174683, 3.006271, 2.83667, 2.790771, 2.741287, 2.761612, 2.856857, 
    3.11824, 3.451385, 3.129837, 3.105621, 3.16362, 2.998001, 2.746826, 
    2.438553, 2.175858, 1.946823, 1.806396, 1.705612, 1.647934, 1.662842, 
    1.749115, 1.903992, 2.153992, 2.463928, 2.752899, 3.061813, 3.428452, 
    3.760101, 4.078461, 4.376724, 4.561127, 4.705994, 4.920959, 5.088776, 
    5.350067, 5.301437, 5.332153, 5.313858, 5.288925, 5.074402, 4.846497, 
    4.72377, 5.491333, 5.797195, 6.241028, 6.329102, 6.291214, 6.104095, 
    6.065308, 6.078125, 6.235092, 6.372391, 6.410233, 6.367844, 6.269928, 
    6.156326, 6.210556, 6.346375, 6.622421, 7.012253,
  11.90143, 12.22017, 12.14725, 11.57364, 10.95683, 10.41968, 9.807556, 
    9.293716, 9.171692, 9.590378, 10.06354, 9.90892, 8.827881, 7.239136, 
    5.770142, 4.595917, 4.033157, 3.865768, 3.86499, 3.890121, 3.961212, 
    3.921555, 3.833801, 3.728134, 3.592072, 3.330933, 3.106659, 2.998703, 
    3.054306, 3.104126, 3.033081, 2.645264, 2.282562, 3.224503, 3.295013, 
    3.576965, 3.394424, 3.109711, 2.698761, 2.414703, 2.239777, 2.11348, 
    1.984833, 1.868042, 1.716583, 1.389832, 0.8083801, -0.02389526, 
    -0.8984375, -1.352814, -1.433685, -1.221344, -0.8445435, -0.4090271, 
    -0.3188782, -0.0730896, 0.7341003, 1.488983, 1.957031, 2.385803, 
    2.569244, 2.929779, 3.437958, 3.802734, 3.879944, 3.781708, 3.699738, 
    3.744965, 3.818115, 3.84314, 3.98465, 4.604156, 5.217438, 5.865234, 
    6.480774, 6.973297, 7.198242, 7.274628, 7.678894, 8.20639, 7.695557, 
    7.352219, 6.933792, 6.602463, 6.462387, 6.527802, 6.612366, 6.727875, 
    6.859497, 7.065353, 7.316864, 7.664993, 8.240768, 9.09993, 10.13002, 
    11.08058,
  11.22937, 11.26746, 11.09662, 10.81335, 10.53592, 10.16559, 9.627289, 
    9.159698, 8.872406, 8.67749, 8.456787, 8.382233, 8.470306, 8.891602, 
    9.366394, 10.03809, 10.44479, 10.6528, 10.49207, 9.63562, 8.80246, 
    8.357162, 7.993622, 7.746735, 7.430603, 6.545258, 5.557892, 4.577026, 
    3.922058, 3.324158, 2.517456, 1.761047, 1.305847, 1.016479, 1.061981, 
    1.219025, 1.629944, 1.601013, 1.540649, 1.601685, 2.018951, 2.359772, 
    2.1297, 1.70224, 1.387238, 1.021667, 0.4837952, -0.08731079, -0.3934326, 
    -0.493866, -0.5217285, -0.5289917, -0.5177917, -0.4451904, -0.3433533, 
    -0.2729187, 0.1400452, 0.4781189, 0.6233215, 0.8130188, 0.9058838, 
    0.9534607, 1.023071, 1.186005, 1.349945, 1.511658, 1.702759, 1.899109, 
    2.039917, 2.119354, 2.191071, 2.308868, 2.446655, 2.551361, 2.672119, 
    2.762756, 2.763733, 2.688599, 2.744293, 3.13269, 4.734528, 6.094269, 
    6.350708, 6.459503, 6.920502, 7.30545, 7.811401, 8.140625, 8.408325, 
    8.61203, 8.694031, 8.838623, 9.138275, 9.627289, 10.22839, 10.82922,
  5.544403, 5.312958, 4.866211, 4.456635, 4.161987, 3.721375, 3.275269, 
    2.792847, 2.52597, 2.451202, 2.431732, 2.490448, 2.556915, 2.66037, 
    2.755096, 2.881287, 3.032654, 3.245331, 3.555634, 3.907104, 4.225555, 
    3.960052, 3.381775, 2.882233, 2.597595, 2.363739, 2.102051, 1.908783, 
    1.711273, 1.551666, 1.45752, 1.344086, 1.188873, 1.041687, 0.9395142, 
    0.916748, 0.9961853, 1.116547, 1.201813, 1.287109, 1.4263, 1.620758, 
    1.801361, 1.909576, 1.910492, 1.779419, 1.413147, 0.9199219, 0.4666138, 
    0.1828308, 0.04107666, -0.04870605, -0.1533203, -0.2441406, -0.2774048, 
    -0.3344116, -0.3288879, -0.1285095, 0.1587219, 0.3883362, 0.5213623, 
    0.6390686, 0.7578735, 0.8744202, 1.030548, 1.263733, 1.527344, 1.722809, 
    1.82077, 1.858185, 1.909882, 1.990753, 2.036346, 2.081268, 2.114716, 
    2.061981, 1.829895, 1.683136, 1.646088, 1.715179, 1.920898, 2.335419, 
    2.787842, 2.912323, 2.54715, 2.598389, 2.926178, 3.681488, 4.625153, 
    4.931915, 4.802368, 4.846832, 4.975128, 5.208832, 5.422852, 5.561188,
  1.983551, 2.058044, 2.121063, 2.153717, 2.141418, 2.115295, 2.056763, 
    1.974731, 1.922211, 1.900635, 1.896606, 1.959625, 2.063477, 2.106903, 
    2.112244, 2.176605, 2.348114, 2.533539, 2.560944, 2.44696, 2.297607, 
    2.143433, 1.96701, 1.812683, 1.753754, 1.876556, 2.090729, 2.205933, 
    2.162231, 2.123688, 2.06955, 1.918488, 1.756287, 1.610931, 1.448395, 
    1.304077, 1.225128, 1.242584, 1.30011, 1.353119, 1.487518, 1.735687, 
    2.03775, 2.186401, 2.186432, 2.185333, 1.958923, 1.445374, 0.8740845, 
    0.491394, 0.3260498, 0.289917, 0.2416077, 0.1531372, 0.1487732, 
    0.2117615, 0.3076782, 0.4469299, 0.5940857, 0.698761, 0.7453613, 
    0.8178406, 0.9130859, 1.011139, 1.140289, 1.342377, 1.541565, 1.64212, 
    1.666412, 1.683228, 1.705231, 1.726624, 1.746033, 1.76297, 1.698242, 1.5, 
    1.5448, 2.10321, 2.099365, 1.695007, 1.614655, 1.675659, 2.011017, 
    1.891937, 1.66095, 1.661591, 1.831635, 2.014282, 2.10321, 2.102142, 
    2.078552, 2.063599, 2.058014, 2.043488, 1.996979, 1.949829,
  1.955902, 2.033966, 2.13504, 2.208649, 2.24707, 2.305206, 2.376495, 
    2.413818, 2.363037, 2.275513, 2.201172, 2.186127, 2.23938, 2.29303, 
    2.352661, 2.510284, 2.75177, 2.929626, 2.869141, 2.722534, 2.743103, 
    2.854156, 2.779938, 2.540802, 2.404938, 2.505615, 2.662292, 2.674347, 
    2.576508, 2.460876, 2.267181, 1.993622, 1.869049, 1.972809, 1.966736, 
    1.760742, 1.544739, 1.415436, 1.437347, 1.655212, 1.950012, 2.146149, 
    2.182831, 2.048767, 2.069916, 2.086121, 2.017914, 1.625763, 1.154175, 
    0.8513794, 0.7600708, 0.8250122, 0.9104309, 0.8769531, 0.8383484, 
    0.8791504, 0.9506531, 1.0495, 1.151367, 1.194458, 1.222839, 1.290863, 
    1.366974, 1.388672, 1.428253, 1.512299, 1.545654, 1.53952, 1.545227, 
    1.588348, 1.627808, 1.614136, 1.604126, 1.573303, 1.477539, 1.512238, 
    1.793945, 1.872711, 1.808044, 1.775208, 1.643616, 1.590973, 1.704803, 
    1.6026, 1.518219, 1.688599, 1.953705, 2.07782, 2.06073, 1.997192, 
    1.987885, 1.996033, 2.014374, 2.037323, 2.016663, 1.957153,
  2.285156, 2.358124, 2.416351, 2.415497, 2.412872, 2.489807, 2.673645, 
    2.809235, 2.837646, 2.914459, 3.040039, 3.085144, 3.063721, 3.012177, 
    2.952423, 2.904999, 2.977539, 3.198639, 3.30072, 3.50705, 3.87851, 
    3.972046, 3.572083, 3.049225, 2.791046, 2.725983, 2.615936, 2.378296, 
    2.152008, 1.890533, 1.616516, 1.530792, 1.63028, 1.747986, 1.741211, 
    1.624817, 1.486938, 1.421143, 1.476196, 1.79007, 2.391968, 2.572144, 
    2.312225, 2.195038, 2.433563, 2.575409, 2.15564, 1.891388, 1.613556, 
    1.391235, 1.450165, 1.575104, 1.664703, 1.687195, 1.663574, 1.592468, 
    1.463104, 1.460022, 1.578064, 1.667511, 1.686249, 1.68573, 1.667816, 
    1.641754, 1.642395, 1.636261, 1.598053, 1.602142, 1.60788, 1.596344, 
    1.591461, 1.587433, 1.590973, 1.546173, 1.489563, 1.514496, 1.681824, 
    1.715668, 1.807098, 1.797668, 1.721741, 1.563721, 1.486847, 1.381897, 
    1.353241, 1.621155, 1.990356, 2.203918, 2.256378, 2.228149, 2.181305, 
    2.183136, 2.183929, 2.156891, 2.159515, 2.21637,
  2.549194, 2.532776, 2.44574, 2.369812, 2.444305, 2.874359, 3.483887, 
    3.854065, 3.987488, 4.121063, 4.197083, 4.025024, 3.653107, 3.342407, 
    3.172699, 3.076324, 3.022339, 3.052246, 3.153015, 3.307343, 3.335388, 
    3.012482, 2.405579, 1.900635, 1.64566, 1.477966, 1.373077, 1.364197, 
    1.417236, 1.494415, 1.63858, 1.697113, 1.673645, 1.596924, 1.565521, 
    1.60611, 1.645844, 1.722565, 1.710327, 2.021973, 2.836029, 3.000153, 
    2.641357, 2.518463, 2.756287, 2.950897, 2.801086, 2.420105, 2.317932, 
    2.401489, 2.605713, 2.557526, 2.355835, 2.209412, 2.109192, 1.873993, 
    1.670746, 1.72287, 1.880615, 1.927399, 1.878632, 1.823944, 1.789886, 
    1.79425, 1.787689, 1.742096, 1.713104, 1.714539, 1.723083, 1.754456, 
    1.771912, 1.738708, 1.686707, 1.644043, 1.587769, 1.50528, 1.43512, 
    1.419525, 1.612152, 1.803162, 1.744629, 1.693085, 1.77121, 1.937256, 
    2.015839, 2.086304, 2.192535, 2.265137, 2.293396, 2.276276, 2.271332, 
    2.341675, 2.39209, 2.363586, 2.376526, 2.466309,
  2.332733, 2.264557, 2.210663, 2.287445, 2.556549, 3.072632, 3.232391, 
    3.373627, 3.470276, 3.366791, 2.875946, 2.437805, 2.082642, 1.863708, 
    1.802063, 1.888397, 1.991058, 2.042816, 2.041046, 1.886292, 1.608612, 
    1.265228, 1.018646, 0.9768066, 1.038513, 1.217194, 1.447235, 1.654999, 
    1.89566, 2.237732, 2.123474, 1.862915, 1.680176, 1.453156, 1.627106, 
    1.92804, 1.849365, 1.876617, 1.945221, 2.09082, 2.601868, 3.247955, 
    3.273804, 2.935791, 2.903992, 2.998016, 2.940918, 2.551056, 2.485748, 
    2.306488, 2.122955, 2.034729, 1.934021, 1.939758, 1.985321, 1.946594, 
    1.906921, 1.977509, 2.040283, 2.040466, 2.023468, 1.999969, 2.007843, 
    1.994843, 1.932953, 1.88382, 1.858368, 1.838776, 1.86142, 1.882324, 
    1.840851, 1.784515, 1.72287, 1.636902, 1.602325, 1.535004, 1.335693, 
    1.569397, 1.826172, 1.798126, 1.729126, 1.935516, 2.358551, 2.597168, 
    2.562531, 2.360901, 2.192871, 2.141174, 2.14801, 2.115265, 2.069641, 
    2.123016, 2.166046, 2.193146, 2.250427, 2.310974,
  2.166107, 2.066193, 1.999847, 2.116821, 2.259491, 2.371124, 2.475159, 
    2.314178, 2.347534, 2.211426, 1.404449, 1.296661, 1.327057, 1.326721, 
    1.301422, 1.37973, 1.500305, 1.529907, 1.438965, 1.277496, 1.27359, 
    1.43042, 1.606628, 1.810516, 1.986938, 2.115326, 2.166687, 2.257385, 
    2.456207, 2.279572, 1.712982, 1.632843, 1.645599, 1.612213, 1.778046, 
    1.886047, 1.75824, 1.8349, 2.097076, 2.333466, 2.646729, 3.140869, 
    3.684357, 3.473938, 3.147827, 3.098724, 2.774109, 2.343109, 1.964355, 
    1.503632, 1.380066, 1.534027, 1.718384, 1.878479, 2.007965, 2.052643, 
    2.079193, 2.124512, 2.112793, 2.113495, 2.111938, 2.071838, 2.043335, 
    2.017822, 1.982147, 1.972351, 1.90213, 1.819061, 1.801605, 1.736237, 
    1.643707, 1.609924, 1.56488, 1.481079, 1.414368, 1.227509, 0.9716492, 
    1.679047, 2.192657, 1.817078, 1.820099, 2.19223, 2.47644, 2.676544, 
    2.303925, 2.032257, 1.897034, 1.928406, 2.094574, 2.146118, 2.094482, 
    2.080627, 2.062469, 2.05011, 2.110626, 2.165802,
  1.846863, 1.775146, 1.737579, 1.780304, 1.826477, 2.765137, 3.267395, 
    3.316406, 3.193726, 2.133881, 1.939819, 2.017029, 1.958435, 1.85733, 
    1.867554, 1.982086, 2.048737, 2.034363, 2.025543, 2.083099, 2.239197, 
    2.339142, 2.347443, 2.34964, 2.342804, 2.339355, 2.347504, 2.334991, 
    2.214752, 1.840546, 1.695282, 1.843842, 1.861084, 1.759125, 2.052094, 
    2.186523, 2.097015, 2.260529, 2.564575, 3.081451, 3.302673, 2.777557, 
    2.661224, 2.697357, 2.647552, 2.482666, 2.128815, 1.804138, 1.630829, 
    1.625214, 1.822601, 1.992432, 2.055756, 2.080566, 2.129395, 2.148926, 
    2.110321, 2.10141, 2.10321, 2.103424, 2.097748, 2.091949, 2.082733, 
    2.050293, 2.007324, 1.899384, 1.710052, 1.54425, 1.429779, 1.340271, 
    1.281158, 1.264282, 1.172241, 1.151093, 1.118073, 0.9682007, 1.231354, 
    2.657471, 3.10437, 2.183014, 2.143127, 2.521576, 2.61145, 2.352753, 
    2.215912, 1.926544, 1.86731, 2.007965, 2.101471, 2.04657, 2.010071, 
    2.006744, 1.966309, 1.969238, 1.952179, 1.905914,
  1.513367, 1.495087, 1.683228, 1.919891, 2.348663, 3.41214, 3.950073, 
    3.786072, 3.536987, 2.283508, 2.012482, 2.146271, 2.201324, 2.147949, 
    2.242218, 2.415466, 2.50885, 2.46579, 2.446869, 2.452576, 2.436737, 
    2.394501, 2.370087, 2.294495, 2.252716, 2.183777, 2.107056, 2.036041, 
    1.974243, 1.95578, 1.964355, 2.214874, 2.375916, 2.486084, 2.504364, 
    2.493866, 2.566711, 2.581696, 2.433167, 3.274994, 3.543762, 2.27652, 
    1.947754, 1.972321, 2.058899, 2.099976, 2.121246, 2.130585, 2.15921, 
    2.209137, 2.213837, 2.153015, 2.11084, 2.089081, 2.088654, 2.087006, 
    2.036346, 2.030884, 2.031342, 2.043671, 2.011993, 1.98526, 1.933105, 
    1.871796, 1.740997, 1.496063, 1.305817, 1.101196, 1.031403, 1.000824, 
    1.00531, 1.073975, 1.066986, 1.009735, 0.8997192, 1.017761, 1.887482, 
    3.634766, 3.44812, 2.750061, 2.639557, 3.0466, 2.901337, 2.72226, 
    2.305756, 2.003693, 1.945557, 2.095612, 2.043854, 1.956757, 1.940338, 
    1.884735, 1.823608, 1.785126, 1.680084, 1.578552,
  1.699402, 1.889404, 2.191376, 2.604553, 3.918793, 4.04834, 4.396149, 
    4.645905, 4.152374, 3.683044, 2.109528, 2.188171, 3.431396, 2.309784, 
    2.309021, 2.325562, 2.309601, 2.320007, 2.305695, 2.313507, 2.264557, 
    2.195099, 2.155884, 2.09079, 2.065918, 2.08493, 2.078308, 2.158478, 
    2.173706, 2.268585, 2.255035, 2.49649, 2.783295, 2.977844, 2.987122, 
    2.76474, 2.688477, 2.453735, 2.874298, 3.430817, 3.158447, 2.279541, 
    2.341248, 2.488525, 2.491425, 2.40921, 2.344574, 2.289398, 2.239166, 
    2.182434, 2.125885, 2.098206, 2.10907, 2.097107, 2.082062, 2.082062, 
    2.117493, 2.119171, 2.081818, 2.083099, 2.02652, 1.952057, 1.842224, 
    1.684723, 1.466705, 1.218567, 1.065552, 0.9737549, 0.9725952, 1.010559, 
    1.070282, 1.07901, 1.055237, 0.9983215, 1.101593, 1.460114, 2.400574, 
    4.003998, 3.70285, 3.392517, 3.186035, 3.547302, 3.789093, 2.934998, 
    2.855042, 2.141266, 1.898834, 1.914093, 1.855835, 1.793213, 1.767365, 
    1.696594, 1.614532, 1.551056, 1.486298, 1.543732,
  2.126465, 2.370148, 2.523071, 2.713531, 4.133057, 3.882843, 4.216034, 
    4.505829, 3.895386, 3.505219, 2.203369, 2.295532, 3.420593, 2.963715, 
    2.263428, 2.306915, 2.244324, 2.236877, 2.272888, 2.278931, 2.295288, 
    2.285309, 2.273071, 2.262451, 2.253662, 2.334473, 2.389038, 2.38031, 
    2.366821, 2.486664, 2.53244, 2.457458, 3.249451, 3.424133, 3.560913, 
    3.456299, 3.380554, 3.396057, 3.902191, 3.477234, 2.360443, 2.561279, 
    2.715454, 2.706482, 2.638275, 2.518646, 2.370941, 2.29071, 2.223877, 
    2.143524, 2.12439, 2.163574, 2.176514, 2.194153, 2.222626, 2.251282, 
    2.261353, 2.226471, 2.182465, 2.157715, 2.054901, 1.95575, 1.817688, 
    1.640594, 1.458954, 1.304504, 1.248993, 1.199249, 1.233429, 1.229858, 
    1.231873, 1.237335, 1.257965, 1.403473, 1.497864, 1.72464, 2.452118, 
    4.426208, 3.277649, 3.539032, 3.714874, 4.042145, 4.4086, 3.271667, 
    3.147186, 3.135254, 1.988068, 1.974976, 1.931061, 1.872437, 1.80304, 
    1.772308, 1.730377, 1.764221, 1.853882, 1.950165,
  2.583038, 2.68689, 2.573547, 2.559784, 4.114197, 4.161438, 4.018982, 
    4.335846, 4.088379, 3.627502, 3.400238, 2.440735, 3.314606, 2.958771, 
    2.143127, 2.123138, 2.113037, 2.126617, 2.210663, 2.30191, 2.34729, 
    2.385834, 2.367401, 2.38559, 2.411926, 2.447235, 2.455231, 2.462128, 
    2.529541, 2.62674, 2.73114, 2.742493, 2.875031, 4.403625, 4.321198, 
    4.044037, 3.62558, 2.849579, 3.060516, 2.479462, 2.544586, 2.76239, 
    2.759796, 2.665924, 2.525574, 2.378601, 2.28595, 2.229736, 2.174957, 
    2.131195, 2.172272, 2.212463, 2.250366, 2.298096, 2.322632, 2.321442, 
    2.279785, 2.242432, 2.210571, 2.17041, 2.100037, 2.035065, 1.933258, 
    1.839233, 1.804138, 1.777313, 1.764099, 1.747345, 1.73996, 1.745911, 
    1.71402, 1.732635, 1.792938, 1.949707, 1.974792, 2.289154, 4.134735, 
    4.721161, 3.327911, 3.553955, 3.991516, 3.543365, 3.434692, 3.171783, 
    3.350616, 2.83136, 1.954651, 2.046722, 2.04715, 2.055298, 2.07785, 
    2.154022, 2.20816, 2.282135, 2.355896, 2.410004,
  2.68277, 2.610107, 2.501221, 2.442749, 3.773132, 3.787598, 3.609283, 
    3.804993, 3.79068, 3.441956, 3.455841, 2.504242, 2.365662, 2.147827, 
    2.046112, 2.11261, 2.124573, 2.181671, 2.215179, 2.343597, 2.316833, 
    2.33493, 2.320862, 2.329193, 2.404205, 2.429077, 2.446716, 2.502502, 
    2.565643, 2.612793, 2.705688, 2.732208, 2.791046, 2.952637, 2.942596, 
    3.524445, 3.388245, 2.603851, 2.762665, 2.423187, 2.525177, 2.667999, 
    2.625366, 2.50531, 2.371307, 2.239868, 2.199707, 2.171387, 2.172424, 
    2.177063, 2.146667, 2.133026, 2.17868, 2.242676, 2.249207, 2.255524, 
    2.224548, 2.227142, 2.218628, 2.180817, 2.180908, 2.176575, 2.147888, 
    2.11911, 2.12973, 2.132446, 2.121765, 2.130432, 2.154388, 2.195465, 
    2.200562, 2.255096, 2.3172, 2.313507, 2.430176, 3.900177, 3.940857, 
    3.676178, 3.445068, 4.036102, 4.020538, 3.60257, 3.493195, 3.18689, 
    3.09436, 2.69046, 2.035889, 2.14621, 2.197479, 2.235138, 2.297546, 
    2.367462, 2.439514, 2.527435, 2.580353, 2.669434,
  2.548187, 2.499237, 2.439178, 2.395935, 3.656799, 3.905914, 3.638062, 
    3.679138, 3.527008, 3.446381, 3.141571, 2.376984, 2.207916, 2.067017, 
    2.091034, 2.218109, 2.173401, 2.230713, 2.274323, 2.346436, 2.364746, 
    2.373779, 2.337585, 2.327454, 2.390411, 2.416809, 2.395508, 2.407745, 
    2.49411, 2.475494, 2.496521, 2.584229, 2.609344, 2.615326, 2.601593, 
    2.588379, 2.480499, 2.440399, 2.867035, 2.385437, 2.458954, 2.521667, 
    2.473663, 2.367035, 2.23526, 2.092407, 2.061035, 2.101654, 2.096436, 
    2.105316, 2.075806, 2.029388, 2.019897, 2.069092, 2.088043, 2.104462, 
    2.112518, 2.128754, 2.171448, 2.179901, 2.192474, 2.20047, 2.202393, 
    2.234222, 2.23819, 2.268158, 2.299774, 2.360962, 2.416962, 2.458954, 
    2.487396, 2.483246, 2.489288, 2.476196, 2.423889, 3.611115, 3.746521, 
    4.494476, 4.33493, 4.112457, 3.810577, 3.868073, 3.325989, 2.976654, 
    2.881348, 2.940979, 2.809479, 2.164185, 2.21756, 2.266327, 2.330322, 
    2.366974, 2.469086, 2.523651, 2.548798, 2.584015,
  2.451935, 2.50766, 2.572601, 2.708557, 3.914612, 3.609497, 3.530701, 
    3.336548, 3.401917, 2.811035, 2.968018, 2.334808, 2.210571, 2.212097, 
    2.222687, 2.316742, 2.419312, 2.461426, 2.48233, 2.449524, 2.419678, 
    2.404846, 2.396271, 2.451752, 2.460785, 2.496674, 2.400604, 2.40506, 
    2.566772, 2.434784, 2.43042, 2.450165, 2.484344, 2.455444, 2.499969, 
    2.359558, 2.213043, 2.403809, 2.672241, 2.760895, 2.358643, 2.333374, 
    2.286865, 2.247955, 2.101288, 2.046387, 2.048737, 2.069092, 2.054565, 
    2.042175, 2.040588, 2.030884, 2.032623, 2.054901, 2.072357, 2.093658, 
    2.098755, 2.106812, 2.134705, 2.159729, 2.191071, 2.22821, 2.237518, 
    2.264221, 2.276764, 2.308868, 2.34314, 2.368134, 2.421906, 2.436951, 
    2.424774, 2.338074, 2.321777, 2.356415, 2.27948, 3.685455, 4.504791, 
    3.717102, 3.754974, 3.857788, 3.993378, 3.343781, 3.160583, 2.956665, 
    2.837189, 3.116577, 2.783173, 2.185242, 2.25061, 2.322174, 2.366302, 
    2.354919, 2.441162, 2.464203, 2.484558, 2.468445,
  2.518188, 2.612396, 2.650879, 3.388702, 3.457245, 2.912811, 2.748138, 
    3.049591, 3.159149, 2.023682, 2.430756, 3.853424, 2.251587, 2.121124, 
    2.240479, 2.321259, 2.440033, 2.50235, 2.529968, 2.482483, 2.414978, 
    2.395905, 2.399353, 2.471161, 2.495117, 2.443542, 2.343842, 3.471771, 
    2.81073, 2.418091, 3.57196, 3.373383, 2.962402, 2.355743, 2.370483, 
    2.829254, 2.911041, 2.676788, 2.667877, 2.247284, 2.303345, 2.235596, 
    2.175537, 2.172089, 2.124054, 2.113068, 2.134277, 2.134338, 2.083435, 
    2.042419, 2.066681, 2.142609, 2.219482, 2.291046, 2.389374, 2.43808, 
    2.43689, 2.452454, 2.441071, 2.436829, 2.409393, 2.37204, 2.333221, 
    2.326843, 2.334869, 2.327637, 2.33551, 2.352386, 2.384583, 2.393127, 
    2.325806, 2.241974, 2.161102, 2.103882, 2.158966, 3.274353, 3.723755, 
    3.194702, 3.181488, 3.393768, 3.090271, 3.34613, 3.869385, 3.110046, 
    2.948853, 2.483704, 2.2117, 2.293549, 2.393372, 2.468018, 2.496063, 
    2.431427, 2.471771, 2.498413, 2.532593, 2.489441,
  2.348328, 2.514404, 2.564301, 2.898102, 2.760864, 2.686615, 2.856812, 
    2.901642, 2.905853, 2.586304, 2.121185, 3.226715, 3.711853, 2.131348, 
    2.182587, 2.366333, 2.469788, 2.503784, 2.413422, 2.33078, 2.260742, 
    2.269989, 2.269226, 2.434692, 2.589081, 2.420898, 2.371338, 3.035187, 
    2.351624, 2.326416, 3.347778, 2.744934, 2.319824, 2.169464, 2.116974, 
    2.097992, 2.029114, 2.073059, 2.164978, 2.203186, 2.138458, 2.130127, 
    2.152893, 2.164764, 2.138336, 2.139679, 2.146851, 2.113037, 2.106628, 
    2.105835, 2.112579, 2.155884, 2.219574, 2.29541, 2.378876, 2.430878, 
    2.435455, 2.438324, 2.44751, 2.466888, 2.439484, 2.403748, 2.388367, 
    2.377136, 2.381622, 2.384491, 2.368408, 2.352905, 2.333557, 2.295197, 
    2.177246, 2.095917, 1.944489, 1.880493, 1.904114, 2.539703, 2.888916, 
    2.834534, 2.915192, 3.048523, 2.931671, 3.750946, 4.008057, 2.444305, 
    2.375763, 2.358612, 2.243652, 2.221771, 2.257446, 2.405945, 2.463654, 
    2.3992, 2.41568, 2.431885, 2.383698, 2.32901,
  2.749054, 2.554382, 2.922638, 2.916779, 2.846588, 2.959351, 3.272614, 
    3.144226, 3.043732, 3.137665, 2.848724, 2.418396, 3.503265, 2.310394, 
    2.166962, 2.340881, 2.491516, 2.507599, 2.432037, 2.382813, 2.282074, 
    2.249908, 2.32901, 2.490021, 2.504028, 2.410431, 3.069244, 2.456726, 
    2.21756, 2.294464, 2.300934, 2.595673, 2.105743, 2.172028, 2.123718, 
    2.098511, 2.118988, 2.180145, 2.202759, 2.169464, 2.156677, 2.155487, 
    2.199982, 2.247314, 2.245331, 2.258881, 2.270691, 2.277374, 2.27887, 
    2.277496, 2.233612, 2.200775, 2.160461, 2.141418, 2.108429, 2.100433, 
    2.06958, 2.05954, 2.085114, 2.099243, 2.112488, 2.162476, 2.194183, 
    2.254211, 2.265015, 2.332642, 2.338318, 2.339081, 2.299561, 2.231659, 
    2.194489, 2.120728, 1.92804, 1.881805, 1.993652, 2.551788, 2.688293, 
    2.921265, 3.32843, 3.803833, 3.998383, 3.992889, 2.521362, 2.08786, 
    2.271912, 2.233826, 2.281494, 2.298645, 2.335449, 2.448669, 2.440247, 
    2.385315, 2.294495, 2.322754, 2.77002, 2.888397,
  2.97345, 2.845612, 2.851257, 2.93512, 2.940674, 2.952423, 2.883301, 
    3.034576, 2.999756, 3.071259, 3.271729, 3.302765, 3.626862, 3.856995, 
    2.270081, 2.220398, 2.463135, 2.568298, 2.54776, 2.472198, 2.39502, 
    1.905579, 2.487793, 2.406738, 2.420502, 2.445831, 2.476959, 2.279541, 
    2.38092, 2.409546, 2.400543, 2.180847, 2.176544, 2.483978, 2.118469, 
    2.104706, 2.141327, 2.121155, 2.159943, 2.151764, 2.152832, 2.151703, 
    2.182129, 2.218781, 2.271057, 2.277496, 2.273865, 2.297882, 2.296265, 
    2.288239, 2.282318, 2.274841, 2.255432, 2.234772, 2.199707, 2.171204, 
    2.12619, 2.094421, 2.082336, 2.089355, 2.115906, 2.13559, 2.115082, 
    2.139557, 2.175964, 2.288513, 2.318298, 2.368073, 2.387238, 2.359436, 
    2.321198, 2.375763, 2.274384, 2.023529, 2.46109, 2.426849, 2.848022, 
    3.445618, 3.9263, 3.542755, 2.330627, 2.365082, 2.226593, 2.151611, 
    2.158691, 2.162354, 2.271118, 2.326385, 2.385864, 2.393372, 2.443604, 
    2.343445, 2.284149, 2.766296, 2.817017, 2.982208,
  2.806152, 2.862427, 2.965668, 3.624542, 4.18335, 4.506317, 4.122437, 
    3.973206, 3.448364, 3.438171, 4.246857, 3.958069, 4.319397, 4.170929, 
    2.518555, 2.216888, 2.399139, 2.501251, 2.579437, 2.508453, 2.42926, 
    1.636444, 2.235535, 2.356781, 2.312103, 2.29837, 2.370361, 2.892731, 
    2.667603, 2.19339, 2.342712, 2.23645, 2.160919, 2.717651, 2.125641, 
    2.129822, 2.071167, 2.072906, 2.156372, 2.157776, 2.189484, 2.192413, 
    2.235992, 2.262451, 2.314941, 2.34259, 2.33728, 2.338318, 2.31488, 
    2.309875, 2.322327, 2.303741, 2.286713, 2.278168, 2.249329, 2.248535, 
    2.224426, 2.225372, 2.211853, 2.234619, 2.250092, 2.275696, 2.271179, 
    2.246857, 2.207916, 2.225281, 2.244629, 2.389191, 2.542694, 2.504547, 
    2.475586, 2.583984, 3.346405, 2.730835, 2.058563, 2.049255, 2.18161, 
    2.200867, 2.212006, 2.216156, 2.135437, 2.162933, 2.083435, 2.051788, 
    2.073669, 2.125824, 2.149261, 2.231476, 2.261627, 2.374847, 2.424896, 
    2.376862, 3.740875, 5.287628, 4.103577, 2.988434,
  3.933868, 4.209717, 4.512939, 4.524475, 4.223816, 3.795563, 3.766937, 
    3.775238, 3.679779, 3.465332, 3.37912, 3.834595, 4.048492, 4.111816, 
    3.088623, 2.349731, 2.420227, 2.472137, 2.594788, 2.508575, 2.312958, 
    1.677521, 2.055328, 2.420502, 2.377869, 2.313202, 2.77063, 2.775238, 
    2.044434, 2.059723, 2.181458, 2.375275, 2.210632, 2.008636, 2.094971, 
    2.118195, 2.051788, 2.076141, 2.133942, 2.171082, 2.190643, 2.125885, 
    2.159485, 2.1745, 2.217224, 2.241455, 2.267334, 2.303955, 2.307526, 
    2.294678, 2.318268, 2.334686, 2.310272, 2.258972, 2.210266, 2.15686, 
    2.10614, 2.079529, 2.062408, 2.11676, 2.171387, 2.258881, 2.313446, 
    2.264801, 2.084076, 1.863586, 1.82608, 2.239594, 2.654816, 2.722168, 
    2.997681, 3.761475, 3.607117, 1.988495, 2.114929, 2.079529, 2.078552, 
    2.090973, 2.029053, 2.059082, 2.077179, 2.027374, 2.017761, 2.069641, 
    2.085632, 2.056549, 2.017273, 2.045013, 2.048798, 2.206879, 2.308105, 
    2.360748, 4.507629, 6.516968, 5.653381, 4.522797,
  4.883423, 4.485107, 4.514587, 4.262909, 3.88974, 3.530609, 3.352295, 
    3.32608, 3.353882, 3.013885, 2.284058, 3.49704, 3.988586, 3.791168, 
    3.312866, 1.940216, 2.367798, 2.608124, 2.595032, 2.520538, 2.655365, 
    1.922363, 0.9897461, 1.605347, 2.463013, 2.508087, 2.450287, 2.233887, 
    2.22049, 2.176697, 2.093384, 2.260254, 2.25769, 2.196777, 2.195099, 
    2.151306, 2.100342, 2.149963, 2.156189, 2.155762, 2.111664, 2.069244, 
    2.055054, 2.024048, 2.011292, 2.02478, 2.04483, 2.060516, 2.058563, 
    2.064758, 2.073853, 2.062988, 2.045563, 2.054718, 2.027496, 1.940704, 
    1.901794, 1.843842, 1.751404, 1.770538, 1.790192, 1.866699, 1.947968, 
    1.997803, 1.805847, 1.444641, 1.34729, 2.078308, 3.538452, 2.998535, 
    3.243591, 4.443604, 4.073364, 2.109619, 2.220917, 2.140594, 2.068329, 
    2.018524, 1.980835, 1.949951, 1.952972, 2.01944, 2.033997, 1.998474, 
    1.943787, 1.941193, 1.892242, 1.821594, 1.772125, 1.822632, 1.976837, 
    2.47464, 4.496429, 5.913116, 6.015533, 5.671967,
  5.025085, 4.691498, 4.753387, 4.64917, 4.168152, 3.790955, 3.490112, 
    3.15741, 3.241425, 3.442596, 2.249664, 3.684662, 4.146667, 3.929016, 
    3.880585, 3.4935, 2.467529, 2.374573, 2.204407, 2.920197, 3.050354, 
    2.076141, 1.441193, 1.227509, 1.610016, 1.895996, 1.741821, 2.087128, 
    2.475983, 2.281494, 2.34549, 2.81839, 2.344238, 2.282928, 2.265137, 
    2.291046, 2.301331, 2.240448, 2.211151, 2.178101, 2.123077, 2.077362, 
    2.023041, 1.971527, 1.933563, 1.893921, 1.897644, 1.897247, 1.91806, 
    1.95636, 1.967804, 1.964355, 1.896454, 1.852325, 1.824921, 1.804871, 
    1.767609, 1.764679, 1.68512, 1.640289, 1.614288, 1.631195, 1.705231, 
    1.742889, 1.595978, 1.3591, 1.735077, 3.254974, 3.901123, 3.460449, 
    2.827515, 2.342926, 2.036102, 2.115326, 2.207123, 1.973938, 1.909607, 
    2.009277, 2.210236, 2.248291, 2.181671, 2.213898, 2.177246, 2.174713, 
    2.161865, 2.098999, 2.020081, 1.961121, 1.858551, 1.801392, 1.692474, 
    1.968323, 3.443634, 4.786102, 5.380737, 5.481567,
  5.011169, 4.861542, 5.058105, 4.855377, 4.465729, 3.964325, 3.785889, 
    3.402252, 2.948059, 3.492188, 3.848114, 4.003601, 3.907806, 3.714233, 
    3.870605, 4.253479, 3.865662, 3.499451, 3.678894, 4.017365, 3.592743, 
    2.099304, 2.137482, 2.887512, 2.32196, 2.409088, 2.537994, 2.647034, 
    3.150146, 3.055878, 2.967804, 3.108704, 3.049591, 2.410583, 2.430054, 
    2.461029, 2.438629, 2.396057, 2.401398, 2.298462, 2.192108, 2.124115, 
    2.109192, 2.10318, 2.084808, 2.06311, 1.996765, 1.932709, 1.915314, 
    1.896576, 1.953491, 2.020477, 2.009399, 1.941162, 1.876404, 1.842804, 
    1.77594, 1.760193, 1.723724, 1.716461, 1.698212, 1.67514, 1.701996, 
    1.61377, 1.413177, 1.592804, 3.10498, 3.838684, 2.830627, 2.026154, 
    2.16922, 2.410461, 2.541504, 2.756104, 2.970062, 1.986359, 1.961029, 
    2.126007, 2.205017, 2.187653, 2.166901, 2.253235, 2.329712, 2.364227, 
    2.343323, 2.27594, 2.238251, 2.165466, 2.038757, 1.951202, 1.751221, 
    1.658966, 2.032104, 3.539856, 4.769714, 5.276672,
  5.281769, 5.471924, 5.161407, 4.338196, 3.622894, 2.503082, 3.323181, 
    3.395691, 2.456207, 3.329681, 4.101379, 3.895355, 3.83728, 3.977814, 
    4.282471, 4.205872, 4.298187, 4.353699, 4.020355, 4.347809, 3.859619, 
    3.905304, 4.071228, 3.604492, 3.672668, 3.045044, 3.186584, 3.080627, 
    3.336426, 3.506592, 3.353027, 3.242584, 3.175507, 2.258942, 2.427063, 
    2.456543, 2.417816, 2.375641, 2.354889, 2.384918, 2.320129, 2.214752, 
    2.209625, 2.207916, 2.207275, 2.256073, 2.227509, 2.213257, 2.199066, 
    2.149719, 2.163666, 2.153748, 2.180176, 2.191559, 2.137329, 2.052185, 
    1.946899, 1.866577, 1.769135, 1.721832, 1.702332, 1.659454, 1.610901, 
    1.505951, 1.56723, 2.185883, 3.090363, 3.562317, 2.527008, 1.368103, 
    2.096375, 3.062683, 3.63974, 3.159851, 2.863708, 2.205383, 1.955231, 
    1.988037, 2.017151, 2.05777, 2.088226, 2.036163, 1.986115, 2.02301, 
    2.11972, 2.223785, 2.259552, 2.234406, 2.206238, 2.158234, 2.017181, 
    1.818634, 1.754791, 2.287994, 4.135193, 5.216644,
  5.61377, 5.484283, 5.118866, 2.86734, 2.305756, 2.189545, 2.43396, 
    2.682251, 2.690094, 2.787994, 3.776825, 3.941742, 4.35556, 5.373993, 
    4.707764, 4.267456, 4.303772, 4.476471, 4.793732, 4.862152, 5.483612, 
    4.190186, 3.721619, 3.236603, 2.910614, 3.013672, 3.307678, 3.839417, 
    3.237061, 3.038635, 2.855255, 2.756927, 2.770782, 2.262604, 2.673462, 
    2.691589, 2.942932, 3.056671, 2.593201, 2.49762, 2.435516, 2.36145, 
    2.330414, 2.34259, 2.332977, 2.334625, 2.303436, 2.345367, 2.394196, 
    2.395599, 2.386414, 2.31488, 2.266357, 2.254791, 2.229401, 2.171753, 
    2.102692, 2.013, 1.854126, 1.737091, 1.689819, 1.637604, 1.629547, 
    1.899902, 3.093323, 3.569885, 3.658813, 3.889679, 3.858551, 3.431274, 
    2.980377, 3.30899, 3.813202, 3.455627, 3.105591, 2.800598, 2.340729, 
    2.096039, 1.87262, 1.828949, 1.862457, 1.893311, 1.831848, 1.702759, 
    1.548126, 1.410645, 1.590393, 1.841766, 1.966766, 2.001587, 2.078918, 
    2.061676, 1.858612, 1.975342, 2.817688, 5.416504,
  4.607788, 2.346985, 2.383148, 2.494812, 2.331299, 2.454987, 4.538574, 
    4.38208, 3.607056, 3.464752, 3.997498, 4.337128, 4.921631, 4.894623, 
    2.942291, 4.300201, 4.53244, 3.925201, 4.176849, 6.123383, 5.232483, 
    4.380005, 4.064423, 3.89267, 3.377899, 3.207581, 3.639252, 3.958801, 
    3.089813, 2.651794, 2.667755, 2.39566, 2.472961, 2.645538, 2.631409, 
    2.455444, 2.39978, 2.643066, 2.596191, 2.663452, 2.78244, 2.828156, 
    2.749329, 2.704315, 2.659576, 2.569183, 2.463837, 2.470551, 2.505554, 
    2.498077, 2.497833, 2.463654, 2.343201, 2.27301, 2.22464, 2.149536, 
    2.074188, 2.036255, 1.890717, 1.744507, 1.725494, 1.646454, 1.781494, 
    3.051086, 3.657501, 3.969238, 3.34729, 3.849457, 4.525543, 4.375488, 
    3.985504, 3.722534, 3.749969, 3.759521, 3.590515, 3.453156, 3.173126, 
    2.676849, 2.237061, 1.921143, 1.86792, 1.954712, 1.875488, 1.518707, 
    1.055634, 0.4911194, 0.4860229, 1.002441, 1.338501, 1.565643, 1.80719, 
    1.901794, 1.957184, 2.425079, 4.614868, 5.400818,
  3.118927, 2.124115, 2.388367, 4.016418, 2.578033, 2.627625, 2.617096, 
    2.216187, 2.159454, 2.41626, 2.55426, 2.56955, 2.868256, 2.610657, 
    3.702179, 4.159576, 4.234467, 3.776642, 3.69809, 4.104462, 4.203094, 
    3.963257, 3.840515, 3.496643, 3.746246, 3.752075, 3.424316, 3.338959, 
    3.154022, 2.88089, 3.242432, 3.058563, 2.775177, 3.013702, 3.112793, 
    2.796661, 2.454468, 2.415527, 2.690155, 3.234924, 3.332153, 3.155151, 
    2.947144, 2.79245, 2.597321, 2.444275, 2.294617, 2.196442, 2.170715, 
    2.177307, 2.27002, 2.324036, 2.294952, 2.251648, 2.233368, 2.131866, 
    1.975037, 1.843353, 1.716705, 1.715271, 1.722626, 1.667023, 1.805023, 
    2.822815, 3.197693, 3.388519, 3.621826, 4.242279, 3.78595, 4.215332, 
    4.607056, 4.599487, 4.403625, 4.423584, 3.705231, 4.090271, 3.748199, 
    3.327911, 3.468628, 3.14267, 2.561676, 2.347565, 2.177887, 1.708252, 
    1.24234, 0.8791809, 0.7190247, 0.8189087, 0.8153992, 0.9944763, 1.371979, 
    1.570862, 1.688049, 2.073914, 3.637909, 3.866394,
  2.26474, 2.084534, 2.110565, 2.128235, 1.722107, 1.904663, 1.88031, 
    1.519592, 1.674377, 2.056793, 1.612274, 1.188782, 1.618073, 2.494446, 
    2.477844, 3.259949, 3.416443, 3.42926, 3.524628, 3.494446, 3.361176, 
    3.222687, 3.361389, 3.125427, 3.35321, 3.858978, 3.817688, 3.581024, 
    3.56485, 3.902832, 3.84671, 3.502258, 3.329987, 3.105042, 3.022766, 
    3.427704, 3.375488, 2.650696, 2.897186, 2.476746, 2.537018, 2.523254, 
    2.501312, 2.474548, 2.3862, 2.238678, 2.113556, 2.073761, 2.067505, 
    2.060394, 2.047119, 2.048492, 2.086334, 2.13092, 2.128754, 2.078979, 
    1.944122, 1.79834, 1.710297, 1.74762, 1.78302, 1.720795, 1.754913, 
    2.423157, 2.638458, 2.83136, 3.054138, 3.368134, 3.511566, 3.979218, 
    3.974854, 4.178162, 4.206879, 3.275726, 4.042023, 3.99762, 3.756439, 
    3.38739, 3.321533, 3.181702, 2.8461, 2.227936, 1.9151, 1.710876, 
    1.418365, 1.179901, 0.9553528, 0.7687988, 0.4782104, 0.4043274, 
    0.9069519, 1.399261, 1.622284, 1.671204, 1.86557, 2.325165,
  1.890839, 1.707336, 1.416321, 1.261688, 1.156403, 1.609528, 1.672485, 
    1.46344, 1.91684, 2.195129, 2.251831, 2.368469, 2.799255, 3.327271, 
    3.447998, 3.417755, 3.634613, 3.723206, 3.664551, 3.364227, 3.059387, 
    3.186432, 3.244934, 3.325592, 3.204559, 3.48468, 3.192657, 3.032104, 
    2.704681, 3.114349, 2.884583, 2.890076, 2.899323, 2.824066, 2.601074, 
    3.090729, 3.453094, 3.476868, 2.228119, 2.54126, 2.88855, 2.797333, 
    2.625854, 2.47937, 2.408905, 2.346039, 2.268951, 2.190613, 2.141968, 
    2.042755, 1.981049, 1.997894, 2.074097, 2.151489, 2.226501, 2.209503, 
    2.063293, 1.921448, 1.861359, 1.846893, 1.800659, 1.798737, 1.967346, 
    2.425354, 2.646027, 2.881805, 3.121643, 3.173584, 3.589264, 3.937012, 
    3.927399, 4.146729, 4.475708, 4.594055, 4.58136, 4.442535, 4.110779, 
    3.988617, 4.193756, 4.0625, 2.908264, 2.942444, 2.045593, 2.117004, 
    1.82135, 1.283203, 0.5863647, -0.07849121, -0.3744507, -0.2500305, 
    0.3361816, 0.9820557, 1.401917, 1.578491, 1.612274, 1.730499,
  1.369873, 1.493408, 1.09436, 1.261566, 1.663177, 1.9104, 2.017426, 
    2.161041, 2.662384, 3.046021, 3.500763, 3.662537, 3.69754, 3.825867, 
    3.801788, 4.07193, 4.134338, 3.941376, 3.685455, 3.087219, 2.672638, 
    2.639954, 2.626251, 2.970154, 2.751373, 2.702942, 2.462006, 2.353333, 
    2.4534, 2.366943, 1.880615, 1.763092, 1.786194, 2.18042, 2.349396, 
    2.342773, 2.561707, 2.855774, 2.06366, 2.414459, 2.977539, 3.004822, 
    3.036865, 2.245758, 2.363739, 2.350067, 2.340881, 2.280975, 2.20282, 
    2.175598, 2.215515, 2.322327, 2.411407, 2.444336, 2.471741, 2.422638, 
    2.257019, 2.102997, 2.002197, 1.905762, 1.739685, 1.801331, 2.010864, 
    2.72049, 2.760986, 2.893951, 2.979645, 2.962402, 3.222687, 3.643402, 
    4.139374, 4.657837, 4.959473, 5.169708, 5.064178, 1.517273, 3.842133, 
    3.741547, 3.758087, 3.646545, 3.204468, 1.8815, 1.657166, 1.527863, 
    1.266266, 1.246033, 0.7845154, -0.06463623, -0.6381226, -0.4885254, 
    0.1817322, 0.8364868, 1.217865, 1.34671, 1.466644, 1.562073,
  1.022278, 1.160828, 1.164429, 1.64502, 2.167816, 2.471405, 2.110962, 
    2.71759, 3.199524, 3.583038, 3.882477, 4.101898, 4.08609, 4.132782, 
    4.100891, 4.013428, 3.767151, 3.849548, 3.644287, 3.275024, 2.836365, 
    2.589417, 2.623993, 2.420959, 2.051727, 2.013519, 1.779663, 1.865814, 
    1.784271, 1.880157, 1.738342, 1.595703, 1.42514, 1.435944, 1.732483, 
    1.719574, 1.74823, 2.0784, 1.861267, 1.777466, 1.851044, 1.664154, 
    2.113281, 2.183075, 1.89505, 2.338409, 2.592834, 2.83313, 3.062042, 
    3.184387, 3.261383, 3.06015, 2.805969, 2.700378, 2.59552, 2.232422, 
    2.146149, 2.072052, 1.998505, 1.833466, 1.830505, 2.421753, 2.792358, 
    2.941071, 2.680023, 2.394836, 2.292023, 2.511688, 3.429504, 4.028229, 
    4.214111, 3.731171, 1.130585, 1.025604, 1.04422, 1.212708, 3.246887, 
    3.188293, 2.736206, 2.809448, 1.331665, 1.369751, 0.9736938, 0.3737488, 
    0.3059998, 0.8779297, 1.081238, 0.7467346, 0.3134766, 0.2705688, 
    0.5382385, 0.8630981, 1.08493, 1.126251, 1.162689, 1.222107,
  0.5961609, 0.7171021, 1.657074, 2.402527, 2.945709, 1.60379, 2.991455, 
    3.486755, 3.812073, 4.23877, 4.496521, 4.425995, 4.400391, 4.353912, 
    4.157959, 3.94577, 3.673065, 3.541595, 3.350189, 3.01709, 2.672882, 
    2.410248, 2.248749, 2.077301, 1.837555, 1.806488, 1.596039, 1.419525, 
    1.468231, 1.539124, 1.560608, 1.766693, 1.818237, 1.711487, 1.607361, 
    1.613861, 1.927094, 1.963867, 1.783905, 1.573425, 1.327148, 1.375732, 
    1.762909, 2.071869, 2.388397, 2.453064, 2.603851, 2.189911, 2.51062, 
    2.724213, 2.760345, 2.677917, 2.798767, 2.733276, 2.772552, 2.79538, 
    2.5784, 2.419006, 2.397736, 2.052856, 2.097321, 2.070831, 2.390625, 
    3.058929, 3.184601, 3.036224, 3.061432, 3.016937, 3.512756, 3.516235, 
    3.00351, 1.153259, 0.9402466, 0.8096313, 0.7902527, 0.8178406, 2.426941, 
    2.621216, 0.9567261, 0.8902283, 0.7988892, 0.8811646, 0.7322388, 
    0.4669189, 0.5968628, 0.2763062, 0.4190369, 0.7016296, 0.9248962, 
    1.07077, 1.093018, 0.7294006, 0.2246094, 0.1602173, 0.4539185, 0.5837708,
  0.09100342, 0.1806641, 0.4667969, 1.96756, 2.444672, 2.75351, 1.236603, 
    3.307739, 3.588013, 3.663025, 3.654877, 3.637329, 3.659088, 3.818817, 
    3.887756, 3.703247, 3.407166, 3.035919, 2.644196, 2.34256, 2.25293, 
    2.132172, 1.843018, 1.575195, 1.664856, 1.637909, 1.526703, 1.255524, 
    0.906189, 0.778595, 0.9562378, 1.179932, 1.364563, 1.375153, 1.604614, 
    1.707092, 1.90625, 2.261719, 2.326324, 2.227478, 1.849548, 1.857269, 
    2.041718, 2.46936, 2.855011, 3.004547, 2.574219, 2.327148, 2.814667, 
    1.874603, 1.599609, 1.36496, 1.935486, 2.26004, 2.338104, 2.215698, 
    1.85733, 1.662201, 1.66922, 1.654938, 1.55719, 1.744537, 1.921936, 
    2.227936, 2.574615, 2.785614, 2.945435, 2.933655, 2.854553, 2.585938, 
    2.606506, 2.90448, 3.324799, 3.463531, 1.165314, 0.8627319, 0.8353271, 
    2.335297, 2.134766, 1.742706, 0.6032715, 0.7949829, 1.174469, 1.718475, 
    1.713409, 1.49057, 0.9794922, 0.5093689, 0.5899658, 1.057556, 1.316803, 
    1.384003, 0.9298706, 0.1486206, -0.1774597, -0.1823425,
  0.3724365, 0.2974548, 0.3129578, 0.1373596, -0.1280518, 2.003387, 2.409821, 
    2.749847, 2.886841, 2.720184, 2.65097, 1.779236, 1.799591, 1.815887, 
    3.070892, 3.219666, 3.276154, 3.177002, 3.069733, 3.024689, 2.8125, 
    2.62384, 2.364258, 2.059723, 1.96698, 2.689728, 2.010864, 1.472137, 
    1.084229, 0.8184814, 0.7026062, 0.5804749, 0.6476746, 0.7832642, 
    0.9858093, 1.091156, 0.9134827, 0.9611206, 1.057892, 1.150055, 1.284851, 
    1.487701, 1.353638, 1.46991, 1.968292, 2.566193, 2.95874, 3.105408, 
    2.788483, 1.039215, 0.7597961, 0.4683838, 0.5831909, 1.377594, 1.596741, 
    1.703918, 1.704102, 1.345245, 1.095978, 1.236786, 1.055847, 1.290497, 
    1.380402, 1.717896, 1.992523, 2.303375, 2.592773, 2.540436, 2.439453, 
    1.127014, 2.392029, 2.791595, 3.17215, 1.421692, 2.514862, 0.9562073, 
    2.422058, 2.431641, 2.173309, 0.734314, 0.5464478, 0.6074219, 1.548187, 
    2.920837, 2.985931, 2.985565, 2.814209, 2.34198, 1.798248, 1.433655, 
    0.7412109, 0.8722839, 0.9934998, 0.913208, 0.8425293, 0.6217346,
  1.423431, 1.19223, 0.863739, 0.6738281, 0.4881592, 0.8925781, 1.722595, 
    2.314697, 2.366333, 2.2164, 1.89621, 1.709717, 1.525452, 1.231476, 
    1.025421, 2.331573, 1.374359, 1.385101, 1.264343, 2.453918, 2.283661, 
    2.239838, 1.937103, 1.857117, 1.853668, 1.703064, 1.591156, 1.349091, 
    1.002411, 0.6846313, 0.6835938, 0.5892029, 0.5583191, 0.5083923, 
    0.5140076, 0.3336487, 0.315094, 0.2956238, 0.993103, 1.175598, 0.6547546, 
    0.7251892, 0.7975464, 0.8820496, 0.9849243, 1.092072, 1.147919, 1.183777, 
    1.176147, 1.130066, 1.019592, 0.8741455, 0.7876892, 0.7677307, 0.7687683, 
    0.814209, 0.8517456, 0.7861633, 0.6587219, 0.5166626, 0.4241638, 
    0.3777466, 0.4953613, 1.947662, 2.400787, 2.694519, 2.904236, 2.790375, 
    2.674988, 1.042419, 2.484711, 2.552856, 1.291931, 3.046448, 3.029297, 
    3.046906, 2.581604, 1.428528, 1.222382, 0.9145813, 0.6497803, 1.890564, 
    2.891205, 3.415405, 3.69812, 3.713806, 3.373657, 2.967316, 2.775146, 
    2.330933, 1.771179, 0.7916565, 0.4963684, 0.6790771, 1.126373, 1.340881,
  1.130951, 1.388336, 1.512939, 1.81958, 2.003418, 1.557495, 1.515137, 
    1.342316, 1.261475, 1.211639, 1.205261, 1.22226, 1.24765, 1.307922, 
    1.380402, 1.472443, 1.508453, 1.504608, 1.442444, 1.32019, 1.102356, 
    0.9403992, 0.7989502, 0.6960449, 0.6428528, 2.236847, 2.325256, 1.557617, 
    1.482727, 1.434906, 1.284698, 0.5682373, 0.5838623, 0.6022949, 0.651825, 
    0.7223816, 0.7712097, 0.8362122, 0.9029846, 0.9794922, 1.038483, 
    1.155609, 1.256714, 1.280151, 1.287964, 1.298431, 1.307861, 1.310486, 
    1.361664, 1.397858, 1.42865, 1.472839, 1.580292, 1.655975, 1.668427, 
    1.654877, 1.610931, 1.539429, 1.448059, 1.351624, 1.277679, 1.204437, 
    1.200867, 1.20462, 1.195465, 3.223663, 3.31192, 3.311279, 3.231201, 
    3.190826, 2.969757, 2.54187, 2.66571, 2.988495, 2.767883, 1.516022, 
    1.592621, 1.509766, 2.659882, 2.833679, 3.092651, 3.292389, 3.516479, 
    3.63443, 3.681519, 3.671814, 3.503601, 3.321014, 3.055511, 2.757599, 
    2.316132, 2.12149, 0.9318237, 0.89505, 0.6530457, 0.683136,
  1.188019, 1.17395, 1.089081, 0.9889221, 1.800781, 1.8172, 1.862579, 
    1.636078, 1.675964, 1.672394, 1.669464, 1.670898, 1.672028, 1.64856, 
    1.64505, 1.611267, 1.560211, 1.518158, 1.495117, 1.442657, 1.354614, 
    1.261871, 1.147125, 1.029724, 0.8371277, 1.515747, 1.508148, 1.158844, 
    1.175262, 1.172974, 1.127289, 1.07312, 1.031006, 1.019989, 1.025208, 
    1.011414, 0.9889526, 1.002106, 1.027985, 1.077332, 1.124817, 1.182098, 
    1.206635, 1.24765, 1.324921, 1.422394, 1.458405, 1.479034, 1.498291, 
    1.515167, 1.520905, 1.500061, 1.506134, 1.4953, 1.496399, 1.511139, 
    1.517517, 1.516327, 1.480286, 1.446472, 1.409119, 1.352814, 1.319977, 
    1.335815, 1.369843, 1.467377, 1.545746, 1.61731, 1.658783, 1.653076, 
    1.587433, 2.907501, 3.379242, 2.761078, 2.906372, 3.013275, 3.038605, 
    3.072845, 3.009827, 3.010834, 2.998779, 3.024475, 3.032166, 3.076447, 
    3.195953, 3.160004, 3.055542, 2.95755, 2.828186, 2.666412, 2.537109, 
    2.343811, 1.452393, 1.35675, 1.340637, 1.262817,
  1.707733, 1.67453, 1.67218, 1.653137, 1.651611, 1.659424, 1.687897, 
    1.728851, 1.780731, 1.829376, 1.864624, 1.882935, 1.910034, 1.917053, 
    1.921722, 1.922638, 1.908478, 1.879028, 1.840607, 1.797607, 1.746094, 
    1.721802, 1.666138, 1.625183, 1.585358, 1.54303, 1.512756, 1.469452, 
    1.424622, 1.397156, 1.368164, 1.336212, 1.307678, 1.287964, 1.288605, 
    1.288635, 1.293182, 1.319855, 1.380402, 1.440582, 1.473877, 1.494598, 
    1.539276, 1.56189, 1.600464, 1.609772, 1.62793, 1.626953, 1.616669, 
    1.590027, 1.563599, 1.540558, 1.506592, 1.49765, 1.492706, 1.487305, 
    1.481842, 1.477325, 1.490234, 1.509705, 1.522705, 1.529663, 1.568604, 
    1.585144, 1.58429, 1.602661, 1.660156, 1.712494, 1.797607, 1.839447, 
    1.868408, 1.886017, 1.937866, 1.991089, 2.049713, 2.049927, 2.106903, 
    2.150726, 2.193176, 2.24646, 2.266937, 2.311584, 2.347015, 2.390106, 
    2.410095, 2.380524, 2.35144, 2.306366, 2.213867, 2.136139, 2.057434, 
    1.976349, 1.919006, 1.850983, 1.777008, 1.725067,
  1.940369, 1.926239, 1.92804, 1.92688, 1.921021, 1.913605, 1.904907, 
    1.898773, 1.908386, 1.932343, 1.952484, 1.956116, 1.958649, 1.969208, 
    1.976837, 1.969788, 1.970703, 1.964111, 1.963562, 1.962433, 1.967438, 
    1.954559, 1.949738, 1.94043, 1.931061, 1.904358, 1.886475, 1.880341, 
    1.871613, 1.851959, 1.838074, 1.823608, 1.815765, 1.829224, 1.826996, 
    1.824036, 1.829376, 1.82547, 1.837036, 1.83728, 1.838165, 1.855408, 
    1.864044, 1.870331, 1.874481, 1.890564, 1.887634, 1.880585, 1.895172, 
    1.898499, 1.90451, 1.917053, 1.928253, 1.940552, 1.956573, 1.954956, 
    1.948761, 1.941101, 1.928131, 1.920898, 1.924133, 1.929443, 1.952454, 
    1.963531, 1.992371, 2.016388, 2.009521, 1.995972, 1.994202, 1.983215, 
    1.983643, 1.994263, 1.990936, 1.995911, 1.996002, 1.998749, 2.006531, 
    2.010651, 2.018616, 2.034637, 2.044617, 2.064453, 2.064392, 2.065308, 
    2.05899, 2.052032, 2.035675, 2.030579, 2.018951, 2.011566, 2.01297, 
    1.998199, 1.973175, 1.958588, 1.953278, 1.944519,
  2.022385, 2.039581, 2.054306, 2.06485, 2.072662, 2.073303, 2.072342, 
    2.065826, 2.059113, 2.048248, 2.030792, 2.012985, 1.99437, 1.972824, 
    1.947952, 1.922562, 1.895081, 1.865326, 1.833099, 1.799973, 1.768204, 
    1.738846, 1.716568, 1.703278, 1.701065, 1.705887, 1.716187, 1.731018, 
    1.748413, 1.771255, 1.794952, 1.818939, 1.844528, 1.869202, 1.899155, 
    1.929886, 1.960678, 1.988602, 2.015427, 2.043762, 2.07103, 2.099548, 
    2.128769, 2.156967, 2.184509, 2.206635, 2.222916, 2.264389, 2.286453, 
    2.299606, 2.305984, 2.314072, 2.349609, 2.378067, 2.36998, 2.391144, 
    2.389328, 2.449219, 2.471939, 2.44133, 2.420761, 2.527527, 2.448502, 
    2.485672, 2.479218, 2.470322, 2.458069, 2.427155, 2.387238, 2.323044, 
    2.278839, 2.216537, 2.124084, 2.239258, 2.1362, 2.086258, 2.072784, 
    2.137894, 1.961517, 1.966537, 1.957413, 1.944397, 1.926956, 1.923248, 
    1.918625, 1.912369, 1.906189, 1.903061, 1.903061, 1.906387, 1.913986, 
    1.927994, 1.949615, 1.967697, 1.985947, 2.005478,
  2.522781, 2.546753, 2.557877, 2.561325, 2.555542, 2.547028, 2.539825, 
    2.532776, 2.526077, 2.517548, 2.505707, 2.493332, 2.484604, 2.464798, 
    2.433548, 2.400223, 2.374969, 2.352249, 2.257523, 2.142288, 1.983688, 
    1.828934, 1.677826, 1.553024, 1.47049, 1.452438, 1.484467, 1.544495, 
    1.617676, 1.690201, 1.751923, 1.789978, 1.812897, 1.838669, 1.882889, 
    1.955276, 2.058456, 2.186401, 2.347397, 2.526749, 2.711136, 2.947403, 
    3.199478, 3.454483, 3.696365, 3.973831, 4.152542, 4.345825, 4.533081, 
    4.714706, 4.788086, 4.820847, 4.849426, 4.83255, 4.829819, 4.715363, 
    4.609192, 4.507935, 4.375061, 4.283142, 4.243423, 4.211197, 4.218826, 
    4.238419, 4.251434, 4.239441, 4.174408, 4.053772, 3.903244, 3.724869, 
    3.477936, 3.287369, 3.15332, 3.088013, 3.042252, 2.899017, 2.794144, 
    2.700714, 2.677353, 2.537048, 2.442581, 2.382736, 2.336197, 2.347076, 
    2.273956, 2.295822, 2.202148, 2.177933, 2.178253, 2.197403, 2.237701, 
    2.29837, 2.364395, 2.43132, 2.483459, 2.510666,
  2.441528, 2.441284, 2.570572, 2.771057, 2.989746, 3.183426, 3.210983, 
    3.168594, 3.110901, 3.074646, 2.938904, 2.765778, 2.578934, 2.385971, 
    2.258041, 2.214676, 2.22699, 2.220215, 2.178101, 2.159805, 2.17041, 
    2.203934, 2.311493, 2.468964, 2.509979, 2.340698, 2.111801, 1.983246, 
    1.912781, 1.855499, 1.828674, 1.838898, 1.903107, 1.988144, 2.041595, 
    2.065887, 2.102539, 2.171875, 2.309891, 2.500259, 2.73764, 3.077866, 
    3.609055, 4.419464, 5.409775, 6.116272, 6.376236, 6.398758, 6.407867, 
    6.393295, 6.386978, 6.473114, 6.635864, 6.822266, 6.938019, 6.973373, 
    6.769989, 6.343948, 5.866013, 5.47142, 5.115356, 4.90358, 4.755539, 
    4.582748, 4.364639, 4.201569, 4.019653, 3.933334, 3.881119, 3.881577, 
    3.878906, 3.847931, 3.735535, 3.586075, 3.430725, 3.30899, 3.234756, 
    3.167572, 3.093094, 2.947067, 2.871674, 2.886337, 2.799026, 2.77388, 
    2.755005, 2.749023, 2.712173, 2.639786, 2.622971, 2.628906, 2.607025, 
    2.580719, 2.579361, 2.556183, 2.512894, 2.473633,
  2.366486, 2.459045, 2.690094, 2.907578, 3.115601, 3.301727, 3.336365, 
    3.17009, 2.987915, 2.795013, 2.60701, 2.49411, 2.467285, 2.428253, 
    2.347458, 2.300583, 2.174469, 2.071289, 2.042313, 1.853836, 1.658737, 
    1.497513, 1.373764, 1.337692, 1.76741, 2.298981, 2.206284, 2.008881, 
    2.034409, 2.242096, 2.540604, 2.804001, 2.918976, 2.832718, 2.600494, 
    2.403351, 2.315155, 2.240295, 2.230927, 2.218811, 2.283142, 2.399872, 
    2.653, 3.191071, 4.245117, 5.723373, 4.236984, 4.471802, 4.542252, 
    4.729492, 4.925919, 5.121231, 5.174545, 5.313354, 5.376694, 5.286194, 
    4.672455, 5.44075, 5.143372, 4.829941, 4.68132, 4.366928, 4.160095, 
    4.035355, 3.960342, 3.87767, 3.762894, 3.714584, 3.656448, 3.635086, 
    3.59668, 3.544464, 3.519531, 3.480408, 3.43222, 3.476044, 3.536316, 
    3.542969, 3.501755, 3.42897, 3.460739, 3.499283, 3.419067, 3.433853, 
    3.421478, 3.438354, 3.553253, 3.532425, 3.74588, 2.827667, 2.720963, 
    2.692505, 2.596802, 2.537689, 2.447647, 2.411652,
  3.011002, 2.980408, 2.955399, 2.959305, 3.044205, 3.127594, 3.149872, 
    3.104431, 3.110352, 2.947525, 2.829102, 2.804565, 2.894531, 2.996811, 
    3.007813, 2.798828, 2.569275, 2.376877, 2.269073, 2.054886, 1.597076, 
    1.525909, 1.630341, 1.611923, 1.423187, 1.307159, 1.288544, 1.353836, 
    1.460556, 1.63913, 1.882233, 2.078583, 2.260666, 2.430145, 2.638412, 
    2.869522, 3.157806, 3.1306, 2.704559, 2.269913, 2.143555, 2.246017, 
    2.504166, 2.969147, 3.710999, 4.829178, 4.548309, 4.86322, 5.001694, 
    5.324738, 5.564453, 5.639648, 5.455399, 5.208984, 4.830841, 4.496277, 
    4.00441, 3.747177, 3.755905, 3.824661, 3.889374, 3.965805, 3.81398, 
    3.717621, 3.613724, 3.510208, 3.400635, 3.455719, 3.507355, 3.478134, 
    3.50943, 2.822311, 3.142822, 3.314514, 3.482025, 3.472839, 4.053116, 
    4.056641, 3.984497, 3.842972, 3.409286, 3.414627, 3.396606, 3.464828, 
    3.556885, 3.624069, 3.707932, 3.791916, 3.917435, 4.145676, 3.957092, 
    3.558594, 3.236649, 3.171158, 3.101685, 3.057358,
  5.800568, 4.909485, 4.803787, 4.376892, 4.106583, 3.91452, 3.855804, 
    3.824539, 3.785873, 3.764511, 3.729691, 3.398621, 3.122986, 2.964905, 
    2.879364, 2.819336, 2.573303, 2.390366, 2.317978, 2.486328, 2.496353, 
    2.2845, 2.064453, 1.878204, 1.689529, 1.604553, 1.558136, 1.484253, 
    1.376892, 1.251694, 1.246475, 1.19902, 1.166931, 1.184509, 1.209045, 
    1.295822, 1.368225, 1.434235, 1.525772, 1.732025, 2.026627, 2.44043, 
    2.920044, 3.525589, 3.844864, 4.284622, 4.422211, 4.266907, 4.214767, 
    4.297562, 4.442505, 4.5354, 4.476578, 4.281006, 4.022079, 3.75705, 
    3.604187, 3.582108, 3.743378, 3.87529, 3.932373, 3.990967, 4.047867, 
    4.02507, 4.022278, 4.041153, 3.952744, 3.955551, 3.980103, 4.011078, 
    3.953964, 3.937943, 4.150833, 4.262421, 4.429474, 4.549591, 4.693863, 
    4.740158, 4.933182, 4.73468, 4.36821, 4.391327, 4.370956, 4.340118, 
    4.433319, 4.521729, 4.544128, 4.496399, 4.422241, 4.230377, 4.107788, 
    4.164627, 4.278961, 4.616852, 5.02153, 5.426422,
  6.49614, 6.635925, 6.555588, 6.35051, 6.141388, 6.092758, 6.036179, 
    5.88501, 5.710083, 5.545044, 5.336182, 5.220032, 5.159164, 5.134613, 
    4.821594, 4.225647, 3.939636, 3.89621, 4.00975, 4.107086, 4.049469, 
    3.870819, 3.548477, 3.209549, 2.901871, 2.724777, 2.695099, 2.683441, 
    2.447311, 2.101746, 1.849136, 1.629883, 1.196365, 1.264374, 1.007599, 
    0.9342346, 1.029434, 1.284164, 1.52916, 1.848953, 2.180527, 2.384872, 
    2.517365, 2.548279, 2.627335, 2.621689, 2.623016, 2.45108, 2.031708, 
    1.450745, 1.075592, 1.193298, 1.246948, 1.2948, 1.455078, 1.490967, 
    1.975922, 2.11377, 2.565887, 3.096039, 3.335388, 3.725281, 4.304443, 
    5.067261, 5.556915, 6.163452, 6.817322, 6.800232, 7.042999, 7.057251, 
    7.134521, 7.661285, 8.090515, 8.444336, 8.257172, 7.706512, 6.727478, 
    6.089142, 5.686981, 5.729767, 5.548645, 5.303986, 5.168961, 5.133484, 
    5.216553, 5.307846, 5.487778, 5.616364, 5.547028, 5.376923, 5.233643, 
    5.122314, 5.063522, 5.212738, 5.549149, 6.064621,
  7.540817, 8.153091, 8.519882, 8.725861, 9.02182, 9.399292, 9.629517, 
    9.535126, 9.333832, 9.138885, 9.300598, 9.638947, 9.829834, 9.967941, 
    9.576447, 9.208084, 8.375259, 7.706589, 7.173523, 6.564148, 5.902344, 
    5.372238, 5.126312, 4.808289, 4.81897, 4.805023, 4.858475, 4.57991, 
    4.481766, 3.839722, 2.788879, 2.73349, 2.261597, 1.832703, 1.416626, 
    1.68811, 2.79303, 2.923523, 2.770264, 2.658691, 2.741028, 3.058502, 
    3.075287, 2.845398, 2.41571, 1.862457, 1.105469, 0.256012, -0.3468628, 
    -0.5829163, -0.7534485, -0.955658, -1.131622, -1.20224, -0.914093, 
    -0.5006409, 0.09063721, 0.4779663, 1.271179, 2.011292, 2.282166, 
    2.459656, 2.430756, 2.215332, 2.185883, 2.227234, 2.309326, 2.447601, 
    2.509857, 2.534546, 2.647949, 2.883911, 3.173248, 3.379303, 3.542145, 
    3.546692, 3.436737, 3.233551, 3.462006, 4.38974, 5.492401, 5.59552, 
    5.749023, 6.002167, 6.137787, 6.257507, 6.413177, 6.464981, 6.470673, 
    6.436737, 6.411148, 6.210968, 6.079117, 6.097427, 6.230606, 6.803467,
  6.51297, 6.321289, 6.220123, 6.148438, 6.216492, 6.209595, 6.041809, 
    5.362457, 4.61792, 4.429901, 4.334839, 4.380157, 4.539734, 4.692261, 
    5.031281, 5.342987, 5.69162, 6.079773, 6.653076, 6.854004, 6.315002, 
    6.332245, 6.264862, 5.784698, 5.170532, 4.782959, 4.324371, 4.059845, 
    3.579315, 3.30658, 2.720215, 1.975952, 1.601959, 1.365387, 1.24054, 
    1.226013, 1.245422, 1.28598, 1.342102, 1.476929, 1.670715, 1.880066, 
    2.147339, 2.334229, 2.250519, 2.114075, 1.744873, 1.100189, 0.5615845, 
    0.3167725, 0.2240295, 0.0930481, -0.07687378, -0.22229, -0.3282471, 
    -0.3548584, -0.2205811, 0.0390625, 0.3606567, 0.6849365, 0.9430237, 
    1.102478, 1.228607, 1.32663, 1.469269, 1.676025, 1.922211, 2.056427, 
    2.074554, 2.046875, 2.03302, 2.096619, 2.1651, 2.150665, 2.122345, 
    1.980988, 1.719482, 1.625336, 1.659515, 1.743622, 1.900055, 2.25943, 
    3.2146, 4.421173, 4.954834, 5.401184, 5.990631, 6.55719, 6.670013, 
    7.087189, 7.394928, 7.206451, 6.843201, 6.248322, 5.989471, 6.261414,
  2.887451, 2.830414, 2.826508, 2.780487, 2.694489, 2.660675, 2.599548, 
    2.402679, 2.263214, 2.180023, 2.135925, 2.119019, 2.12326, 2.179291, 
    2.299103, 2.454529, 2.716736, 3.072266, 3.269684, 3.237305, 3.138275, 
    2.778931, 2.396301, 2.26413, 2.208405, 2.307159, 2.481506, 2.541809, 
    2.485931, 2.406036, 2.273438, 2.018402, 1.825287, 1.814789, 1.905792, 
    1.88562, 1.724426, 1.540833, 1.442383, 1.4888, 1.740356, 2.104828, 
    2.453979, 2.443726, 2.251099, 2.104889, 2.036987, 1.765106, 1.275452, 
    0.8185425, 0.553772, 0.417572, 0.2877502, 0.2209778, 0.2329407, 0.281311, 
    0.4210205, 0.563324, 0.7066956, 0.8311157, 0.9489136, 1.067322, 1.145569, 
    1.208344, 1.309753, 1.447479, 1.592316, 1.679443, 1.723694, 1.774689, 
    1.822845, 1.871826, 1.881653, 1.78299, 1.555267, 1.336792, 1.41922, 
    2.031311, 2.034821, 1.510162, 1.493866, 1.675323, 2.343018, 2.441345, 
    2.234436, 2.226837, 2.425201, 2.673981, 2.792572, 2.800446, 2.61499, 
    2.518829, 2.49292, 2.601837, 2.841949, 2.945587,
  2.134399, 2.257172, 2.40033, 2.450592, 2.42038, 2.436676, 2.505585, 
    2.548767, 2.523682, 2.487549, 2.463104, 2.436157, 2.444519, 2.470184, 
    2.498871, 2.614655, 2.883606, 3.168427, 3.104889, 2.962494, 2.964172, 
    3.114868, 3.0466, 2.808075, 2.659241, 2.733856, 2.889771, 2.922516, 
    2.815704, 2.629791, 2.369415, 2.044403, 1.847382, 1.897339, 2.124176, 
    2.171875, 1.90448, 1.622681, 1.478729, 1.610413, 2.026184, 2.365295, 
    2.355988, 2.208069, 2.205597, 2.171814, 2.134247, 1.957611, 1.416138, 
    0.97995, 0.8715515, 0.9330139, 0.9836426, 0.9898987, 0.957489, 0.9609985, 
    1.01532, 1.101135, 1.199341, 1.232147, 1.26828, 1.363983, 1.393738, 
    1.360168, 1.357422, 1.368805, 1.359711, 1.371368, 1.384888, 1.398254, 
    1.430267, 1.469269, 1.476501, 1.394135, 1.240631, 1.379883, 1.997009, 
    2.147095, 1.935699, 1.835297, 1.661316, 1.545258, 1.874756, 1.782166, 
    1.628235, 1.742828, 1.98468, 2.146637, 2.141052, 2.085999, 2.012695, 
    1.957825, 1.971039, 2.031769, 2.060822, 2.074097,
  2.241943, 2.387512, 2.507294, 2.574402, 2.611633, 2.702942, 2.872223, 
    3.040436, 3.128906, 3.259338, 3.425201, 3.467041, 3.399292, 3.291016, 
    3.133667, 2.975983, 3.028503, 3.35376, 3.542145, 3.748108, 4.13974, 
    4.344025, 3.979431, 3.391663, 3.068024, 2.959259, 2.885559, 2.759033, 
    2.580139, 2.305786, 1.990753, 1.808716, 1.757965, 1.767334, 1.777466, 
    1.664734, 1.475891, 1.337433, 1.272736, 1.454895, 2.154053, 2.53775, 
    2.326477, 2.200378, 2.507751, 2.832245, 2.295441, 2.073395, 1.808075, 
    1.506561, 1.580811, 1.78537, 1.851807, 1.799988, 1.729675, 1.657318, 
    1.560486, 1.502991, 1.558655, 1.590454, 1.58078, 1.557434, 1.517181, 
    1.504059, 1.52533, 1.489075, 1.430481, 1.432281, 1.444794, 1.419922, 
    1.39682, 1.367889, 1.3703, 1.376648, 1.34256, 1.372986, 1.747467, 
    1.841888, 1.871674, 1.808197, 1.689056, 1.557495, 1.532928, 1.420258, 
    1.422272, 1.633911, 1.941528, 2.151825, 2.18573, 2.067444, 1.938934, 
    1.923004, 1.956116, 1.968109, 1.995697, 2.100128,
  2.398682, 2.478241, 2.491882, 2.487579, 2.554047, 2.931854, 3.605591, 
    4.071686, 4.262054, 4.432281, 4.562714, 4.414795, 3.938324, 3.474152, 
    3.183655, 3.040192, 3.0112, 3.127289, 3.322845, 3.51651, 3.584656, 
    3.30542, 2.733398, 2.240356, 2.010925, 1.871094, 1.719055, 1.580078, 
    1.501404, 1.454407, 1.525574, 1.594208, 1.562103, 1.452148, 1.375519, 
    1.399017, 1.434113, 1.506714, 1.55014, 1.763916, 2.524353, 2.855225, 
    2.575012, 2.447205, 2.747528, 3.041901, 3.053192, 2.440369, 2.367188, 
    2.426636, 2.655212, 2.664642, 2.45697, 2.266022, 2.158386, 1.981781, 
    1.737885, 1.658081, 1.717194, 1.737885, 1.727997, 1.700134, 1.65863, 
    1.647797, 1.646301, 1.597137, 1.541473, 1.550903, 1.527283, 1.480743, 
    1.466217, 1.484253, 1.507111, 1.516083, 1.44458, 1.262299, 1.214996, 
    1.466492, 1.64389, 1.738739, 1.684784, 1.62146, 1.696228, 1.87381, 
    1.98938, 2.087585, 2.19101, 2.248718, 2.249664, 2.160736, 2.058716, 
    2.0867, 2.134827, 2.130615, 2.166931, 2.268219,
  2.247406, 2.20401, 2.141998, 2.200409, 2.5513, 3.190613, 3.409058, 
    3.467712, 3.522644, 3.398895, 2.977295, 2.569611, 2.138611, 1.828064, 
    1.705261, 1.77063, 1.912048, 2.02713, 2.03476, 1.892853, 1.652222, 
    1.343018, 1.076508, 0.9563293, 0.9033203, 0.944397, 1.055145, 1.223114, 
    1.555725, 2.134857, 2.1698, 1.833008, 1.532684, 1.152924, 1.157349, 
    1.6427, 1.682465, 1.69455, 1.790741, 1.930542, 2.330841, 2.973297, 
    3.172546, 2.90686, 2.902222, 3.072418, 3.01413, 2.997253, 2.595306, 
    2.401825, 2.214142, 2.136963, 2.00592, 1.896423, 1.912933, 1.876556, 
    1.807617, 1.787506, 1.819519, 1.818481, 1.823822, 1.831909, 1.83197, 
    1.85965, 1.853729, 1.832031, 1.821289, 1.800262, 1.778442, 1.745514, 
    1.71991, 1.674164, 1.623444, 1.543945, 1.450317, 1.298645, 1.200653, 
    1.347076, 1.596802, 1.608612, 1.673615, 1.937958, 2.344543, 2.629944, 
    2.85318, 2.691864, 2.463348, 2.307678, 2.23407, 2.201569, 2.200104, 
    2.220306, 2.172852, 2.11264, 2.116119, 2.182373,
  2.090698, 2.015564, 1.94989, 2.082184, 2.314453, 2.410095, 2.474945, 
    2.311401, 2.457825, 2.2789, 1.494293, 1.336548, 1.314697, 1.251495, 
    1.180847, 1.217773, 1.298126, 1.291687, 1.160797, 0.9263611, 0.8235168, 
    0.8709717, 0.9971313, 1.225525, 1.475311, 1.700317, 1.911499, 2.170959, 
    2.53772, 2.449432, 1.796753, 1.65271, 1.629425, 1.552612, 1.640564, 
    1.781647, 1.68335, 1.726959, 1.972015, 2.025513, 2.112183, 3.027161, 
    3.792175, 3.639648, 3.336212, 3.268494, 2.854431, 2.420105, 2.05072, 
    1.518494, 1.303558, 1.379883, 1.507233, 1.667633, 1.822449, 1.871307, 
    1.865234, 1.881561, 1.90683, 1.92981, 1.966553, 1.979431, 2.004608, 
    2.034576, 2.025665, 2.001495, 1.952606, 1.893341, 1.834961, 1.716095, 
    1.574951, 1.519867, 1.423187, 1.309845, 1.242767, 1.081909, 1.000153, 
    1.514648, 2.093964, 2.018677, 2.120636, 2.601379, 2.815369, 2.971283, 
    2.514954, 2.265228, 2.142853, 1.996033, 1.985413, 2.046356, 2.034576, 
    2.030487, 1.986511, 1.955719, 1.99765, 2.058807,
  1.880219, 1.806122, 1.768768, 1.797516, 1.898773, 3.098633, 3.765106, 
    3.884064, 3.908661, 2.23053, 1.995697, 1.997131, 1.889954, 1.717957, 
    1.639771, 1.733337, 1.785675, 1.73288, 1.691742, 1.7005, 1.862823, 
    2.016449, 2.098053, 2.206818, 2.329773, 2.433411, 2.515778, 2.555725, 
    2.423309, 1.954102, 1.69278, 1.858978, 2.007477, 2.009308, 2.248169, 
    2.395355, 2.304688, 2.169708, 2.338562, 2.38092, 2.548248, 2.779236, 
    2.648621, 2.762115, 2.775848, 2.62616, 2.213867, 1.779755, 1.538879, 
    1.397583, 1.523956, 1.724792, 1.859711, 1.906982, 1.960724, 1.997589, 
    1.989471, 2.008057, 2.009186, 2.027039, 2.045959, 2.028961, 2.028137, 
    2.04187, 2.036652, 1.959503, 1.825653, 1.684357, 1.547974, 1.376831, 
    1.252808, 1.21933, 1.132874, 1.060272, 1.02005, 0.9065552, 1.106567, 
    2.51767, 3.048309, 2.451904, 2.344086, 2.98114, 3.370178, 2.606445, 
    2.329346, 1.994537, 1.878967, 1.90567, 2.00885, 1.998962, 1.959717, 
    1.97467, 1.963867, 1.958221, 1.967682, 1.930298,
  1.679016, 1.643616, 1.76239, 1.974213, 2.497864, 4.022308, 4.659302, 
    4.174713, 3.904236, 2.374878, 2.098694, 2.197937, 2.216736, 2.172943, 
    2.23288, 2.393433, 2.446472, 2.391602, 2.387451, 2.418427, 2.436829, 
    2.453552, 2.463745, 2.436462, 2.39621, 2.322388, 2.233795, 2.115173, 
    2.013885, 1.927216, 1.871155, 2.357819, 2.270264, 2.318237, 2.319611, 
    2.381073, 2.495972, 2.31955, 2.170349, 2.643799, 3.039429, 2.242584, 
    1.899414, 1.893951, 1.967896, 1.978119, 1.992859, 1.984131, 2.002258, 
    2.045898, 2.049225, 1.98587, 1.939331, 1.914337, 1.928802, 1.912445, 
    1.870697, 1.875183, 1.911652, 1.951447, 1.941193, 1.916412, 1.875519, 
    1.870514, 1.863342, 1.732544, 1.572784, 1.386719, 1.214935, 1.074677, 
    1.003632, 0.9882813, 0.9535828, 0.8786011, 0.7873535, 0.885498, 1.65033, 
    3.346344, 3.592682, 2.96347, 2.726044, 3.548828, 3.772339, 3.349365, 
    2.420319, 2.028778, 1.907623, 1.994202, 1.973328, 1.91687, 1.912781, 
    1.905334, 1.902618, 1.871307, 1.789581, 1.727356,
  1.744781, 1.914337, 2.1698, 2.635559, 4.175446, 4.587128, 5.069153, 
    5.028046, 4.396759, 4.043243, 2.248718, 2.279633, 3.383606, 2.339722, 
    2.327209, 2.42691, 2.380127, 2.333618, 2.293365, 2.300781, 2.250275, 
    2.176636, 2.12854, 2.076813, 2.055023, 2.044586, 2.055725, 2.083008, 
    2.069427, 2.100708, 2.113464, 2.473694, 2.5289, 2.56366, 2.54422, 
    2.319794, 2.360443, 2.349213, 2.725586, 2.933197, 2.887024, 2.084595, 
    2.083923, 2.239502, 2.28595, 2.242859, 2.201996, 2.184235, 2.164581, 
    2.066071, 1.983856, 1.920319, 1.873138, 1.81192, 1.785797, 1.797211, 
    1.825592, 1.861145, 1.879669, 1.919006, 1.933319, 1.900909, 1.849274, 
    1.794342, 1.684967, 1.49231, 1.338287, 1.180664, 1.0755, 1.011169, 
    1.004944, 0.9602356, 0.8969421, 0.8147888, 0.9334412, 1.353638, 2.273193, 
    3.873688, 4.231506, 3.503113, 3.372223, 4.047913, 4.453766, 3.31958, 
    3.141235, 2.234161, 1.897064, 1.908936, 1.924164, 1.872131, 1.85321, 
    1.792358, 1.713409, 1.651245, 1.610748, 1.657806,
  2.055573, 2.350128, 2.504578, 2.838409, 4.626312, 4.457153, 4.567566, 
    4.610809, 4.018097, 3.717529, 2.361267, 2.45694, 3.35202, 2.882874, 
    2.246887, 2.255676, 2.155792, 2.156311, 2.1651, 2.166809, 2.176819, 
    2.174103, 2.169342, 2.166351, 2.230194, 2.323059, 2.373505, 2.322174, 
    2.262238, 2.282227, 2.290833, 2.254883, 2.940216, 3.09552, 2.87442, 
    2.690826, 2.681, 2.983856, 3.315735, 2.985413, 2.251312, 2.397125, 
    2.539063, 2.61673, 2.546356, 2.43576, 2.319336, 2.241669, 2.148682, 
    1.986328, 1.927338, 1.923889, 1.875458, 1.841278, 1.899353, 1.958527, 
    1.974091, 2.006714, 2.011627, 2.052429, 2.058411, 2.024536, 1.9328, 
    1.806305, 1.665436, 1.506714, 1.414276, 1.270264, 1.204559, 1.157227, 
    1.112244, 1.079865, 1.043427, 1.203278, 1.449066, 1.702087, 2.500824, 
    4.448517, 3.743439, 3.635223, 3.940765, 4.879547, 4.943359, 3.863281, 
    3.388153, 3.221344, 1.97467, 1.960632, 1.930542, 1.872681, 1.809174, 
    1.75885, 1.744904, 1.767395, 1.815369, 1.885864,
  2.532227, 2.622925, 2.584717, 2.725067, 4.575439, 4.278198, 3.995209, 
    4.173584, 4.016602, 3.623383, 3.429291, 2.518768, 3.26062, 3.069458, 
    2.107178, 2.088165, 2.068054, 2.099609, 2.163666, 2.238678, 2.270233, 
    2.298645, 2.33725, 2.381622, 2.430817, 2.450836, 2.417572, 2.385864, 
    2.398376, 2.456573, 2.517914, 2.467957, 2.571747, 3.874237, 3.696228, 
    3.476166, 3.023834, 2.656708, 3.137238, 2.422394, 2.532928, 2.765106, 
    2.770386, 2.719727, 2.592194, 2.442261, 2.313812, 2.192688, 2.092194, 
    2.002289, 1.991272, 1.977264, 1.98053, 2.021027, 2.076447, 2.136261, 
    2.130127, 2.168488, 2.172791, 2.187317, 2.179108, 2.149811, 2.077667, 
    1.978058, 1.936462, 1.888519, 1.852997, 1.795441, 1.763062, 1.743744, 
    1.656464, 1.717926, 1.836639, 1.950714, 1.932465, 2.20108, 4.210236, 
    4.613739, 3.566406, 3.786591, 4.485413, 4.48465, 4.43866, 4.084045, 
    3.657104, 2.928711, 2.02005, 2.108856, 2.096344, 2.09552, 2.093231, 
    2.149506, 2.197479, 2.238739, 2.301819, 2.363007,
  2.670135, 2.583588, 2.578125, 2.616486, 3.976959, 4.036865, 3.65332, 
    3.808136, 3.810852, 3.531891, 3.494476, 2.447388, 2.235809, 2.133514, 
    2.065094, 2.085876, 2.087891, 2.157104, 2.203644, 2.302643, 2.302338, 
    2.364105, 2.359161, 2.407349, 2.422852, 2.365356, 2.403961, 2.424957, 
    2.439453, 2.53183, 2.66803, 2.731842, 2.784119, 2.849365, 2.851959, 
    3.738922, 3.627808, 2.659637, 3.233002, 2.491669, 2.667267, 2.764709, 
    2.6651, 2.529541, 2.421082, 2.263733, 2.169189, 2.0867, 2.046539, 
    2.05011, 2.028442, 2.033203, 2.072388, 2.118561, 2.145447, 2.199615, 
    2.242584, 2.287292, 2.286926, 2.296234, 2.31543, 2.289917, 2.244781, 
    2.202393, 2.218933, 2.188538, 2.163879, 2.173126, 2.159058, 2.148712, 
    2.179626, 2.266052, 2.316284, 2.238678, 2.295227, 3.841125, 4.401489, 
    3.678192, 3.608673, 4.912292, 4.58667, 4.534058, 4.526428, 3.932281, 
    3.436005, 2.856903, 2.056335, 2.177002, 2.192078, 2.24115, 2.309631, 
    2.371155, 2.415436, 2.512299, 2.554504, 2.649628,
  2.551636, 2.5578, 2.578705, 2.484955, 3.786713, 3.956207, 3.511993, 
    3.577911, 3.568878, 3.366425, 3.040619, 2.365814, 2.153137, 2.103851, 
    2.116943, 2.204681, 2.192963, 2.277802, 2.347992, 2.396942, 2.40274, 
    2.442719, 2.451233, 2.486908, 2.432281, 2.390442, 2.396179, 2.396545, 
    2.446228, 2.494141, 2.592316, 2.642639, 2.653961, 2.649689, 2.579956, 
    2.538269, 2.489258, 2.44162, 2.84433, 2.486847, 2.573181, 2.539337, 
    2.477081, 2.367004, 2.236969, 2.117645, 2.053528, 2.033661, 2.012054, 
    2.048645, 2.050049, 2.082336, 2.080536, 2.103638, 2.124481, 2.156311, 
    2.193817, 2.228577, 2.270142, 2.300446, 2.336456, 2.319977, 2.328003, 
    2.345978, 2.336792, 2.359833, 2.397156, 2.403931, 2.419128, 2.412384, 
    2.448181, 2.402588, 2.432159, 2.408997, 2.404755, 3.805756, 3.767334, 
    4.5961, 4.620728, 4.736511, 4.311676, 4.601959, 4.07016, 3.445374, 
    2.92926, 2.926636, 2.710999, 2.23288, 2.23761, 2.324982, 2.389587, 
    2.429749, 2.472137, 2.556183, 2.580414, 2.586548,
  2.539185, 2.742004, 2.833771, 2.959442, 4.315094, 4.191406, 3.766449, 
    3.5242, 3.196045, 2.300385, 2.432098, 2.274933, 2.213531, 2.219482, 
    2.26062, 2.30304, 2.351746, 2.437164, 2.489014, 2.487701, 2.482147, 
    2.476868, 2.465942, 2.503174, 2.450775, 2.459503, 2.390045, 2.389252, 
    2.679596, 2.479797, 2.465363, 2.502533, 2.51178, 2.505035, 2.601105, 
    2.392914, 2.234314, 2.274017, 2.826782, 2.911224, 2.579376, 2.382935, 
    2.27948, 2.187561, 2.069458, 2.032043, 1.991089, 1.943665, 1.927338, 
    1.948242, 1.967773, 2.039856, 2.111847, 2.173767, 2.2117, 2.273804, 
    2.31308, 2.344391, 2.367004, 2.38736, 2.40033, 2.398193, 2.386475, 
    2.363983, 2.356171, 2.382751, 2.395966, 2.397522, 2.440247, 2.40332, 
    2.396545, 2.350922, 2.423492, 2.43808, 2.351105, 3.791351, 4.492462, 
    3.977753, 3.821747, 4.074951, 4.286316, 3.964966, 3.758331, 3.556122, 
    3.407654, 3.045776, 2.816925, 2.226807, 2.225861, 2.367584, 2.433258, 
    2.475586, 2.547913, 2.590576, 2.5784, 2.540558,
  2.762909, 2.878448, 2.918121, 3.817902, 4.139771, 3.543793, 3.327271, 
    3.231842, 3.025635, 1.634888, 2.265747, 3.476044, 2.262634, 2.231689, 
    2.382355, 2.34082, 2.409515, 2.478699, 2.4664, 2.377014, 2.341217, 
    2.351929, 2.366028, 2.42337, 2.433075, 2.408478, 2.328766, 2.903137, 
    2.755341, 2.419922, 2.953125, 2.8078, 2.734497, 2.372314, 2.464172, 
    2.642181, 2.509827, 2.292084, 2.659241, 2.459198, 2.498505, 2.30777, 
    2.178253, 2.117859, 2.058746, 2.07251, 2.033142, 1.980988, 1.957031, 
    2.015564, 2.135345, 2.323242, 2.534973, 2.686188, 2.786926, 2.81192, 
    2.782959, 2.739777, 2.638947, 2.544342, 2.439362, 2.360199, 2.297485, 
    2.26297, 2.289917, 2.2901, 2.325714, 2.348694, 2.377747, 2.395599, 
    2.366333, 2.321136, 2.3367, 2.310028, 2.265411, 3.328888, 4.054321, 
    3.486115, 3.198425, 3.884827, 3.354095, 3.500977, 3.921539, 3.419159, 
    3.305725, 2.450714, 2.229218, 2.300323, 2.305145, 2.452942, 2.492645, 
    2.546082, 2.633942, 2.653259, 2.637756, 2.636902,
  2.520325, 2.679291, 2.628265, 3.041473, 2.884613, 2.797394, 2.999603, 
    2.996399, 3.11673, 2.793091, 2.618347, 3.447723, 3.375702, 2.229828, 
    2.422607, 2.446808, 2.397247, 2.385864, 2.320465, 2.248291, 2.211395, 
    2.214325, 2.205841, 2.32663, 2.402008, 2.298767, 2.306183, 2.655548, 
    2.367767, 2.314575, 3.043579, 2.291992, 2.177277, 2.186005, 2.133667, 
    2.065704, 2.00116, 2.030334, 2.196228, 2.335815, 2.320648, 2.209045, 
    2.141541, 2.105011, 2.095306, 2.090485, 2.073883, 2.033203, 2.04837, 
    2.120514, 2.211517, 2.385742, 2.571686, 2.7323, 2.829163, 2.869354, 
    2.847321, 2.808136, 2.742462, 2.624146, 2.514587, 2.4216, 2.352844, 
    2.309509, 2.284576, 2.264099, 2.276276, 2.27774, 2.27359, 2.253967, 
    2.14621, 2.062317, 1.947968, 1.91037, 1.881775, 2.486725, 3.102722, 
    3.079559, 2.892059, 3.259766, 3.047638, 3.454285, 3.45932, 2.51413, 
    2.431427, 2.43573, 2.323395, 2.275757, 2.217255, 2.280151, 2.390228, 
    2.442657, 2.486908, 2.493103, 2.439575, 2.412354,
  2.713348, 2.638428, 2.698639, 2.719971, 2.624603, 2.579285, 2.744995, 
    2.770508, 2.917511, 3.142303, 2.878571, 2.882813, 3.426575, 2.388947, 
    2.271301, 2.408539, 2.361847, 2.498291, 2.479095, 2.407379, 2.318939, 
    2.229858, 2.208862, 2.413239, 2.422943, 2.30899, 2.989441, 2.428009, 
    2.282745, 2.258728, 2.326996, 2.482361, 2.037476, 2.189514, 2.177094, 
    2.115021, 2.137634, 2.152527, 2.137299, 2.126343, 2.184631, 2.227142, 
    2.241608, 2.211639, 2.198578, 2.186127, 2.212769, 2.190887, 2.18219, 
    2.192169, 2.157227, 2.125519, 2.12207, 2.12851, 2.140045, 2.173248, 
    2.16217, 2.163605, 2.194336, 2.191406, 2.261902, 2.302155, 2.317383, 
    2.357025, 2.30014, 2.309967, 2.250061, 2.274017, 2.231171, 2.13501, 
    2.040619, 1.929901, 1.776703, 1.847321, 2.024292, 2.564178, 2.653046, 
    2.900146, 3.434387, 3.714386, 3.961761, 3.953674, 2.62558, 2.17746, 
    2.319458, 2.347412, 2.397919, 2.420624, 2.418243, 2.428528, 2.452972, 
    2.397125, 2.316223, 2.31604, 2.803528, 2.897705,
  2.719635, 2.805359, 2.862183, 2.925934, 2.758331, 2.683655, 2.677094, 
    2.739258, 2.933258, 3.377869, 3.240173, 3.319611, 3.392456, 2.967773, 
    2.45105, 2.417114, 2.273376, 2.350464, 2.528717, 2.489532, 2.424408, 
    2.279633, 2.420959, 2.32547, 2.350769, 2.355194, 2.460815, 2.195313, 
    2.5047, 2.436249, 2.455536, 2.354126, 2.235077, 2.300323, 2.205597, 
    2.154572, 2.146332, 2.127563, 2.129364, 2.168427, 2.256531, 2.303833, 
    2.282349, 2.28363, 2.313141, 2.250641, 2.259583, 2.296478, 2.264435, 
    2.26828, 2.264313, 2.244934, 2.230621, 2.197998, 2.191071, 2.15976, 
    2.122467, 2.087646, 2.061798, 2.072784, 2.101868, 2.155151, 2.16391, 
    2.187317, 2.203857, 2.259552, 2.324738, 2.501373, 2.55896, 2.550385, 
    2.389587, 2.25351, 2.250153, 2.099152, 2.621948, 2.650696, 2.961395, 
    3.731964, 4.963135, 3.784943, 2.363342, 2.387238, 2.326599, 2.248199, 
    2.226105, 2.255981, 2.330536, 2.374084, 2.440765, 2.456299, 2.479034, 
    2.358582, 2.38797, 2.869598, 2.926605, 2.97168,
  2.864014, 2.811218, 2.600372, 2.767395, 2.943359, 3.352478, 3.75412, 
    3.333801, 2.890686, 3.417389, 4.139923, 4.430664, 4.191803, 3.546417, 
    2.352173, 2.221039, 2.270691, 2.286133, 2.415222, 2.376953, 2.495941, 
    2.027802, 2.182159, 2.185181, 2.250916, 2.288757, 2.440033, 2.971527, 
    2.907684, 2.422272, 2.482697, 2.433319, 2.349091, 2.27417, 2.138672, 
    2.117188, 2.103516, 2.099792, 2.139801, 2.160034, 2.1828, 2.168671, 
    2.204834, 2.228729, 2.285614, 2.284363, 2.28064, 2.31958, 2.316071, 
    2.308838, 2.307739, 2.278931, 2.282288, 2.297516, 2.285858, 2.278442, 
    2.259979, 2.273438, 2.276306, 2.333649, 2.346008, 2.354828, 2.300781, 
    2.278198, 2.277161, 2.332611, 2.525909, 2.737061, 2.814728, 2.774292, 
    2.597992, 2.703644, 4.582703, 3.786652, 2.00827, 2.101166, 2.245697, 
    2.21048, 2.219604, 2.253143, 2.220978, 2.188477, 2.088623, 2.087006, 
    2.092255, 2.148895, 2.159393, 2.242981, 2.254669, 2.378326, 2.395386, 
    2.315277, 3.950409, 4.74942, 3.932037, 2.940948,
  3.523254, 4.121277, 3.845032, 3.773773, 3.671661, 3.591553, 3.381531, 
    3.237061, 3.29068, 3.453003, 3.612244, 3.791229, 4.412262, 4.634766, 
    3.117889, 2.194336, 2.311584, 2.262238, 2.33255, 2.328125, 2.409637, 
    2.24649, 2.313202, 2.337372, 2.255585, 2.272675, 2.736206, 3.136108, 
    2.738739, 2.276642, 2.300079, 2.563416, 2.433441, 2.091797, 2.069794, 
    2.124878, 2.067505, 2.080017, 2.15683, 2.177734, 2.137634, 2.09668, 
    2.156311, 2.213593, 2.260498, 2.299347, 2.341248, 2.313599, 2.306488, 
    2.321869, 2.309814, 2.31427, 2.301422, 2.305145, 2.244781, 2.248566, 
    2.220093, 2.231323, 2.28772, 2.330933, 2.368683, 2.455658, 2.415436, 
    2.267212, 2.108459, 2.027466, 2.17511, 2.532074, 2.737671, 2.844086, 
    3.576233, 5.054047, 4.418671, 2.065369, 2.061401, 2.148254, 2.127289, 
    2.074921, 2.039063, 2.104736, 2.113464, 2.031311, 2.012939, 2.081451, 
    2.073578, 2.032928, 2.004822, 2.056641, 2.066345, 2.241211, 2.278076, 
    2.278198, 4.074158, 5.839447, 4.988464, 3.635406,
  3.869324, 3.974091, 4.115448, 3.835999, 3.729431, 3.45105, 3.474365, 
    3.443512, 3.585236, 3.519592, 2.337952, 3.612823, 4.425446, 4.091858, 
    3.562408, 2.204346, 2.140411, 2.41153, 2.472565, 2.338562, 1.996185, 
    2.623169, 2.714508, 2.684845, 2.412109, 2.429993, 2.346344, 2.624878, 
    2.627167, 2.297058, 2.116852, 2.348969, 2.380737, 2.224945, 2.183807, 
    2.183655, 2.135864, 2.156097, 2.180237, 2.164276, 2.132294, 2.132233, 
    2.112244, 2.103516, 2.105591, 2.116028, 2.158325, 2.155701, 2.168243, 
    2.17749, 2.172729, 2.182922, 2.156342, 2.194672, 2.146484, 2.102844, 
    2.087494, 2.062958, 2.052429, 2.096008, 2.099792, 2.151947, 2.124237, 
    1.987885, 1.732544, 1.304291, 1.406586, 2.282104, 2.894989, 3.043701, 
    4.316345, 5.567261, 3.654144, 2.162903, 2.275726, 2.188202, 2.08548, 
    2.025848, 2.004944, 1.982544, 1.998352, 2.044647, 2.053192, 2.024994, 
    1.986206, 1.996338, 1.940125, 1.89447, 1.869751, 1.939758, 2.026306, 
    2.264984, 4.292847, 5.798615, 5.597931, 4.674622,
  4.52655, 4.352875, 4.043549, 3.842438, 3.43985, 3.197845, 3.360626, 
    3.346741, 3.455994, 3.601105, 2.480927, 3.949158, 4.678497, 3.971039, 
    3.422455, 2.329712, 2.169403, 2.361786, 1.628204, 1.538727, 1.6651, 
    2.31015, 2.444275, 2.286987, 2.430267, 2.012878, 1.992493, 2.802551, 
    2.815247, 2.371552, 2.197113, 2.51355, 2.329834, 2.352814, 2.314056, 
    2.310669, 2.296631, 2.207764, 2.204254, 2.203461, 2.184784, 2.131836, 
    2.085663, 2.045715, 2.0112, 1.997772, 1.984375, 1.956299, 1.968292, 
    1.985809, 2.00827, 2.005432, 1.961395, 1.92688, 1.930969, 1.934967, 
    1.920898, 1.925476, 1.878662, 1.907959, 1.914673, 1.904938, 1.942902, 
    1.854889, 1.652618, 1.224762, 1.757599, 5.081329, 4.106659, 3.020386, 
    2.668884, 2.215759, 1.904144, 2.139435, 2.188416, 2.022461, 1.967773, 
    2.033478, 2.19754, 2.203125, 2.174866, 2.179321, 2.146484, 2.169525, 
    2.134308, 2.079956, 2.008667, 1.972076, 1.911255, 1.891846, 1.786346, 
    2.195313, 3.952789, 5.275116, 5.231384, 4.911438,
  4.975311, 4.431244, 3.920135, 3.429749, 3.048615, 2.842896, 3.357941, 
    3.536407, 3.30658, 3.467957, 3.825653, 4.501129, 4.621033, 4.316528, 
    4.472992, 4.115173, 3.879242, 3.187897, 1.370636, 0.5042725, 1.046295, 
    1.921539, 2.365936, 2.728851, 2.933685, 2.74469, 2.42572, 2.891663, 
    3.102875, 2.81543, 2.876434, 2.988342, 2.921265, 2.495911, 2.451263, 
    2.480713, 2.418274, 2.352081, 2.332214, 2.268372, 2.194275, 2.09668, 
    2.084045, 2.111969, 2.11499, 2.08078, 2.00592, 1.928558, 1.85965, 
    1.829559, 1.909882, 2.003693, 2.025574, 2.006775, 1.956787, 1.926697, 
    1.861481, 1.872406, 1.820831, 1.828308, 1.857025, 1.853607, 1.903381, 
    1.697327, 1.471039, 1.685486, 3.354431, 4.584076, 3.187775, 1.629425, 
    1.774597, 2.30365, 2.430939, 2.565186, 2.570313, 1.953003, 1.949982, 
    2.127747, 2.257629, 2.194916, 2.189972, 2.240692, 2.287628, 2.304291, 
    2.260498, 2.211121, 2.1745, 2.087708, 2.012756, 1.966736, 1.801178, 
    1.761383, 2.396484, 4.292206, 5.275635, 5.407043,
  5.861328, 5.411072, 4.542053, 3.542389, 2.834229, 2.368622, 3.379425, 
    3.427368, 2.50415, 3.105988, 4.028168, 4.272522, 4.264465, 4.707367, 
    4.921661, 4.967834, 4.542633, 4.113983, 3.689728, 1.871765, 1.705383, 
    2.691162, 4.320496, 3.313171, 3.684296, 3.399139, 3.040436, 3.516754, 
    3.681641, 3.244781, 3.000397, 3.022003, 3.213043, 2.46106, 2.345978, 
    2.440338, 2.393158, 2.347656, 2.282623, 2.28125, 2.378052, 2.320129, 
    2.275757, 2.271088, 2.277161, 2.303131, 2.236603, 2.156708, 2.079163, 
    2.0224, 2.080719, 2.117767, 2.167206, 2.198853, 2.171356, 2.109314, 
    2.01886, 1.924011, 1.832581, 1.819733, 1.855316, 1.816284, 1.734161, 
    1.564453, 1.713593, 2.700439, 3.686279, 3.47995, 1.851563, 1.491669, 
    2.542328, 3.38266, 3.728058, 3.466187, 3.037048, 2.201752, 1.899017, 
    1.956329, 2.060028, 2.117645, 2.190826, 2.164978, 2.070831, 2.040375, 
    2.101501, 2.15918, 2.172729, 2.143402, 2.136047, 2.076294, 1.994263, 
    1.869324, 1.808319, 2.471985, 4.436676, 5.659515,
  5.993225, 5.972565, 5.135803, 2.842896, 2.250275, 2.312836, 2.741394, 
    2.788483, 2.801056, 2.956329, 4.140991, 4.392975, 4.654358, 4.953033, 
    4.965027, 4.921692, 4.515411, 4.430542, 4.519073, 4.531189, 4.26062, 
    4.998688, 4.964752, 4.080933, 4.192017, 3.976379, 3.487976, 3.6875, 
    3.55722, 3.056122, 2.838348, 2.601257, 2.655853, 2.57428, 2.594666, 
    2.776825, 2.808777, 2.618896, 2.364655, 2.351837, 2.388214, 2.324921, 
    2.338654, 2.41452, 2.430084, 2.405273, 2.374634, 2.37851, 2.361664, 
    2.326874, 2.354218, 2.35434, 2.346375, 2.358734, 2.371368, 2.355225, 
    2.262573, 2.142395, 1.968384, 1.871552, 1.874146, 1.77597, 1.786865, 
    2.114075, 3.629028, 4.177155, 4.188812, 3.894623, 3.297638, 2.266876, 
    2.589844, 3.357208, 4.20282, 3.624603, 2.908203, 2.497528, 2.32312, 
    2.144989, 1.985168, 2.0047, 2.008392, 2.00885, 1.987091, 1.866333, 
    1.696411, 1.486511, 1.584442, 1.881897, 2.081512, 2.109955, 2.112701, 
    2.073303, 1.827667, 1.988983, 2.753387, 5.164795,
  5.117981, 2.56073, 2.569214, 2.703796, 2.676575, 3.082306, 5.190033, 
    4.833527, 4.801575, 5.055817, 4.702942, 4.72644, 4.68457, 4.192444, 
    2.739838, 4.169006, 4.265167, 3.865417, 3.992584, 4.772125, 5.418213, 
    4.674622, 4.486176, 4.230286, 4.405853, 4.276581, 3.694275, 3.53302, 
    3.074677, 2.674805, 2.718475, 2.618347, 2.484283, 2.562042, 2.781311, 
    2.978119, 2.792725, 2.657959, 2.512115, 2.503143, 2.545685, 2.598114, 
    2.602295, 2.626312, 2.682495, 2.657013, 2.582428, 2.563171, 2.567535, 
    2.550781, 2.492188, 2.452393, 2.397278, 2.311249, 2.293091, 2.266937, 
    2.212189, 2.164642, 1.996429, 1.856903, 1.872528, 1.776764, 2.180725, 
    3.966217, 5.179321, 4.574219, 3.753448, 3.958069, 3.805481, 3.308716, 
    3.354492, 3.6026, 3.451019, 3.019806, 2.654236, 2.765411, 3.026154, 
    2.926819, 2.542725, 2.248169, 2.203247, 2.306824, 2.237549, 1.84967, 
    1.314392, 0.6134644, 0.3781738, 0.8864746, 1.417908, 1.786652, 2.023102, 
    1.978516, 1.967834, 2.643677, 5.227234, 6.238647,
  4.440613, 2.497009, 2.974762, 5.234436, 3.018188, 4.600128, 4.348297, 
    3.898438, 3.766418, 3.161865, 3.30246, 3.008698, 3.233063, 2.399078, 
    3.071533, 3.273804, 3.509491, 3.188873, 3.294617, 3.634979, 3.954773, 
    4.554565, 4.66629, 4.58905, 4.584839, 4.464844, 4.316162, 4.32605, 
    4.03183, 3.443939, 2.984497, 2.649872, 2.485352, 2.70575, 2.734253, 
    2.686676, 2.615112, 2.628387, 2.662567, 3.232422, 3.192535, 3.014252, 
    2.68692, 2.555725, 2.474884, 2.406982, 2.353119, 2.294342, 2.295197, 
    2.340637, 2.403717, 2.370819, 2.289398, 2.183868, 2.133148, 2.141724, 
    2.129303, 2.051758, 1.900909, 1.901825, 1.898743, 1.757813, 2.106323, 
    4.152008, 4.880066, 4.501038, 3.664764, 3.918091, 3.613403, 3.205078, 
    3.458008, 3.48941, 3.18158, 3.271545, 3.433411, 3.644989, 3.693237, 
    3.859497, 3.625153, 3.343109, 2.853149, 2.622406, 2.479095, 2.040955, 
    1.579376, 1.004028, 0.6270142, 0.708313, 0.9026184, 1.176392, 1.656708, 
    1.803528, 1.775146, 2.498749, 5.56543, 5.715485,
  3.850128, 3.875854, 3.874481, 3.584229, 2.556976, 2.534241, 2.62735, 
    2.737823, 3.11499, 3.158081, 2.872131, 2.424683, 2.377411, 2.818573, 
    2.227753, 2.483521, 2.540802, 2.798431, 3.186768, 3.384155, 3.492065, 
    3.625122, 3.650116, 3.683716, 3.650696, 3.672974, 3.028564, 2.914764, 
    3.103394, 2.984375, 2.605927, 2.605865, 2.743835, 2.696442, 2.601105, 
    2.456238, 2.292603, 2.470306, 2.840576, 2.677429, 2.565308, 2.66745, 
    2.539856, 2.43985, 2.352997, 2.227936, 2.073242, 2.088867, 2.16275, 
    2.172668, 2.181976, 2.170227, 2.112885, 2.093811, 2.072601, 2.070435, 
    2.049103, 1.990021, 1.913879, 1.935303, 1.955139, 1.833191, 2.023712, 
    3.302673, 3.952026, 4.114655, 4.056122, 4.252014, 3.697601, 3.291718, 
    3.004211, 3.198486, 3.484253, 3.254089, 3.857819, 3.858398, 3.676086, 
    3.730347, 3.825562, 3.737244, 3.146027, 2.518616, 1.904968, 1.691284, 
    1.513672, 1.302216, 0.9184265, 0.6837769, 0.5253906, 0.4834595, 1.012878, 
    1.618286, 1.797211, 1.838776, 2.314514, 3.774078,
  3.217987, 3.387177, 3.129822, 2.695648, 2.056702, 2.00174, 1.923309, 
    2.216553, 2.464111, 2.750061, 2.475189, 1.906067, 1.941803, 2.23053, 
    2.483978, 2.631378, 2.517883, 2.526428, 2.593109, 2.477539, 2.750854, 
    3.065308, 3.071899, 3.057739, 3.5047, 3.204742, 3.058838, 2.671204, 
    2.7547, 2.507935, 2.421021, 2.407501, 2.475403, 2.229614, 2.239197, 
    2.396942, 2.249084, 2.071106, 1.863373, 2.38266, 2.813599, 2.814697, 
    2.645905, 2.485168, 2.461182, 2.417572, 2.337372, 2.266907, 2.257813, 
    2.204285, 2.148956, 2.117493, 2.155853, 2.233978, 2.302887, 2.308319, 
    2.21347, 2.112671, 2.020844, 1.951233, 1.8685, 1.922668, 2.67807, 
    3.10202, 3.190369, 3.448914, 4.191284, 4.494659, 4.378632, 4.062805, 
    3.678711, 3.589325, 3.619354, 3.802734, 3.848846, 3.82016, 3.693542, 
    3.536652, 3.550995, 3.588806, 3.035736, 3.244537, 2.183746, 2.144196, 
    1.781769, 1.279297, 0.5627747, -0.1034546, -0.3509216, -0.1983032, 
    0.3695984, 1.09494, 1.589447, 1.709625, 1.776245, 2.031067,
  2.698883, 1.976227, 2.544128, 2.57605, 2.579102, 2.456635, 1.957825, 
    1.581573, 1.829254, 1.906128, 1.95462, 1.779358, 1.491272, 1.344025, 
    1.28653, 1.241425, 1.811737, 2.390808, 2.795959, 3.020203, 3.096222, 
    3.110992, 3.158325, 3.157959, 3.099426, 2.984222, 2.659637, 2.744263, 
    2.942444, 2.948242, 3.358856, 3.202667, 2.824921, 2.522644, 2.786072, 
    2.851624, 2.516144, 2.177155, 1.700653, 2.239014, 2.960693, 3.101746, 
    3.073059, 2.392517, 2.437714, 2.40799, 2.379425, 2.349213, 2.308075, 
    2.277069, 2.323517, 2.419403, 2.468597, 2.509399, 2.522339, 2.474091, 
    2.341583, 2.2117, 2.077728, 1.951233, 1.805725, 2.161652, 2.489716, 
    2.846741, 2.899109, 3.028168, 3.209961, 3.450836, 3.44278, 3.343353, 
    3.240875, 3.401764, 3.467773, 3.755188, 4.264038, 2.921936, 3.448761, 
    3.308899, 3.486206, 3.664459, 3.365295, 1.983246, 1.774475, 1.555267, 
    1.185822, 1.058014, 0.663269, -0.1086731, -0.6504517, -0.5123596, 
    0.138092, 0.8434143, 1.333008, 1.591919, 2.187256, 2.578369,
  1.439545, 1.50885, 1.288788, 2.063873, 2.400848, 2.397797, 1.913208, 
    1.594147, 1.738647, 1.77597, 1.680145, 1.701477, 1.482178, 1.249207, 
    1.214111, 1.515747, 1.940826, 2.702667, 3.300507, 3.613617, 3.828003, 
    3.831757, 3.863617, 3.742432, 3.287323, 2.692139, 2.675537, 2.868561, 
    3.042511, 3.357025, 3.571106, 3.550537, 3.336914, 3.318512, 3.471222, 
    3.298645, 2.945831, 2.685791, 1.789246, 1.810944, 1.961456, 1.917114, 
    3.204956, 3.289215, 2.061523, 2.41687, 2.627197, 2.836517, 3.009827, 
    3.144989, 3.259705, 3.194855, 2.998962, 2.814697, 2.690033, 2.400513, 
    2.318726, 2.224548, 2.114319, 1.897278, 2.270966, 2.537292, 2.948547, 
    2.920685, 2.706696, 2.831787, 2.892517, 2.840881, 3.010742, 3.064789, 
    3.084625, 3.248962, 1.781189, 1.634521, 1.794525, 2.088623, 2.97937, 
    3.272278, 3.37674, 3.165863, 1.741272, 1.47876, 1.063843, 0.5244751, 
    0.5201111, 0.9404297, 1.019409, 0.7524109, 0.3791809, 0.3467712, 
    0.6171875, 0.9226074, 1.124329, 1.253845, 1.466064, 2.011444,
  0.8901062, 1.038086, 1.645386, 2.039215, 2.157471, 1.550385, 1.971497, 
    1.820496, 1.958801, 1.994843, 2.141144, 2.280396, 2.442261, 2.651825, 
    2.869263, 3.189575, 3.740021, 4.295319, 4.724792, 4.749237, 4.717773, 
    4.413513, 4.390961, 4.270233, 3.961731, 4.128906, 3.686401, 3.455017, 
    3.342194, 3.300262, 3.140106, 2.921356, 2.7948, 2.758636, 2.745422, 
    2.863434, 2.9599, 2.973419, 2.685486, 2.68573, 2.857605, 2.968811, 
    3.474365, 3.402924, 3.481323, 3.362488, 3.467773, 2.482666, 2.764648, 
    3.02655, 3.096008, 2.926941, 2.832092, 2.656647, 2.580719, 2.78717, 
    3.182617, 4.026764, 4.025208, 3.705353, 3.647278, 3.695557, 3.497681, 
    3.173767, 2.574493, 2.504822, 2.712036, 2.765625, 2.742767, 2.750061, 
    2.597931, 2.008209, 1.909698, 1.498718, 1.225403, 1.1586, 2.303589, 
    2.468506, 1.218109, 1.32193, 1.208221, 0.9768677, 0.7662659, 0.4697266, 
    0.4057312, 0.2389832, 0.3777466, 0.6996155, 0.9581299, 1.07547, 1.103638, 
    0.8674622, 0.4921875, 0.4130859, 0.7339783, 0.8890076,
  0.3127136, 0.3846741, 0.6375427, 1.475586, 1.567566, 1.648773, 1.061005, 
    2.119202, 2.3508, 2.478729, 2.532013, 2.674408, 2.966339, 3.308868, 
    3.536469, 3.737366, 4.152435, 4.662354, 4.867828, 4.933014, 4.759064, 
    4.615173, 4.408203, 4.257355, 4.391388, 4.459442, 4.264008, 3.769928, 
    3.173248, 3.126495, 2.735413, 2.831635, 2.733795, 2.549957, 2.789459, 
    2.94635, 2.333282, 2.383331, 2.022522, 1.966675, 2.698639, 2.343384, 
    2.600647, 2.566864, 2.272217, 2.186462, 2.471344, 2.725128, 2.565491, 
    2.854034, 2.76651, 2.500519, 2.613953, 2.693878, 2.88028, 3.132874, 
    3.376953, 3.564117, 3.537231, 3.469452, 3.331573, 3.282379, 2.789703, 
    2.300995, 2.455811, 2.807434, 2.970184, 2.988281, 2.816406, 2.326508, 
    2.340698, 2.725739, 2.84082, 2.511078, 0.5821533, 0.7887573, 1.041321, 
    1.958771, 1.952728, 1.54068, 0.9759216, 0.8684082, 1.336975, 1.454773, 
    1.685364, 1.458984, 0.7946167, 0.6294861, 0.6238708, 0.9335022, 1.066559, 
    1.31842, 0.9282532, 0.3959656, 0.136261, 0.07427979,
  0.5612183, 0.5365906, 0.4850464, 0.2998657, -0.02441406, 1.389771, 
    1.918091, 2.427094, 2.803711, 2.943695, 2.903381, 2.013031, 2.02356, 
    2.126617, 3.576233, 3.711151, 4.061005, 4.311523, 4.633972, 4.941589, 
    5.069336, 4.95813, 4.7771, 4.569122, 4.285156, 3.786926, 3.561005, 
    3.713013, 3.608002, 3.4823, 3.180023, 2.932037, 2.706116, 2.649994, 
    2.089661, 2.164581, 2.353912, 1.876221, 1.636597, 1.155273, 0.538147, 
    0.3616333, 0.1906433, 0.2266541, 0.6664124, 0.9206848, 1.094727, 
    1.413727, 1.700653, 0.4614563, 0.7635498, 1.217438, 1.438293, 2.128967, 
    2.339478, 2.489471, 2.414398, 2.219147, 2.278381, 1.762695, 1.277802, 
    1.020294, 0.9492188, 1.434113, 2.115875, 2.73056, 3.427551, 3.298828, 
    2.993866, 1.648376, 2.514984, 2.474152, 2.332886, 0.8902283, 1.916351, 
    0.4662781, 1.784698, 1.787842, 1.161285, 0.3115234, 0.6384277, 0.8151855, 
    1.2388, 2.699097, 2.874756, 3.075623, 2.807251, 2.519531, 2.197601, 
    1.651245, 1.229431, 1.324341, 1.018494, 0.9809265, 0.8881531, 0.7484131,
  1.51355, 1.341797, 1.08197, 0.8447876, 0.6324158, 0.9013672, 1.680664, 
    2.267944, 2.397308, 2.296692, 2.072723, 1.961639, 1.867889, 1.706757, 
    1.399811, 2.017181, 0.8376465, 0.8947144, 0.9639587, 3.627167, 4.352539, 
    4.386658, 4.316803, 4.243256, 4.161469, 4.127075, 4.012451, 4.055878, 
    4.066528, 3.708862, 3.571869, 3.063263, 2.582153, 2.159363, 1.808472, 
    0.4347534, 0.4810486, 0.5532532, 1.831055, 1.665771, 0.2625122, 
    0.2036438, 0.15625, 0.1540222, 0.1553955, 0.1705627, 0.2061157, 0.210022, 
    0.2121277, 0.2208557, 0.2085876, 0.1899719, 0.1568909, 0.1586609, 
    0.1708374, 0.1806641, 0.2133484, 0.2169495, 0.2080078, 0.1587219, 
    0.2110596, 0.3679504, 0.6528015, 2.313995, 2.847534, 3.202362, 3.517212, 
    3.443359, 3.15918, 1.493866, 2.002197, 1.638611, 0.7561035, 1.690369, 
    1.874664, 2.722382, 1.66095, 0.5757141, 0.3772583, 0.4113464, 0.6968689, 
    1.336456, 2.901886, 3.371582, 3.618561, 3.465759, 3.320862, 3.176178, 
    2.999573, 2.757629, 2.007233, 0.5357361, 0.9477234, 1.167664, 1.285828, 
    1.463013,
  1.465759, 1.544159, 1.746613, 2.052155, 2.139465, 2.053711, 2.003815, 
    1.701904, 1.398712, 1.050537, 0.8057556, 0.6414795, 0.5319824, 0.3910217, 
    0.3045654, 0.308136, 0.3449402, 0.4195251, 0.4816589, 0.5389099, 
    0.6360779, 0.7453918, 0.8305969, 0.8903503, 1.088928, 2.519073, 2.547791, 
    2.769012, 2.681763, 2.329559, 2.029053, 0.5246582, 0.4689331, 0.3735657, 
    0.3339233, 0.3251953, 0.3471375, 0.3856201, 0.4299316, 0.4550781, 
    0.4597473, 0.4611511, 0.468689, 0.456604, 0.4270935, 0.4276123, 0.412384, 
    0.4267578, 0.433075, 0.4335938, 0.4253235, 0.4220886, 0.3929443, 
    0.3754272, 0.4011841, 0.433075, 0.481842, 0.5196838, 0.5151672, 
    0.4832764, 0.4215698, 0.3299561, 0.2570496, 0.2840576, 0.3411865, 
    1.492706, 1.669281, 1.685547, 1.792145, 2.007935, 1.995056, 0.8450317, 
    0.8979187, 1.051239, 1.433258, 0.1911316, 0.3716125, 0.4096069, 2.082062, 
    2.388824, 2.629578, 3.010162, 3.369873, 3.707001, 3.850494, 3.688019, 
    3.400787, 3.25, 2.986877, 2.664001, 2.330963, 1.414703, 0.2166138, 
    0.0916748, 0.4359436, 1.182434,
  0.3288574, 0.2875977, 0.3639526, 0.3862915, 1.316162, 1.294952, 1.260498, 
    0.406189, 0.4598999, 0.4867859, 0.4285278, 0.385437, 0.3296204, 
    0.3161316, 0.3566589, 0.3821106, 0.4286499, 0.454895, 0.4316101, 
    0.3827209, 0.3503418, 0.3300781, 0.3503418, 0.3681946, 0.4099731, 
    1.186157, 1.148254, 0.386261, 0.3632813, 0.3374939, 0.3266296, 0.3244019, 
    0.352417, 0.3492432, 0.3345337, 0.3270569, 0.3540649, 0.369812, 
    0.3812561, 0.3826599, 0.3778076, 0.3956604, 0.4006653, 0.416687, 
    0.4729309, 0.5170288, 0.5769653, 0.6427307, 0.6864929, 0.6941528, 
    0.6983337, 0.7376404, 0.7320251, 0.7168579, 0.6763306, 0.6802979, 
    0.7017822, 0.7159729, 0.7651672, 0.7734375, 0.8180542, 0.8522339, 
    0.8710022, 0.8933105, 0.9109497, 0.9041138, 0.870697, 0.7617798, 
    0.6539917, 0.5945435, 0.5379639, 1.554413, 2.483795, 1.798004, 1.966095, 
    2.147156, 2.28479, 2.481201, 2.704102, 2.92691, 3.053986, 3.208679, 
    3.348053, 3.405884, 3.440125, 3.453705, 3.37738, 3.212341, 2.96701, 
    2.705872, 2.392792, 2.081207, 0.6045532, 0.513092, 0.4386902, 0.3668213,
  0.9762573, 0.9598999, 0.9448547, 0.8901062, 0.8929138, 0.865448, 0.8268433, 
    0.7798462, 0.7329102, 0.6729736, 0.6230469, 0.5984497, 0.6004944, 
    0.612793, 0.6190186, 0.6080322, 0.5895996, 0.5806885, 0.5506592, 
    0.5247803, 0.492218, 0.4666748, 0.4273682, 0.3809509, 0.3587341, 
    0.3381653, 0.3179626, 0.3132324, 0.3051453, 0.3165894, 0.3209839, 
    0.3302307, 0.3489685, 0.3676453, 0.4160767, 0.4150391, 0.4226685, 
    0.4420471, 0.4658203, 0.4675293, 0.4781189, 0.4820557, 0.5101318, 
    0.548584, 0.5873718, 0.6165466, 0.6271667, 0.6358948, 0.6602783, 
    0.6632385, 0.6673279, 0.6802979, 0.6898499, 0.7163696, 0.7171326, 
    0.7325745, 0.7375793, 0.7840576, 0.8283997, 0.8798523, 0.9347229, 
    0.9612732, 0.9845886, 1.01413, 1.016876, 1.004547, 0.957489, 0.916626, 
    0.8948059, 0.8955078, 0.9273376, 0.9701538, 1.029968, 1.055023, 1.1362, 
    1.250366, 1.399231, 1.577026, 1.770447, 1.913757, 2.031158, 2.138153, 
    2.203339, 2.191742, 2.14032, 2.075836, 1.854706, 1.682068, 1.512512, 
    1.373657, 1.206451, 1.073853, 1.02066, 1.02417, 1.00061, 0.9955444,
  1.024323, 1, 0.9891968, 0.9721375, 0.9533997, 0.9277344, 0.9074402, 
    0.8754883, 0.8504028, 0.8233337, 0.803772, 0.7772827, 0.7454834, 
    0.7225952, 0.6968994, 0.6746826, 0.6528931, 0.6340027, 0.630249, 
    0.625061, 0.6237183, 0.5985718, 0.5894775, 0.5992432, 0.5957642, 
    0.5951538, 0.5808105, 0.5649109, 0.5470276, 0.5374451, 0.5411682, 
    0.541626, 0.5527649, 0.571106, 0.591095, 0.6101074, 0.6313477, 0.6433105, 
    0.6572876, 0.6635437, 0.6764526, 0.6808167, 0.693573, 0.6930237, 
    0.7002563, 0.7220154, 0.7429199, 0.7644043, 0.7860107, 0.8008728, 
    0.8041382, 0.7991028, 0.791748, 0.8052368, 0.8035278, 0.8195496, 
    0.8363953, 0.8451233, 0.8695068, 0.8972778, 0.9386292, 0.9881592, 
    1.031616, 1.060822, 1.071808, 1.089325, 1.099091, 1.133392, 1.145721, 
    1.18576, 1.230347, 1.256317, 1.254578, 1.269684, 1.268494, 1.234467, 
    1.209625, 1.194611, 1.187256, 1.185547, 1.183411, 1.183533, 1.150665, 
    1.139008, 1.128021, 1.129883, 1.115387, 1.096497, 1.092712, 1.109314, 
    1.114319, 1.094604, 1.072357, 1.086853, 1.07547, 1.061157,
  2.595551, 2.585526, 2.573166, 2.556625, 2.537155, 2.514694, 2.491394, 
    2.468613, 2.449188, 2.427841, 2.403702, 2.383118, 2.364441, 2.345627, 
    2.326492, 2.308517, 2.290878, 2.274536, 2.258774, 2.243027, 2.227707, 
    2.215668, 2.207474, 2.204605, 2.204086, 2.207993, 2.215668, 2.225433, 
    2.235397, 2.244904, 2.253174, 2.259094, 2.260788, 2.257599, 2.255005, 
    2.244247, 2.235535, 2.227188, 2.220169, 2.212021, 2.204544, 2.195999, 
    2.18898, 2.179672, 2.169647, 2.161041, 2.154266, 2.150375, 2.14093, 
    2.139053, 2.124725, 2.125702, 2.144455, 2.126678, 2.114166, 2.110855, 
    2.118668, 2.107925, 2.12999, 2.157288, 2.1259, 2.204468, 2.199265, 
    2.256683, 2.293015, 2.335144, 2.37532, 2.431427, 2.480972, 2.483521, 
    2.491333, 2.518082, 2.586578, 2.700302, 2.506546, 2.502975, 2.491394, 
    2.679871, 2.543472, 2.510529, 2.507858, 2.513657, 2.520752, 2.527649, 
    2.528183, 2.53775, 2.548431, 2.560211, 2.572708, 2.584167, 2.595169, 
    2.609756, 2.617691, 2.618286, 2.614624, 2.603561,
  2.635727, 2.648422, 2.657135, 2.670547, 2.682602, 2.676819, 2.642944, 
    2.582794, 2.529663, 2.492172, 2.468338, 2.476883, 2.535141, 2.625168, 
    2.730515, 2.822891, 2.871658, 2.855515, 2.763, 2.622452, 2.468475, 
    2.320694, 2.201996, 2.122375, 2.104736, 2.122711, 2.167419, 2.222244, 
    2.269958, 2.305969, 2.323166, 2.314102, 2.277588, 2.233566, 2.195755, 
    2.165085, 2.143402, 2.13501, 2.137955, 2.146927, 2.190292, 2.240051, 
    2.288223, 2.315033, 2.343811, 2.400787, 2.359177, 2.340103, 2.304688, 
    2.285019, 2.22142, 2.100983, 2.03978, 1.90834, 1.996872, 1.68782, 
    1.603714, 1.547791, 1.490753, 1.460938, 1.435547, 1.405655, 1.428787, 
    1.502213, 1.643799, 1.815033, 2.064316, 2.365616, 2.642441, 2.875824, 
    3.068802, 3.1651, 3.1427, 3.111969, 2.992447, 2.916397, 2.84491, 
    2.803589, 2.776291, 2.692245, 2.675003, 2.720184, 2.595764, 2.608139, 
    2.524338, 2.478119, 2.366913, 2.359299, 2.376434, 2.419067, 2.473251, 
    2.529892, 2.562759, 2.593094, 2.611374, 2.622833,
  2.638855, 2.667496, 2.667236, 2.56926, 2.452255, 2.33931, 2.239822, 
    2.267426, 2.32576, 2.389771, 2.484695, 2.548996, 2.58136, 2.549072, 
    2.492889, 2.422562, 2.383911, 2.384552, 2.45253, 2.610077, 2.921921, 
    3.339767, 3.693863, 3.675629, 3.323822, 2.887939, 2.574402, 2.513, 
    2.555466, 2.618866, 2.635605, 2.583176, 2.498352, 2.409164, 2.313263, 
    2.252731, 2.247696, 2.287018, 2.331177, 2.388077, 2.441071, 2.517319, 
    2.608597, 2.813599, 3.229752, 3.551102, 3.78363, 3.81398, 3.686386, 
    3.478043, 3.215027, 2.955734, 2.758087, 2.632294, 2.522644, 2.534058, 
    2.504227, 2.275513, 1.939713, 1.6026, 1.351044, 1.256516, 1.243301, 
    1.328186, 1.361328, 1.386002, 1.564377, 1.866852, 2.169785, 2.450577, 
    2.563919, 2.537888, 2.47467, 2.457169, 2.492508, 2.605133, 2.797653, 
    2.988144, 3.063812, 3.081833, 3.140549, 3.249023, 3.202347, 3.148178, 
    3.008591, 2.9888, 2.88855, 2.669724, 2.549942, 2.43013, 2.373825, 
    2.356064, 2.368881, 2.427078, 2.501862, 2.572632,
  1.920105, 2.112946, 2.235413, 2.284286, 2.24646, 2.175964, 2.127319, 
    2.161819, 2.238266, 2.292816, 2.341644, 2.395157, 2.407074, 2.332535, 
    2.146988, 2.023102, 1.922318, 1.889694, 1.882538, 1.86731, 1.957214, 
    2.057281, 2.149918, 2.167114, 2.100571, 2.01619, 1.915024, 1.958191, 
    2.142685, 2.401474, 2.618469, 2.747177, 2.783569, 2.727859, 2.601028, 
    2.412811, 2.273361, 2.210266, 2.163452, 2.178436, 2.270844, 2.373108, 
    2.449615, 2.48085, 2.619919, 3.165115, 2.007355, 2.216736, 2.382095, 
    2.244202, 2.192383, 2.314896, 2.354874, 2.348251, 2.27774, 2.213684, 
    2.344009, 2.367126, 2.125198, 1.804092, 1.541718, 1.28743, 1.217697, 
    1.209045, 1.294601, 1.427353, 1.66217, 1.791992, 1.923294, 2.088608, 
    2.21315, 2.336014, 2.458267, 2.600845, 2.830536, 3.05957, 3.162628, 
    3.128784, 3.085678, 3.153259, 3.091537, 3.365952, 3.416351, 3.45755, 
    3.540695, 3.627472, 3.731125, 3.681442, 3.673569, 3.109177, 2.743942, 
    2.42598, 2.125717, 1.919662, 1.833725, 1.840286,
  2.368805, 2.338806, 2.333588, 2.301758, 2.239258, 2.227341, 2.186722, 
    2.160217, 2.17897, 2.231308, 2.242432, 2.191589, 2.095825, 1.913971, 
    2.087479, 2.247055, 1.990738, 1.843918, 1.710068, 1.397705, 1.14682, 
    1.480865, 1.690689, 1.816833, 1.978699, 2.181961, 2.112549, 2.155594, 
    2.273163, 2.401154, 2.590271, 2.913071, 3.110275, 3.079086, 2.92804, 
    2.803375, 2.814178, 2.847443, 2.799789, 2.492645, 2.24231, 2.072327, 
    2.014511, 2.138153, 2.441467, 2.992188, 2.309387, 2.6987, 2.678253, 
    2.793289, 2.78685, 2.612564, 2.445435, 2.340363, 2.328064, 2.343033, 
    2.352219, 2.324997, 2.2509, 2.171356, 1.972076, 1.820633, 1.605011, 
    1.485153, 1.428131, 1.341919, 1.350204, 1.312363, 1.507034, 1.687424, 
    1.624283, 1.366028, 1.686401, 2.078583, 2.400467, 2.709183, 3.194672, 
    3.308075, 3.280273, 3.153656, 3.186722, 3.232803, 3.391144, 3.667831, 
    3.873383, 3.953705, 3.978394, 3.942047, 3.888733, 3.649734, 3.181839, 
    3.135803, 2.746552, 2.587357, 2.561066, 2.423752,
  4.110291, 3.704178, 3.731888, 3.406387, 3.22702, 3.067459, 3.105133, 
    3.105728, 3.389908, 3.556519, 3.547928, 3.150848, 2.71666, 2.320251, 
    2.142517, 2.11615, 1.747589, 1.592636, 1.581314, 1.57103, 1.466858, 
    1.41713, 1.242371, 1.180344, 1.213531, 1.332809, 1.488083, 1.591736, 
    1.615692, 1.571472, 1.520905, 1.667252, 1.86673, 2.053635, 2.089584, 
    2.093491, 2.120377, 2.149673, 2.116806, 2.118347, 2.221542, 2.504227, 
    2.95723, 3.397079, 3.138931, 3.423035, 3.527863, 3.3974, 3.299149, 
    3.137497, 2.884674, 2.696732, 2.590942, 2.536514, 2.507141, 2.488068, 
    2.431168, 2.261398, 2.091019, 1.953781, 1.848831, 1.749161, 1.717377, 
    1.636063, 1.658386, 1.67038, 1.686981, 1.761261, 1.853836, 1.983978, 
    2.018036, 2.061401, 2.360748, 2.637161, 2.958069, 3.050064, 3.173889, 
    3.255264, 4.060349, 4.184891, 4.216599, 4.210159, 4.340179, 4.370636, 
    4.346619, 4.383072, 4.43782, 4.376297, 4.389984, 4.38678, 4.236984, 
    4.038086, 3.745392, 3.688675, 3.751572, 3.905533,
  4.381775, 4.394012, 4.316269, 4.121811, 3.848572, 3.681778, 3.638733, 
    3.74707, 3.940094, 4.115356, 4.339127, 4.4888, 4.461975, 4.35527, 
    3.936462, 3.277466, 2.849945, 2.728973, 2.866531, 3.134567, 3.306061, 
    3.223694, 2.929169, 2.521866, 2.134247, 1.801117, 1.818817, 1.707886, 
    1.367386, 1.119003, 1.091339, 1.327148, 1.365158, 2.030594, 2.302933, 
    2.699738, 2.833527, 3.12207, 3.352707, 3.556686, 3.735397, 3.956375, 
    4.202469, 4.509247, 4.651855, 4.481812, 4.042145, 3.419983, 2.746735, 
    2.339905, 2.031158, 1.837555, 1.799011, 1.881897, 1.821472, 1.881958, 
    2.062622, 2.05246, 2.111176, 2.192291, 2.213959, 2.452026, 2.797775, 
    3.202728, 3.782516, 4.462875, 5.105591, 5.933167, 6.649963, 7.352173, 
    7.704773, 8.263885, 8.087143, 7.959824, 7.528107, 6.995575, 6.06781, 
    5.360977, 5.005783, 5.360535, 5.726349, 5.611832, 5.511368, 5.374924, 
    5.154877, 4.955719, 4.856888, 4.839828, 4.836639, 4.701889, 4.512634, 
    4.242188, 3.993881, 3.878845, 3.974869, 4.225388,
  5.007294, 5.316589, 5.363327, 5.443222, 5.389511, 5.146591, 5.057465, 
    5.069916, 5.262619, 5.409744, 5.646271, 5.936905, 6.046616, 6.159698, 
    6.338333, 6.248413, 5.933197, 5.762497, 5.58313, 5.31041, 5.001694, 
    4.649277, 4.265427, 3.854553, 3.599213, 3.148376, 2.857941, 2.454758, 
    2.003769, 1.396149, 0.8649902, 1.216217, 1.4534, 2.239685, 2.308899, 
    2.575287, 3.148956, 3.358459, 3.420502, 3.000061, 3.073029, 3.00589, 
    3.071655, 3.58548, 4.137482, 4.195496, 3.077271, 1.725525, 0.02108765, 
    -0.9257202, -1.240143, -1.361481, -1.292206, -1.315887, -1.177429, 
    -1.126923, -0.8879089, -0.4977417, 0.4694519, 1.34256, 2.399475, 
    2.836395, 3.243225, 3.712158, 3.981812, 3.878571, 3.585266, 3.408112, 
    3.553223, 3.750519, 4.131683, 4.30545, 4.617645, 4.965363, 5.124329, 
    5.029724, 4.810608, 4.691254, 4.699921, 4.695374, 5.05072, 5.536163, 
    6.053558, 6.161102, 5.953156, 5.709869, 5.516922, 5.317169, 5.121017, 
    4.92485, 4.808441, 4.69458, 4.464233, 4.212479, 4.178558, 4.489746,
  5.101685, 5.400299, 5.828552, 5.987793, 6.310211, 6.47171, 6.156494, 
    5.699768, 5.429932, 5.324463, 4.908966, 4.784302, 5.232391, 5.766785, 
    6.372894, 6.99588, 6.961365, 7.370758, 7.694763, 6.67038, 5.728973, 
    5.114105, 4.489899, 4.039368, 3.874664, 3.8927, 3.621033, 3.701202, 
    3.685913, 3.452637, 2.825165, 2.038971, 1.398926, 1.110413, 1.054871, 
    1.207733, 1.463776, 1.573425, 1.631805, 1.781342, 2.040039, 2.435547, 
    2.90094, 3.060425, 2.813812, 2.612457, 2.466248, 1.797943, 0.8056335, 
    0.2864075, 0.07403564, -0.03683472, -0.1463928, -0.3079224, -0.4786682, 
    -0.6708069, -0.6809387, -0.3209839, 0.2051086, 0.7070007, 1.074921, 
    1.255493, 1.429504, 1.640717, 1.779724, 1.908478, 2.138733, 2.268066, 
    2.298523, 2.401306, 2.439941, 2.42392, 2.493958, 2.52301, 2.455719, 
    2.276062, 1.941711, 1.814331, 1.840271, 1.890564, 1.991302, 2.268585, 
    2.781677, 3.524994, 3.779144, 4.429016, 4.851532, 5.262115, 5.39505, 
    5.367371, 5.466736, 5.435211, 5.440216, 5.01535, 4.497833, 4.72406,
  3.460602, 3.524017, 3.405518, 3.285126, 3.191101, 3.10611, 3.09613, 
    2.999725, 2.678955, 2.518738, 2.507019, 2.534607, 2.598053, 2.721527, 
    2.929626, 3.180145, 3.497894, 3.887939, 4.300873, 4.475311, 4.372986, 
    3.827667, 2.980896, 2.519257, 2.278564, 2.296326, 2.380127, 2.415588, 
    2.35965, 2.272888, 2.067474, 1.746765, 1.470093, 1.37854, 1.486816, 
    1.732513, 1.910278, 1.970276, 1.871002, 1.815765, 2.081085, 2.611755, 
    2.990723, 2.831421, 2.35907, 2.171722, 2.140198, 1.974518, 1.52597, 
    1.097473, 0.7958679, 0.5966492, 0.4376831, 0.3260193, 0.2579651, 
    0.2532654, 0.3517151, 0.534668, 0.7653198, 0.9194946, 0.9629822, 
    1.011292, 1.081024, 1.164429, 1.257141, 1.384033, 1.524963, 1.636902, 
    1.70166, 1.766113, 1.819092, 1.864807, 1.847168, 1.746277, 1.54892, 
    1.366791, 1.489288, 2.393799, 2.285522, 1.470886, 1.422028, 1.536102, 
    2.020996, 2.047729, 2.007874, 2.215149, 2.598419, 3.310791, 3.820557, 
    4.019012, 4.014709, 3.777161, 3.705322, 3.482086, 3.182007, 3.209351,
  2.120544, 2.22998, 2.355072, 2.434143, 2.454315, 2.477386, 2.553436, 
    2.638641, 2.654144, 2.665802, 2.748657, 2.813263, 2.78244, 2.71814, 
    2.715973, 2.802124, 3.081024, 3.443329, 3.54834, 3.399902, 3.320923, 
    3.369171, 3.245789, 2.95816, 2.749054, 2.73349, 2.802246, 2.828156, 
    2.763458, 2.580109, 2.288574, 1.936737, 1.710907, 1.70343, 1.839691, 
    1.98114, 1.959686, 1.779083, 1.619507, 1.716125, 2.121857, 2.559326, 
    2.637115, 2.381805, 2.32074, 2.26416, 2.123016, 2.046906, 1.756409, 
    1.325348, 1.102173, 1.045166, 1.031006, 1.033997, 1.003235, 0.9901123, 
    1.016968, 1.147034, 1.302094, 1.343079, 1.308167, 1.306091, 1.290527, 
    1.269165, 1.271271, 1.308746, 1.326141, 1.319824, 1.307465, 1.301849, 
    1.31012, 1.318756, 1.288239, 1.205841, 1.136566, 1.357086, 2.276703, 
    2.453888, 2.040344, 1.817749, 1.548187, 1.487671, 1.991089, 2.011749, 
    1.780304, 1.76825, 1.97049, 2.204254, 2.34729, 2.434021, 2.402832, 
    2.290009, 2.202515, 2.130127, 2.071442, 2.051849,
  2.100281, 2.236359, 2.379333, 2.486115, 2.56311, 2.685944, 2.906158, 
    3.113129, 3.219238, 3.360382, 3.565125, 3.664154, 3.570923, 3.456207, 
    3.328674, 3.157196, 3.160187, 3.443207, 3.625153, 3.808044, 4.258118, 
    4.476257, 4.091248, 3.472351, 3.102783, 2.957306, 2.860565, 2.748322, 
    2.595276, 2.348724, 2.0354, 1.808105, 1.742432, 1.751068, 1.75412, 
    1.681366, 1.506989, 1.306732, 1.193665, 1.334991, 1.993256, 2.550507, 
    2.513062, 2.366364, 2.608826, 2.770203, 2.250549, 2.052185, 1.928406, 
    1.771576, 1.79364, 1.882172, 1.846069, 1.73941, 1.663269, 1.632538, 
    1.591827, 1.597015, 1.679596, 1.699249, 1.675812, 1.595123, 1.455505, 
    1.380249, 1.366119, 1.319183, 1.282196, 1.281921, 1.267853, 1.24826, 
    1.254791, 1.282135, 1.30304, 1.264221, 1.217102, 1.314819, 1.836304, 
    2.05365, 2.065582, 1.809662, 1.609283, 1.563812, 1.759277, 1.659607, 
    1.561462, 1.692993, 1.903687, 2.083038, 2.147827, 2.090607, 1.98996, 
    1.924652, 1.902893, 1.862671, 1.871582, 1.963318,
  2.323853, 2.437592, 2.473999, 2.450409, 2.49588, 2.934937, 3.680237, 
    4.170868, 4.344177, 4.486816, 4.621338, 4.483154, 4.03891, 3.629333, 
    3.358582, 3.161377, 3.089752, 3.150238, 3.332886, 3.527313, 3.587189, 
    3.356598, 2.841827, 2.338318, 2.084534, 1.96402, 1.861511, 1.731232, 
    1.614288, 1.519897, 1.507935, 1.56488, 1.496155, 1.333435, 1.224121, 
    1.21405, 1.225891, 1.292877, 1.496063, 1.686218, 2.255737, 2.758545, 
    2.593781, 2.462402, 2.711212, 2.920197, 2.539429, 2.293854, 2.395294, 
    2.533752, 2.668762, 2.617432, 2.372955, 2.09729, 1.956299, 1.893127, 
    1.737213, 1.635071, 1.686035, 1.72998, 1.693909, 1.622833, 1.529419, 
    1.503632, 1.492798, 1.424225, 1.400604, 1.39267, 1.358368, 1.4151, 
    1.482849, 1.484039, 1.454376, 1.406036, 1.343201, 1.243378, 1.218445, 
    1.438568, 1.693329, 1.761292, 1.690735, 1.694458, 1.816437, 1.960114, 
    2.088043, 2.199066, 2.250641, 2.27652, 2.298859, 2.201477, 2.042084, 
    1.984039, 1.968689, 1.950867, 2.017029, 2.165405,
  2.091919, 2.078888, 2.024841, 2.077637, 2.421967, 3.153595, 3.437927, 
    3.48703, 3.567627, 3.414673, 2.991516, 2.615265, 2.243134, 1.98526, 
    1.849579, 1.841095, 1.902252, 1.977814, 2.023315, 1.949646, 1.756287, 
    1.476593, 1.209076, 1.061584, 0.9942322, 0.9796448, 0.9926147, 1.028351, 
    1.268127, 1.866943, 2.043762, 1.74411, 1.449585, 1.064941, 0.943573, 
    1.406219, 1.621185, 1.64679, 1.772034, 2.037537, 2.237091, 2.799957, 
    3.013062, 2.755493, 2.749664, 2.869873, 2.789032, 2.536041, 2.539154, 
    2.40799, 2.186951, 2.051727, 1.929993, 1.779205, 1.711945, 1.695679, 
    1.633881, 1.613373, 1.716949, 1.764618, 1.75473, 1.773468, 1.734283, 
    1.733185, 1.719299, 1.673218, 1.673889, 1.630768, 1.625427, 1.689941, 
    1.699829, 1.65744, 1.605042, 1.525238, 1.420532, 1.233826, 1.095093, 
    1.390198, 1.865387, 1.76416, 1.677979, 1.891235, 2.331726, 2.648132, 
    2.923004, 2.844238, 2.676178, 2.518127, 2.352234, 2.18454, 2.066986, 
    2.01767, 1.985626, 1.975616, 1.977509, 2.004669,
  1.903534, 1.888885, 1.856354, 1.991058, 2.264435, 2.376709, 2.363129, 
    2.235382, 2.518127, 2.27597, 1.515045, 1.385986, 1.405762, 1.348541, 
    1.246307, 1.234253, 1.267456, 1.226074, 1.094635, 0.8550415, 0.7055664, 
    0.7267456, 0.8103638, 0.9691467, 1.187012, 1.401093, 1.586945, 1.86615, 
    2.350677, 2.391785, 1.722046, 1.615082, 1.614349, 1.563324, 1.612549, 
    1.727234, 1.695953, 2.009399, 2.060455, 2.083801, 2.055695, 2.967163, 
    3.666046, 3.45694, 3.12381, 3.060852, 2.718323, 2.292816, 1.986542, 
    1.504456, 1.225739, 1.216095, 1.255646, 1.35022, 1.496185, 1.603149, 
    1.682404, 1.775299, 1.885315, 1.937164, 1.971985, 2.003998, 1.979218, 
    1.961365, 1.929413, 1.879395, 1.839294, 1.755249, 1.701416, 1.67157, 
    1.59613, 1.555817, 1.451141, 1.328674, 1.270416, 1.042358, 1.037659, 
    1.923096, 2.295288, 2.036682, 2.018982, 2.437134, 2.803284, 2.943604, 
    2.514587, 2.276398, 2.166046, 2.01709, 1.883698, 1.90451, 1.891846, 
    1.87439, 1.805786, 1.726318, 1.738708, 1.820618,
  1.736298, 1.681213, 1.659149, 1.691071, 1.815613, 2.731415, 3.299225, 
    3.418579, 3.303741, 2.226929, 2.009399, 1.963562, 1.880341, 1.731903, 
    1.612335, 1.660522, 1.690002, 1.646179, 1.635651, 1.656403, 1.814209, 
    1.977051, 2.059875, 2.171204, 2.30014, 2.378174, 2.467072, 2.578156, 
    2.452332, 1.912781, 1.648071, 1.701935, 1.641815, 1.862396, 2.023254, 
    2.041199, 2.002899, 2.055176, 2.000763, 2.242798, 2.374176, 2.636108, 
    2.519012, 2.667542, 2.697357, 2.602112, 2.160034, 1.629974, 1.342468, 
    1.163452, 1.232391, 1.424713, 1.610962, 1.729462, 1.810364, 1.845856, 
    1.870789, 1.943909, 1.981598, 2.029541, 2.051666, 2.016693, 1.963501, 
    1.942047, 1.912262, 1.83786, 1.721924, 1.557343, 1.437286, 1.356232, 
    1.273254, 1.225891, 1.144318, 1.114227, 1.102051, 0.9201965, 1.209473, 
    3.239807, 3.690002, 2.486633, 2.106018, 2.794617, 2.977753, 2.541473, 
    2.231903, 1.935944, 1.815247, 1.80365, 1.926544, 1.950623, 1.896057, 
    1.860931, 1.834015, 1.791779, 1.791046, 1.776337,
  1.549133, 1.525482, 1.67746, 1.938599, 2.29364, 3.218079, 4.047821, 
    4.428009, 3.747742, 2.373077, 2.158875, 2.241638, 2.252716, 2.155975, 
    2.257477, 2.401672, 2.472717, 2.484192, 2.497192, 2.519684, 2.525848, 
    2.518036, 2.495819, 2.45639, 2.425079, 2.33316, 2.230682, 2.05481, 
    1.900269, 1.779419, 1.768555, 2.266815, 2.018311, 2.03891, 2.060913, 
    2.064667, 2.079651, 2.088379, 1.8396, 2.000854, 2.249847, 1.991089, 
    1.70343, 1.726746, 1.824677, 1.796021, 1.755615, 1.778717, 1.79892, 
    1.8927, 1.933472, 1.908905, 1.895111, 1.865356, 1.845032, 1.792328, 
    1.759979, 1.786804, 1.81485, 1.859894, 1.83667, 1.773315, 1.738342, 
    1.72525, 1.685089, 1.582642, 1.449127, 1.272827, 1.157227, 1.080536, 
    1.010498, 1.021332, 1.029144, 0.9564819, 0.8557739, 0.9222412, 1.68161, 
    3.937408, 4.780426, 3.050446, 2.702026, 3.442352, 3.577179, 3.231262, 
    2.357788, 1.96814, 1.875549, 2.004486, 1.997009, 1.927673, 1.91275, 
    1.85321, 1.792664, 1.748779, 1.682007, 1.625641,
  1.624634, 1.795105, 2.053711, 2.450439, 3.609924, 3.676392, 4.649506, 
    5.337402, 4.990997, 4.235046, 2.306793, 2.398865, 3.65683, 2.288391, 
    2.320404, 2.489746, 2.438629, 2.432281, 2.37146, 2.328278, 2.247772, 
    2.176453, 2.124634, 2.08786, 2.039459, 2.009552, 1.987823, 1.933167, 
    1.907867, 1.96756, 2.028473, 2.993011, 2.711853, 2.30069, 2.268829, 
    2.038574, 1.81546, 1.78949, 2.068909, 2.106415, 2.103119, 1.85611, 
    1.942871, 2.066956, 2.141113, 2.112061, 2.076599, 2.091949, 2.042236, 
    1.970551, 1.888702, 1.806427, 1.77829, 1.712402, 1.672974, 1.672485, 
    1.657074, 1.688782, 1.732635, 1.778198, 1.776001, 1.776276, 1.740784, 
    1.690277, 1.585083, 1.399292, 1.257507, 1.139038, 1.048737, 0.9929504, 
    0.9747925, 0.97995, 0.9462585, 0.8565369, 0.9987488, 1.37204, 2.300385, 
    4.42157, 5.03479, 3.6185, 4.072968, 4.636719, 4.694275, 3.436432, 
    3.416779, 2.173462, 1.852844, 1.879395, 1.886688, 1.787079, 1.759064, 
    1.698914, 1.597748, 1.538879, 1.477081, 1.535614,
  2.001587, 2.221161, 2.38092, 2.600311, 4.429047, 4.794464, 5.05072, 
    5.177673, 4.846161, 4.371552, 2.386505, 2.496582, 3.729462, 2.927765, 
    2.164612, 2.256042, 2.209656, 2.188263, 2.17215, 2.147644, 2.108826, 
    2.080322, 2.064484, 2.056152, 2.093719, 2.110046, 2.108826, 2.056488, 
    2.04657, 2.143127, 2.204712, 2.128357, 2.515045, 2.631287, 2.417145, 
    2.142456, 1.90921, 2.260925, 2.891937, 2.59317, 2.080414, 2.163055, 
    2.32309, 2.394836, 2.333374, 2.225433, 2.1203, 2.032257, 1.926117, 
    1.813629, 1.775879, 1.751923, 1.710846, 1.668579, 1.7258, 1.78949, 
    1.816528, 1.875549, 1.906403, 1.945801, 1.979279, 1.995209, 1.916382, 
    1.820282, 1.681671, 1.499359, 1.384552, 1.275085, 1.190735, 1.136169, 
    1.078094, 1.042816, 1.041016, 1.210419, 1.45163, 1.616425, 2.543579, 
    4.830658, 4.397614, 3.772949, 4.826416, 5.832672, 4.611359, 4.112091, 
    3.948792, 3.45163, 1.93576, 1.888428, 1.889435, 1.818848, 1.746582, 
    1.673096, 1.628601, 1.643005, 1.724792, 1.871674,
  2.437469, 2.444366, 2.482452, 2.570404, 4.627197, 4.844574, 4.964111, 
    4.927795, 4.739319, 4.512238, 3.74646, 2.558502, 3.791931, 3.186188, 
    2.115601, 2.133362, 2.143646, 2.14801, 2.166382, 2.186035, 2.190643, 
    2.214691, 2.231018, 2.26886, 2.283356, 2.272949, 2.233887, 2.207245, 
    2.279724, 2.36853, 2.401855, 2.336578, 2.451141, 3.85083, 3.390503, 
    3.084564, 2.906891, 2.562012, 3.063324, 2.348816, 2.424774, 2.643188, 
    2.625641, 2.597015, 2.442871, 2.262054, 2.147156, 2.031158, 1.955444, 
    1.894836, 1.874756, 1.853546, 1.856781, 1.914703, 2.006012, 2.082214, 
    2.156158, 2.21344, 2.212646, 2.243011, 2.251617, 2.251465, 2.195679, 
    2.07724, 2.015198, 1.961304, 1.864868, 1.774445, 1.714447, 1.654144, 
    1.595642, 1.648193, 1.807068, 1.894257, 1.899689, 2.141357, 4.233246, 
    4.821136, 3.457001, 4.104095, 4.86377, 4.840576, 4.374786, 3.758118, 
    4.117554, 2.957886, 1.97699, 2.0177, 1.989349, 1.979614, 1.998413, 
    2.049194, 2.101135, 2.148193, 2.244293, 2.345398,
  2.613495, 2.554016, 2.595673, 2.600372, 4.473999, 4.987488, 4.506042, 
    4.587372, 4.497009, 4.113373, 3.899658, 2.378235, 2.196198, 2.093445, 
    2.058167, 2.136566, 2.176483, 2.231598, 2.271576, 2.338837, 2.354004, 
    2.380219, 2.376404, 2.392212, 2.326202, 2.310852, 2.345947, 2.358826, 
    2.438629, 2.558167, 2.651917, 2.703735, 2.7258, 2.793274, 2.809479, 
    3.771332, 3.478271, 2.728149, 3.251984, 2.465332, 2.61554, 2.672882, 
    2.562592, 2.480286, 2.350494, 2.217957, 2.114502, 2.044495, 2.03363, 
    2.039093, 2.043152, 2.05835, 2.116364, 2.188965, 2.24585, 2.32132, 
    2.377625, 2.447571, 2.452637, 2.470032, 2.47757, 2.454987, 2.406097, 
    2.359467, 2.335205, 2.255768, 2.181213, 2.177124, 2.146057, 2.130096, 
    2.184662, 2.245148, 2.251862, 2.111389, 2.219757, 3.511627, 4.122986, 
    3.600403, 3.576508, 5.106354, 4.493652, 4.503082, 4.504059, 3.645874, 
    3.64032, 3.027405, 2.051025, 2.147491, 2.151031, 2.238464, 2.276642, 
    2.330566, 2.383423, 2.47113, 2.545593, 2.628723,
  2.597443, 2.665741, 2.691559, 2.544678, 3.93396, 4.392151, 3.923187, 
    3.865143, 3.983459, 3.91333, 3.560974, 2.308777, 2.134735, 2.120392, 
    2.168213, 2.254272, 2.284668, 2.361145, 2.37854, 2.398621, 2.398193, 
    2.415771, 2.38443, 2.373718, 2.371582, 2.400269, 2.410889, 2.406738, 
    2.425415, 2.544312, 2.65213, 2.673218, 2.658569, 2.686615, 2.60791, 
    2.598663, 2.527191, 2.496582, 2.654205, 2.485626, 2.554413, 2.485138, 
    2.4422, 2.363586, 2.260986, 2.192566, 2.093201, 2.067963, 2.07016, 
    2.093262, 2.118988, 2.151672, 2.167938, 2.205688, 2.237457, 2.310242, 
    2.364471, 2.426941, 2.476593, 2.501404, 2.511017, 2.514618, 2.491241, 
    2.486023, 2.435333, 2.408478, 2.400818, 2.38858, 2.387482, 2.394897, 
    2.404541, 2.343567, 2.3255, 2.289825, 2.349304, 3.042877, 3.584412, 
    4.652344, 4.241455, 4.334381, 4.202576, 4.256744, 4.402191, 4.039948, 
    3.439819, 3.149658, 2.719177, 2.239685, 2.286682, 2.363525, 2.396912, 
    2.446716, 2.478271, 2.589355, 2.602203, 2.64566,
  2.73233, 2.939819, 2.893585, 2.926605, 4.100037, 4.045868, 3.583618, 
    3.473999, 3.321259, 2.727783, 2.76944, 2.264374, 2.183746, 2.242096, 
    2.300354, 2.359497, 2.448639, 2.49939, 2.466431, 2.432922, 2.403503, 
    2.395355, 2.374329, 2.397491, 2.396515, 2.478149, 2.442017, 2.393005, 
    2.654968, 2.496002, 2.472015, 2.537262, 2.537201, 2.587402, 2.653534, 
    2.440002, 2.288574, 2.561707, 2.914612, 2.88501, 2.563049, 2.320221, 
    2.249573, 2.187653, 2.099365, 2.053162, 1.982269, 1.939026, 1.947083, 
    2.004791, 2.080505, 2.203674, 2.302612, 2.389069, 2.462463, 2.507324, 
    2.557068, 2.561035, 2.541656, 2.544434, 2.534271, 2.531494, 2.510254, 
    2.476471, 2.483887, 2.494293, 2.454071, 2.445251, 2.432709, 2.396118, 
    2.360016, 2.351898, 2.382385, 2.486877, 2.438965, 3.231995, 4.104919, 
    3.878906, 3.20578, 3.794678, 4.142517, 4.283203, 4.281219, 4.4841, 
    4.145416, 3.360626, 3.224365, 2.332642, 2.397034, 2.490326, 2.544312, 
    2.624115, 2.65921, 2.69281, 2.680817, 2.693909,
  2.918335, 3.016632, 2.963715, 3.549713, 4.019958, 3.07666, 2.860382, 
    3.132477, 3.347656, 2.343689, 2.587036, 3.39093, 2.237091, 2.279785, 
    2.442505, 2.462006, 2.559906, 2.541382, 2.4245, 2.32489, 2.307831, 
    2.316833, 2.349243, 2.396576, 2.39859, 2.449585, 2.43396, 2.65274, 
    2.695465, 2.481628, 2.54541, 2.734222, 2.914093, 2.457397, 2.594482, 
    2.617035, 2.54483, 2.876617, 3.124512, 2.557251, 2.447693, 2.252563, 
    2.134796, 2.087585, 2.015656, 1.984924, 1.956757, 1.977112, 2.045929, 
    2.222626, 2.451477, 2.697296, 2.816681, 2.83725, 2.796204, 2.721832, 
    2.640472, 2.581421, 2.537598, 2.493652, 2.469574, 2.476868, 2.502808, 
    2.511292, 2.546844, 2.522095, 2.52594, 2.559204, 2.494293, 2.476288, 
    2.408813, 2.376801, 2.336304, 2.319366, 2.208038, 3.094757, 3.497681, 
    3.240601, 2.976257, 3.288025, 3.443329, 4.414734, 4.754944, 4.289307, 
    3.623962, 2.475616, 2.372833, 2.354645, 2.475922, 2.632843, 2.714355, 
    2.762726, 2.768829, 2.794647, 2.812683, 2.813965,
  2.705048, 2.797241, 2.671387, 2.885071, 2.812744, 2.666718, 2.794312, 
    2.953339, 3.193512, 3.104645, 3.049591, 4.046356, 3.388428, 2.310913, 
    2.505219, 2.564087, 2.609406, 2.501404, 2.297668, 2.163025, 2.147369, 
    2.171112, 2.20874, 2.267426, 2.306549, 2.299622, 2.353424, 2.587677, 
    2.484314, 2.382751, 2.551208, 2.389618, 2.555054, 2.240479, 2.162262, 
    2.032898, 1.915192, 2.038116, 2.283264, 2.436829, 2.331146, 2.192047, 
    2.089508, 2.070068, 2.00351, 2.030609, 2.095978, 2.126526, 2.240417, 
    2.407562, 2.60791, 2.824463, 2.953827, 3.022247, 2.978882, 2.916504, 
    2.797791, 2.715088, 2.658691, 2.585571, 2.561035, 2.543335, 2.536804, 
    2.557648, 2.52951, 2.507904, 2.498993, 2.459351, 2.394684, 2.330444, 
    2.176331, 2.081482, 1.985718, 1.884735, 1.817017, 2.588379, 3.049103, 
    3.104584, 2.707642, 2.788422, 3.372101, 4.295441, 4.334686, 2.575531, 
    2.484589, 2.485504, 2.406464, 2.367401, 2.310486, 2.369507, 2.49826, 
    2.563416, 2.575684, 2.559021, 2.564545, 2.565002,
  2.80368, 2.695557, 2.837006, 2.767151, 2.676819, 2.847748, 3.093994, 
    2.994568, 3.01297, 3.258698, 3.389526, 4.407623, 3.765381, 2.460968, 
    2.408447, 2.530579, 2.626251, 2.672913, 2.524994, 2.400055, 2.229462, 
    2.087341, 2.08905, 2.239288, 2.427582, 2.302612, 2.788177, 2.437714, 
    2.418518, 2.332306, 2.356323, 2.438782, 1.995209, 2.259491, 2.238831, 
    2.159119, 2.173615, 2.167877, 2.242859, 2.269135, 2.220917, 2.154327, 
    2.098999, 2.043915, 2.006805, 2.031036, 2.085449, 2.008362, 2.02301, 
    2.027313, 2.044373, 2.095276, 2.119995, 2.200623, 2.242279, 2.284271, 
    2.280579, 2.323547, 2.346802, 2.373688, 2.421051, 2.44046, 2.427094, 
    2.455109, 2.394043, 2.37973, 2.251068, 2.263123, 2.249237, 2.088318, 
    2.042084, 1.919434, 1.792999, 1.881866, 2.034607, 2.746979, 2.707764, 
    2.80127, 3.152496, 3.258514, 4.074036, 4.069672, 2.707886, 2.289948, 
    2.480408, 2.555878, 2.537659, 2.406799, 2.297089, 2.287262, 2.30368, 
    2.295288, 2.271057, 2.313507, 2.718597, 2.767029,
  2.861572, 2.835205, 2.962646, 2.877228, 2.677521, 2.812988, 2.905304, 
    2.89917, 3.033356, 3.316071, 3.567566, 3.984619, 3.908264, 2.982758, 
    2.594818, 2.631561, 2.473083, 2.479858, 2.485077, 2.434937, 2.403656, 
    2.410919, 2.251526, 2.115204, 2.240204, 2.403015, 2.453918, 2.596832, 
    2.596924, 2.465393, 2.41571, 2.430206, 2.306458, 2.627441, 2.328552, 
    2.247284, 2.263428, 2.237549, 2.216339, 2.149933, 2.149567, 2.151611, 
    2.109192, 2.111176, 2.165527, 2.146393, 2.176086, 2.156006, 2.13028, 
    2.156219, 2.158905, 2.147888, 2.132721, 2.131714, 2.133362, 2.121063, 
    2.101593, 2.123657, 2.112946, 2.153107, 2.133881, 2.245941, 2.328918, 
    2.354553, 2.37677, 2.426788, 2.461304, 2.606537, 2.616516, 2.583557, 
    2.463959, 2.230103, 2.389557, 2.263062, 2.669098, 2.772217, 2.626678, 
    2.983612, 4.407379, 3.539703, 2.369629, 2.351685, 2.350739, 2.36618, 
    2.356873, 2.362732, 2.400177, 2.37027, 2.376526, 2.408234, 2.453491, 
    2.402954, 2.369232, 2.734985, 2.853668, 2.819031,
  2.81131, 2.707855, 2.593048, 2.577423, 2.626129, 3.095337, 3.408508, 
    3.309479, 3.136841, 3.326324, 4.807404, 4.921539, 4.454498, 3.784698, 
    2.599274, 2.581757, 2.59845, 2.466522, 2.423523, 2.381042, 2.657013, 
    2.447357, 2.288361, 2.263519, 2.333221, 2.457672, 2.522583, 2.739655, 
    2.590393, 2.427887, 2.518005, 2.557068, 2.547272, 2.426666, 2.277405, 
    2.25705, 2.233795, 2.20697, 2.191772, 2.112, 2.107941, 2.099762, 
    2.098602, 2.109863, 2.20575, 2.198669, 2.155701, 2.175659, 2.156738, 
    2.180908, 2.184784, 2.177826, 2.232971, 2.282593, 2.282471, 2.288055, 
    2.302826, 2.328491, 2.375824, 2.431732, 2.406097, 2.455048, 2.419189, 
    2.444183, 2.504547, 2.569458, 2.760071, 2.939087, 2.867645, 2.782013, 
    2.585571, 2.706055, 5.314148, 4.416351, 1.990448, 2.123016, 2.281403, 
    2.261475, 2.292603, 2.326324, 2.255829, 2.219635, 2.168243, 2.149323, 
    2.131226, 2.199127, 2.198029, 2.269501, 2.310516, 2.453796, 2.511108, 
    2.324097, 3.146759, 3.264496, 2.914093, 2.689423,
  2.80603, 3.336395, 3.4422, 3.516144, 3.468689, 3.536224, 3.499146, 
    3.872711, 4.031128, 4.309631, 4.759766, 4.473053, 4.676544, 4.452362, 
    2.944916, 2.343262, 2.598419, 2.469055, 2.438446, 2.360046, 2.555237, 
    2.558807, 2.462158, 2.35321, 2.313782, 2.381409, 2.634888, 2.764618, 
    2.338531, 2.30191, 2.290924, 2.577301, 2.647583, 2.257416, 2.161407, 
    2.249695, 2.177673, 2.161713, 2.156708, 2.054749, 2.030823, 2.063751, 
    2.102051, 2.125854, 2.160004, 2.191071, 2.169037, 2.136871, 2.14502, 
    2.164246, 2.187012, 2.217529, 2.271393, 2.308563, 2.287811, 2.31366, 
    2.30542, 2.331085, 2.417206, 2.44632, 2.498077, 2.533936, 2.450836, 
    2.302368, 2.196442, 2.288361, 2.500763, 2.694336, 2.722656, 2.735107, 
    3.430054, 5.48999, 5.201538, 2.055817, 2.119446, 2.264069, 2.188629, 
    2.165192, 2.111938, 2.145721, 2.139008, 2.07608, 2.048462, 2.085968, 
    2.06189, 2.041687, 2.020935, 2.081207, 2.110504, 2.305481, 2.314148, 
    2.202332, 4.593414, 4.853699, 3.255188, 2.751404,
  3.971832, 3.803192, 3.893219, 3.933136, 3.977142, 3.77832, 3.896881, 
    3.918365, 3.949432, 3.527283, 2.591125, 3.86615, 4.8125, 4.367584, 
    4.189056, 2.707611, 2.30661, 2.399506, 2.478241, 2.306, 2.455963, 
    2.669495, 2.640533, 2.563507, 2.365509, 2.611542, 2.570801, 2.662537, 
    2.763062, 2.683838, 2.195282, 2.380096, 2.523193, 2.336975, 2.254089, 
    2.243896, 2.241974, 2.230408, 2.154633, 2.059998, 2.067719, 2.133118, 
    2.094818, 2.092468, 2.087524, 2.096313, 2.115387, 2.152466, 2.178619, 
    2.180695, 2.183868, 2.220154, 2.245148, 2.271912, 2.233429, 2.201843, 
    2.167938, 2.161316, 2.194763, 2.200867, 2.232727, 2.253479, 2.158051, 
    1.952057, 1.666229, 1.401001, 1.724396, 2.442902, 2.801514, 3.309387, 
    4.964508, 5.565033, 4.033264, 2.158386, 2.300659, 2.21994, 2.114105, 
    2.093323, 2.089935, 2.080963, 2.041107, 2.062469, 2.059204, 2.036743, 
    2.00296, 2.000488, 1.960266, 1.947876, 1.892487, 1.948273, 2.012451, 
    2.402252, 4.918304, 5.532623, 4.482819, 4.05838,
  4.348511, 4.535736, 4.10495, 3.89859, 3.749542, 3.49234, 3.685669, 
    3.797974, 4.120728, 4.136658, 2.695496, 4.395233, 4.996033, 4.237152, 
    4.195007, 3.609924, 2.277405, 2.226959, 1.480865, 1.001343, 1.496521, 
    1.908081, 2.335175, 2.54834, 2.649963, 2.657013, 2.653137, 2.587189, 
    2.443909, 2.584656, 2.691895, 2.847229, 2.450989, 2.369843, 2.364197, 
    2.375122, 2.330475, 2.219055, 2.187469, 2.153473, 2.169373, 2.173798, 
    2.135651, 2.103363, 2.031982, 2.044678, 2.078674, 2.083557, 2.097229, 
    2.106537, 2.144775, 2.128937, 2.081146, 2.021393, 2.026337, 2.048096, 
    2.039429, 1.997742, 1.989624, 2.018707, 2.025024, 2.044067, 2.036743, 
    1.865845, 1.530029, 1.094818, 1.733704, 4.672333, 3.693939, 3.430695, 
    3.668365, 2.181213, 1.900146, 2.19339, 2.235199, 2.054932, 2.077271, 
    2.09494, 2.18869, 2.170715, 2.142548, 2.177826, 2.151398, 2.160004, 
    2.128113, 2.087006, 2.033234, 1.991302, 1.955444, 1.898407, 1.798859, 
    2.245026, 3.930939, 5.067261, 4.958771, 4.431702,
  4.557739, 4.241272, 4.011261, 3.89505, 3.812958, 3.482086, 3.788452, 
    3.897705, 3.930664, 4.197662, 4.500641, 4.799591, 4.919983, 4.650208, 
    4.853119, 4.540436, 4.235352, 3.871674, 2.431396, 0.7085266, 1.085114, 
    2.101715, 2.747009, 2.890808, 2.810272, 2.816193, 2.635651, 2.239227, 
    2.141418, 2.626007, 2.927551, 3.033875, 2.883881, 2.490601, 2.405334, 
    2.508636, 2.473816, 2.383362, 2.36618, 2.324768, 2.254089, 2.191742, 
    2.212341, 2.175354, 2.09613, 2.090149, 2.048645, 2.00882, 1.949829, 
    1.938354, 2.023529, 2.092621, 2.081909, 2.022827, 2.000885, 1.978485, 
    1.939301, 1.977509, 1.919006, 1.929352, 1.912903, 1.932251, 1.945923, 
    1.676208, 1.432648, 1.689789, 4.21347, 5.284698, 3.589294, 2.789063, 
    2.398895, 2.261353, 2.370605, 2.517395, 2.991516, 2.0354, 2.012512, 
    2.181793, 2.310059, 2.234009, 2.192932, 2.212341, 2.184326, 2.200043, 
    2.157471, 2.155823, 2.153564, 2.089722, 2.052887, 1.958954, 1.82132, 
    1.765717, 2.180389, 3.888733, 5.175842, 4.769318,
  5.666412, 5.484833, 5.041412, 4.318298, 3.639191, 2.634277, 3.679535, 
    3.613617, 2.686615, 3.589752, 4.769531, 4.766479, 4.543701, 4.857086, 
    4.805054, 5.277802, 4.923767, 4.304169, 3.483307, 2.381653, 2.293335, 
    2.599457, 3.190002, 2.797485, 2.908295, 2.701935, 2.444122, 2.065857, 
    2.301636, 2.508698, 2.618195, 2.814941, 2.845215, 2.378021, 2.288055, 
    2.420807, 2.485535, 2.453796, 2.397308, 2.393646, 2.434937, 2.321381, 
    2.256348, 2.249146, 2.255035, 2.295471, 2.274109, 2.211121, 2.130707, 
    2.084381, 2.086884, 2.085846, 2.138702, 2.171661, 2.191101, 2.145355, 
    2.070435, 2.033173, 1.954529, 1.953278, 1.940521, 1.911407, 1.811066, 
    1.61438, 1.811493, 3.360199, 4.452271, 4.110138, 2.808868, 2.451416, 
    2.003723, 2.458405, 3.279999, 3.531372, 3.396088, 2.22226, 1.944061, 
    2.024384, 2.131989, 2.221893, 2.32843, 2.282257, 2.141754, 2.072815, 
    2.069824, 2.095398, 2.115906, 2.154602, 2.150665, 2.088562, 2.004395, 
    1.869171, 1.751221, 2.238007, 4.049744, 5.263153,
  6.169067, 6.353455, 5.901245, 3.101532, 2.459137, 2.423157, 2.687988, 
    2.90506, 3.012787, 3.213593, 4.425903, 4.544281, 4.456818, 4.382629, 
    4.71405, 5.242188, 5.027924, 4.756409, 4.462067, 4.549469, 3.908752, 
    4.061676, 3.730957, 3.123474, 3.023132, 2.731171, 2.440796, 2.400055, 
    2.585205, 2.635559, 2.438812, 2.462799, 2.47522, 2.271698, 2.347504, 
    2.586609, 2.598267, 2.609131, 2.377686, 2.369537, 2.510986, 2.44519, 
    2.336029, 2.33194, 2.366638, 2.384338, 2.416412, 2.395081, 2.348022, 
    2.334656, 2.338318, 2.308563, 2.276123, 2.254211, 2.33075, 2.403351, 
    2.317352, 2.24353, 2.132324, 2.044617, 2.013214, 1.864197, 1.879181, 
    2.137146, 3.232788, 4.162262, 4.481842, 4.054962, 3.685638, 2.734497, 
    2.128174, 2.70755, 3.547668, 3.224976, 2.846375, 2.637146, 2.324768, 
    2.166809, 2.050995, 2.161163, 2.149323, 2.136688, 2.182861, 2.090851, 
    1.928864, 1.672821, 1.660431, 1.954193, 2.182007, 2.223236, 2.12973, 
    2.009033, 1.759735, 1.792542, 2.535645, 4.975128,
  4.811035, 2.803925, 2.843658, 2.84314, 2.831604, 3.25061, 5.145325, 
    4.933411, 5.287964, 4.988251, 4.386505, 4.406616, 4.227844, 3.721466, 
    2.691071, 4.18042, 4.655548, 4.635071, 4.633484, 4.835205, 4.925873, 
    4.62085, 4.578186, 4.4505, 4.294373, 4.181366, 3.934418, 3.771454, 
    3.523987, 3.27002, 2.973053, 2.657166, 2.473206, 2.441895, 2.473846, 
    2.752502, 2.689178, 2.637573, 2.470032, 2.518829, 2.747955, 2.895813, 
    2.932007, 2.866211, 2.806061, 2.725403, 2.612518, 2.517487, 2.426483, 
    2.406708, 2.409515, 2.448181, 2.44635, 2.34967, 2.349213, 2.332947, 
    2.276184, 2.295593, 2.219391, 2.103729, 2.048889, 1.877045, 2.266754, 
    3.649719, 4.452576, 4.309662, 4.184479, 3.916779, 3.49704, 3.09079, 
    2.062805, 2.389374, 2.976257, 2.979706, 2.939667, 3.093018, 3.023621, 
    2.889404, 2.632599, 2.409546, 2.270935, 2.463501, 2.533112, 2.253143, 
    1.873322, 1.216125, 0.7588806, 1.037018, 1.549896, 1.947968, 2.129791, 
    1.972137, 1.836792, 2.320221, 4.276093, 5.513611,
  4.230286, 2.711578, 3.135651, 4.287598, 3.195709, 5.168945, 5.240631, 
    4.420593, 3.988892, 3.778809, 3.708618, 4.020233, 3.466309, 2.446838, 
    2.959259, 3.478302, 3.820313, 3.790894, 4.118744, 4.65799, 5.001892, 
    5.121033, 5.181702, 4.909149, 4.903656, 5.033295, 4.722137, 4.716736, 
    4.70462, 4.096497, 3.20993, 2.988342, 2.807953, 2.680023, 2.614471, 
    2.580994, 2.51239, 2.547028, 2.886627, 3.239685, 3.245972, 3.277435, 
    3.156403, 2.976074, 2.862579, 2.71579, 2.543213, 2.397797, 2.289948, 
    2.231873, 2.264862, 2.319122, 2.294647, 2.261536, 2.262115, 2.272552, 
    2.296326, 2.26474, 2.146118, 2.182465, 2.177368, 1.934998, 2.353485, 
    4.278473, 4.58905, 4.146362, 3.12793, 3.470306, 3.170319, 2.664948, 
    2.408356, 2.680023, 2.872437, 2.985504, 3.440125, 3.676147, 3.729065, 
    3.703003, 3.523651, 3.217529, 2.79541, 2.618439, 2.474762, 2.105438, 
    1.824463, 1.336761, 0.7746887, 0.7262878, 0.9660034, 1.289795, 1.758545, 
    1.857208, 1.739441, 2.259644, 4.339233, 4.705688,
  3.564423, 3.752197, 3.670135, 3.453278, 2.887909, 2.705902, 2.713837, 
    2.828888, 3.253113, 3.292236, 3.214203, 2.918518, 2.734985, 2.687866, 
    2.436035, 2.92868, 3.122284, 3.306915, 3.915985, 4.318909, 4.481201, 
    4.781677, 5.202789, 5.029846, 4.808197, 4.857697, 4.501617, 4.205872, 
    3.870209, 3.723389, 3.301971, 2.813904, 2.92926, 2.992889, 2.861847, 
    2.914795, 2.917023, 2.618713, 2.798248, 2.819519, 2.548859, 2.634125, 
    2.595093, 2.543457, 2.507904, 2.437531, 2.30246, 2.193909, 2.179535, 
    2.194702, 2.192657, 2.186096, 2.12149, 2.105194, 2.111938, 2.098145, 
    2.117249, 2.11911, 2.09964, 2.187378, 2.194183, 2.022217, 2.346893, 
    3.96582, 4.245605, 3.907318, 3.319427, 3.549652, 3.126434, 3.007446, 
    2.784302, 2.741425, 3.100739, 3.318176, 3.494476, 3.518677, 3.567627, 
    3.587799, 3.638794, 3.587677, 3.164551, 2.610443, 1.827759, 1.576599, 
    1.574646, 1.47998, 1.05661, 0.7655334, 0.6500549, 0.6164246, 1.069244, 
    1.640137, 1.788574, 1.81427, 2.280121, 3.663177,
  2.676147, 2.850281, 2.808014, 2.533844, 1.801666, 1.831879, 1.696106, 
    2.03952, 2.036133, 2.215759, 2.224945, 2.322296, 2.37262, 2.201599, 
    2.028259, 2.344238, 2.749969, 3.036163, 3.441132, 3.927185, 4.180573, 
    4.449249, 4.66626, 4.483093, 4.389679, 4.066956, 3.686157, 3.436157, 
    3.309143, 3.029938, 2.985962, 2.88028, 2.883484, 2.772278, 2.705231, 
    2.922821, 2.991821, 2.780426, 2.11319, 2.42627, 2.775604, 2.835968, 
    2.698517, 2.536743, 2.526978, 2.522186, 2.480591, 2.407562, 2.35321, 
    2.300751, 2.280945, 2.265015, 2.29364, 2.326996, 2.328156, 2.266296, 
    2.202911, 2.19754, 2.161377, 2.110962, 2.076141, 2.188507, 3.172241, 
    3.56369, 3.55246, 3.516174, 3.506622, 3.572998, 3.531433, 3.631256, 
    3.402405, 3.227386, 3.179199, 3.295197, 3.310638, 3.36618, 3.340332, 
    3.127625, 3.064758, 3.164276, 3.071106, 2.894684, 2.077026, 2.028351, 
    1.805878, 1.38208, 0.7254333, 0.09854126, -0.1687622, -0.04782104, 
    0.4468689, 1.084595, 1.522034, 1.637268, 1.795532, 2.059631,
  2.235321, 1.96521, 2.173859, 2.022217, 1.993591, 1.951782, 1.724274, 
    1.18103, 0.9786682, 1.02951, 1.146271, 1.567078, 1.922668, 1.981171, 
    1.88092, 2.061432, 2.593597, 2.936737, 3.417847, 3.800537, 4.142578, 
    4.377472, 4.21106, 4.04306, 3.994446, 3.808746, 3.486176, 3.515717, 
    3.531738, 3.520416, 3.46228, 3.326904, 3.179932, 3.020721, 3.120544, 
    3.324066, 3.322418, 3.143188, 2.118134, 2.33551, 2.860657, 3.121002, 
    3.263763, 2.572021, 2.523712, 2.54541, 2.524048, 2.467224, 2.425476, 
    2.425568, 2.459808, 2.534149, 2.629791, 2.706085, 2.670807, 2.515991, 
    2.374115, 2.313965, 2.212982, 2.131073, 2.09259, 2.703491, 3.019775, 
    3.16214, 3.150818, 3.071259, 3.146851, 3.214172, 3.147827, 3.201263, 
    3.156097, 2.891357, 2.817871, 2.798859, 3.086243, 3.765686, 2.613312, 
    2.402557, 2.461365, 2.617554, 2.467102, 1.989166, 1.661255, 1.340912, 
    1.093079, 1.074188, 0.7827759, 0.1031189, -0.3944397, -0.2924805, 
    0.2831116, 0.8978271, 1.305786, 1.5354, 1.81723, 2.119263,
  1.390137, 1.571991, 1.38797, 1.983368, 2.17453, 2.34079, 2.003204, 
    1.749969, 1.768799, 1.72699, 1.367615, 1.155365, 1.250275, 1.393463, 
    1.729126, 1.923981, 2.307373, 2.76001, 3.338379, 3.660065, 3.753632, 
    3.897797, 3.90094, 4.107239, 4.316101, 3.959595, 3.883881, 3.69931, 
    3.727386, 3.772125, 3.795349, 3.610901, 3.47525, 3.451965, 3.486633, 
    3.749695, 3.704468, 3.563263, 2.188629, 2.150238, 2.215118, 2.188904, 
    3.067596, 3.049896, 2.186768, 2.526611, 2.728546, 2.83374, 2.948181, 
    3.100433, 3.232605, 3.225037, 3.158752, 3.107147, 3.045776, 2.538116, 
    2.38266, 2.344543, 2.298279, 2.16098, 2.614044, 2.819122, 3.007751, 
    2.892883, 2.565399, 2.662079, 2.862122, 2.657104, 2.611633, 2.523743, 
    2.366058, 2.451324, 2.654327, 2.778442, 2.987488, 3.154419, 2.051636, 
    1.973297, 2.119507, 2.169952, 1.600861, 1.364594, 0.9707947, 0.5310059, 
    0.5891418, 0.9031677, 1.023315, 0.8419495, 0.4814758, 0.4241333, 
    0.673645, 0.9885254, 1.177917, 1.279266, 1.465393, 1.792999,
  0.9830017, 1.235168, 1.664185, 1.91864, 1.967682, 1.723877, 2.006927, 
    1.889435, 2.064758, 2.004669, 1.823334, 1.728027, 1.934418, 2.207397, 
    2.478363, 2.728363, 2.925293, 3.169037, 3.530365, 3.80719, 4.060913, 
    3.886993, 3.945923, 3.892609, 3.897308, 4.063782, 4.069397, 3.919891, 
    3.785583, 3.852966, 3.786926, 3.901276, 4.048218, 3.907867, 3.665924, 
    3.695801, 3.721466, 3.72348, 3.952759, 3.847046, 3.67984, 3.84256, 
    3.623474, 3.502441, 3.47998, 3.699341, 3.24353, 2.417267, 2.75531, 
    3.103333, 3.280701, 3.23941, 3.323547, 3.283112, 3.258026, 3.214172, 
    3.13266, 3.200531, 3.129089, 2.974884, 2.943909, 3.151123, 3.154846, 
    2.863373, 2.36618, 2.249725, 2.494629, 2.551727, 2.501343, 2.273865, 
    2.003418, 2.277222, 2.382843, 2.345428, 2.240479, 2.058044, 1.76825, 
    2.012329, 1.989929, 1.738403, 1.3367, 0.9928589, 0.740509, 0.571991, 
    0.639801, 0.4050903, 0.6620178, 0.9717712, 1.151184, 1.23233, 1.209229, 
    1.003632, 0.697052, 0.5619507, 0.7999573, 0.9501038,
  0.3583679, 0.3652649, 0.6296387, 1.518188, 1.835968, 2.021667, 1.359802, 
    2.152496, 2.119171, 2.08551, 1.984406, 1.893158, 1.982727, 2.229004, 
    2.476257, 2.723846, 2.882507, 3.068542, 3.18634, 3.257019, 3.319214, 
    3.410767, 3.52771, 3.583344, 3.840393, 4.287903, 4.522736, 4.581818, 
    4.37027, 4.011475, 3.88916, 3.786316, 3.724121, 3.686249, 3.766571, 
    3.763794, 3.669495, 3.886505, 3.17868, 3.217407, 3.597076, 3.683228, 
    3.371307, 3.355499, 3.1922, 3.131683, 3.292603, 3.284424, 3.052917, 
    3.117279, 3.067627, 2.813049, 3.139862, 3.187439, 3.276855, 3.380371, 
    3.468842, 3.662811, 3.646515, 3.412384, 3.084473, 3.033478, 2.926636, 
    2.781616, 2.667358, 2.549744, 2.53064, 2.492035, 2.294617, 2.115448, 
    2.22998, 2.335327, 2.663574, 2.72757, 1.524323, 1.503937, 1.417664, 
    2.201019, 2.411621, 2.262604, 1.263062, 1.070618, 1.807068, 2.125336, 
    2.47757, 2.512238, 1.797699, 1.015442, 0.9535522, 1.103302, 1.096527, 
    1.359009, 0.8012695, 0.4092102, 0.2433777, 0.1968994,
  0.7383728, 0.6754761, 0.5969849, 0.4753418, 0.208313, 1.621521, 1.92569, 
    2.13266, 2.272888, 2.183899, 2.086334, 1.622345, 1.630249, 1.704987, 
    2.505493, 2.70575, 2.99295, 3.146088, 3.251587, 3.453949, 3.652313, 
    3.701447, 3.858765, 4.027466, 4.104004, 4.366241, 4.539612, 4.520538, 
    4.362793, 4.319214, 4.133484, 3.918701, 3.573273, 3.462921, 3.240601, 
    3.35199, 3.434906, 3.374573, 3.197693, 2.867432, 2.331665, 2.026062, 
    1.750488, 1.687469, 1.817566, 2.010132, 2.125488, 2.161987, 2.188171, 
    1.578613, 1.891113, 2.105835, 2.207733, 2.837006, 2.940338, 3.056824, 
    3.180176, 3.279419, 3.465729, 2.935822, 2.758057, 2.666565, 2.546906, 
    2.481476, 2.534454, 2.582123, 2.622894, 2.679901, 2.577301, 1.743073, 
    2.558044, 2.49234, 2.483246, 1.233246, 2.256958, 1.178955, 1.885773, 
    2.009613, 1.811951, 1.233215, 1.223785, 1.188171, 2.176392, 3.937866, 
    4.045929, 4.212677, 3.935211, 3.61853, 3.229675, 2.340515, 1.499054, 
    1.299774, 0.9437866, 0.9256592, 0.9025574, 0.8735352,
  1.43576, 1.279633, 1.117157, 0.9373169, 0.7488708, 0.9204102, 1.485443, 
    1.983368, 2.172821, 2.124908, 1.945221, 1.852814, 1.774689, 1.706177, 
    1.552185, 2.02124, 1.544067, 1.678864, 1.810059, 2.914764, 3.301025, 
    3.483368, 3.619629, 3.874847, 4.127258, 4.363831, 4.468842, 4.548859, 
    4.538574, 4.188721, 3.956146, 3.577057, 3.206879, 2.987793, 2.704315, 
    0.9868774, 1.071564, 1.085114, 2.133209, 1.86969, 0.9072876, 0.7790222, 
    0.6445618, 0.6174316, 0.5911865, 0.5834961, 0.6156006, 0.6564941, 
    0.7218018, 0.7592773, 0.8694458, 0.9210815, 0.8680115, 0.8225098, 
    0.8540955, 0.8892517, 0.9293518, 0.9804993, 1.033081, 1.065033, 1.09436, 
    1.229126, 1.445496, 2.178162, 2.323395, 2.521851, 2.703369, 2.662872, 
    2.549713, 1.52948, 2.023071, 1.718201, 0.918396, 1.44809, 1.545166, 
    1.793518, 1.822632, 1.522461, 1.451874, 1.477051, 1.448456, 2.206421, 
    3.943268, 4.249207, 4.682007, 5.089752, 4.695084, 4.150818, 3.870605, 
    3.593658, 2.485931, 1.733307, 1.505585, 1.332794, 1.345001, 1.456818,
  1.457703, 1.442291, 1.674255, 1.951508, 2.005676, 2.061951, 2.208374, 
    2.225952, 2.088348, 1.904144, 1.762878, 1.684814, 1.645996, 1.562347, 
    1.419006, 1.312134, 1.260345, 1.172577, 1.139435, 1.137238, 1.141602, 
    1.189362, 1.244659, 1.298096, 1.427673, 2.555634, 2.677124, 2.892426, 
    2.845978, 2.611877, 2.419891, 1.164001, 1.137024, 1.029938, 1.048767, 
    0.9980469, 0.9378052, 0.9051208, 0.9231567, 0.8785095, 0.8141174, 
    0.7926941, 0.7842407, 0.7952881, 0.817627, 0.8480225, 0.8780823, 
    0.894043, 0.8948364, 0.9119263, 0.9495239, 1.021332, 1.101685, 1.15213, 
    1.18399, 1.223877, 1.269196, 1.33728, 1.364044, 1.315491, 1.217041, 
    1.149323, 1.166382, 1.3479, 1.590881, 1.770081, 1.832611, 1.845215, 
    1.900482, 1.818909, 1.676605, 1.467407, 1.505646, 1.641815, 1.750732, 
    1.798553, 1.963013, 1.85141, 3.374512, 3.405853, 3.552277, 3.877869, 
    4.256226, 4.507919, 4.487488, 4.549591, 4.639053, 4.394073, 4.156097, 
    3.989044, 3.756042, 2.48175, 1.674835, 1.44223, 1.476227, 1.510193,
  1.513458, 1.507874, 1.670685, 1.691956, 2.455322, 2.482666, 2.477997, 
    1.88385, 1.740112, 1.624512, 1.514954, 1.383759, 1.274475, 1.212524, 
    1.177216, 1.149719, 1.128021, 1.085602, 1.06073, 1.06723, 1.057587, 
    1.07132, 1.062408, 1.084625, 1.114105, 2.219513, 2.204742, 1.360077, 
    1.372833, 1.390747, 1.351654, 1.285522, 1.204407, 1.172211, 1.168915, 
    1.177307, 1.235992, 1.303101, 1.344818, 1.351685, 1.324554, 1.322815, 
    1.33902, 1.35025, 1.375702, 1.413513, 1.446472, 1.491974, 1.544983, 
    1.592255, 1.61795, 1.666992, 1.711548, 1.736511, 1.783173, 1.838959, 
    1.882141, 1.93338, 1.993927, 2.112213, 2.19986, 2.248413, 2.291534, 
    2.331482, 2.325836, 2.291077, 2.221985, 2.173279, 2.152802, 2.221802, 
    2.114563, 2.631836, 3.123993, 3.279755, 3.314819, 3.222565, 3.191193, 
    3.271606, 3.39856, 3.601349, 3.68631, 3.752502, 3.85434, 3.848389, 
    3.845459, 3.826904, 3.703735, 3.575043, 3.60376, 3.650055, 3.799927, 
    3.807251, 2.20993, 1.962067, 1.693787, 1.579987,
  2.98703, 2.844727, 2.741608, 2.669434, 2.644043, 2.54184, 2.42453, 
    2.307556, 2.227203, 2.138458, 2.100067, 2.073883, 2.040955, 2.001892, 
    1.968475, 1.95871, 1.957733, 1.97226, 1.965363, 1.942444, 1.918152, 
    1.875061, 1.858856, 1.841248, 1.835999, 1.833893, 1.811951, 1.802002, 
    1.770233, 1.707092, 1.644958, 1.621185, 1.621063, 1.636261, 1.655243, 
    1.684906, 1.727386, 1.790741, 1.831116, 1.845703, 1.856445, 1.86438, 
    1.890869, 1.919067, 1.94342, 1.956299, 1.95343, 1.945251, 1.907745, 
    1.882477, 1.871399, 1.838806, 1.843994, 1.870056, 1.915985, 1.998077, 
    2.081757, 2.200623, 2.291962, 2.401367, 2.509796, 2.597229, 2.708191, 
    2.808502, 2.875427, 2.92099, 2.93161, 2.876038, 2.806427, 2.809998, 
    2.895752, 3.010986, 3.109283, 3.162933, 3.333649, 3.444458, 3.609375, 
    3.808838, 4.091064, 4.308105, 4.580109, 4.78363, 5.036194, 5.187012, 
    5.271423, 5.261505, 5.240784, 5.133118, 4.940735, 4.649597, 4.297363, 
    3.807922, 3.533508, 3.41449, 3.288086, 3.168915,
  3.13208, 3.079865, 3.087097, 3.11731, 3.088074, 3.057678, 3.006409, 
    2.931732, 2.872375, 2.800964, 2.741852, 2.680206, 2.631561, 2.598541, 
    2.545166, 2.494385, 2.452911, 2.421967, 2.397247, 2.365204, 2.334015, 
    2.310211, 2.287354, 2.289429, 2.257721, 2.229919, 2.220551, 2.21228, 
    2.198669, 2.202667, 2.194794, 2.206177, 2.214691, 2.251984, 2.247955, 
    2.243195, 2.232605, 2.245544, 2.229736, 2.234253, 2.237701, 2.236572, 
    2.254669, 2.262787, 2.287079, 2.298553, 2.339844, 2.350708, 2.379761, 
    2.397369, 2.426025, 2.449402, 2.489716, 2.541077, 2.582092, 2.649597, 
    2.721191, 2.765656, 2.792816, 2.836639, 2.877625, 2.941315, 3.012543, 
    3.068604, 3.159821, 3.233398, 3.292358, 3.328491, 3.383118, 3.437286, 
    3.496704, 3.541595, 3.577911, 3.638336, 3.686249, 3.742371, 3.806519, 
    3.888458, 3.939789, 3.972626, 4.031555, 4.043732, 4.006165, 4.006378, 
    4.004822, 3.972321, 3.90564, 3.839813, 3.747131, 3.6427, 3.569, 3.478119, 
    3.415009, 3.340942, 3.277466, 3.220306,
  1.768158, 1.774033, 1.785797, 1.803329, 1.824081, 1.848831, 1.877808, 
    1.913086, 1.953186, 1.995255, 2.04335, 2.094009, 2.151169, 2.206451, 
    2.261261, 2.313339, 2.362366, 2.409515, 2.449097, 2.487045, 2.521027, 
    2.550079, 2.57663, 2.598953, 2.619278, 2.636124, 2.649933, 2.657684, 
    2.658203, 2.652664, 2.640503, 2.623764, 2.605728, 2.584702, 2.554749, 
    2.52597, 2.497925, 2.469666, 2.439835, 2.411392, 2.38118, 2.350067, 
    2.321426, 2.292892, 2.265945, 2.240814, 2.233398, 2.203186, 2.185944, 
    2.180801, 2.16803, 2.16745, 2.20639, 2.241867, 2.217712, 2.259369, 
    2.287964, 2.289642, 2.290939, 2.238602, 2.267975, 2.306442, 2.286652, 
    2.312241, 2.32103, 2.321945, 2.336197, 2.350845, 2.367706, 2.34967, 
    2.343033, 2.349152, 2.380783, 2.489258, 2.31517, 2.270309, 2.271286, 
    2.314651, 2.194077, 2.145889, 2.114777, 2.089584, 2.071091, 2.045181, 
    2.017578, 1.994461, 1.969589, 1.945435, 1.920624, 1.893677, 1.868607, 
    1.846939, 1.819794, 1.798111, 1.78392, 1.771622,
  1.656067, 1.6931, 1.73764, 1.789063, 1.876556, 1.993103, 2.138489, 
    2.310028, 2.470581, 2.601166, 2.705017, 2.78392, 2.836334, 2.8638, 
    2.879623, 2.89856, 2.914261, 2.936127, 2.971222, 3.011841, 3.03157, 
    3.038086, 3.023239, 2.980087, 2.911331, 2.836517, 2.796738, 2.767181, 
    2.731628, 2.680405, 2.616669, 2.557617, 2.501877, 2.451172, 2.410675, 
    2.383591, 2.365234, 2.350906, 2.342056, 2.341599, 2.362167, 2.393494, 
    2.432281, 2.478394, 2.540878, 2.640228, 2.678909, 2.731964, 2.776169, 
    2.822266, 2.836975, 2.851563, 2.836777, 2.811523, 2.808334, 2.714706, 
    2.673767, 2.637115, 2.577087, 2.52507, 2.465622, 2.432617, 2.417068, 
    2.428452, 2.455399, 2.498703, 2.589966, 2.673431, 2.740494, 2.772324, 
    2.779617, 2.732483, 2.592911, 2.44368, 2.294403, 2.149933, 2.034241, 
    1.912369, 1.89389, 1.841476, 1.7677, 1.704041, 1.597855, 1.514252, 
    1.323639, 1.233459, 1.256638, 1.24942, 1.257431, 1.293747, 1.348892, 
    1.409958, 1.472214, 1.533401, 1.587448, 1.62532,
  1.111786, 1.211914, 1.433655, 1.694778, 2.020889, 2.325775, 2.586517, 
    2.762695, 2.813477, 2.753067, 2.671356, 2.653763, 2.598694, 2.538483, 
    2.53093, 2.555923, 2.57637, 2.586838, 2.567261, 2.527863, 2.543365, 
    2.693024, 2.941223, 3.085556, 3.00116, 2.843826, 2.846359, 2.937378, 
    3.0065, 2.995575, 2.88588, 2.700394, 2.479935, 2.315887, 2.24382, 
    2.232422, 2.249741, 2.256256, 2.265045, 2.28418, 2.294266, 2.36145, 
    2.504227, 2.748108, 3.24205, 3.602081, 3.768494, 3.769135, 3.778778, 
    3.758194, 3.708908, 3.676041, 3.682037, 3.725006, 3.671814, 3.515701, 
    3.34993, 3.041672, 2.632095, 2.357742, 2.239334, 2.259308, 2.424149, 
    2.665375, 2.929688, 3.135605, 3.184235, 3.205734, 3.127151, 2.99173, 
    2.663025, 2.362961, 2.098633, 1.921555, 1.817841, 1.752853, 1.758133, 
    1.778519, 1.821487, 1.89238, 1.980789, 2.026428, 1.930344, 1.807159, 
    1.597855, 1.487961, 1.406708, 1.29628, 1.265564, 1.243423, 1.298248, 
    1.33548, 1.372787, 1.322723, 1.239059, 1.143951,
  1.570847, 1.590958, 1.701492, 1.919083, 2.185745, 2.368027, 2.372986, 
    2.260742, 2.180466, 2.183792, 2.188934, 2.217377, 2.276367, 2.361206, 
    2.516083, 2.761795, 2.986389, 3.247452, 3.306519, 2.744003, 1.982544, 
    1.589523, 1.50592, 1.61412, 1.732162, 1.782486, 2.017776, 2.232361, 
    2.350647, 2.353134, 2.280472, 2.195053, 2.111908, 1.952271, 1.703644, 
    1.339447, 1.103897, 1.105988, 1.282288, 1.453583, 1.613998, 1.751297, 
    1.872269, 1.974731, 2.108734, 2.497864, 1.989334, 1.696152, 1.668884, 
    1.574142, 1.719543, 1.867447, 2.048828, 2.152863, 2.287567, 2.407623, 
    2.206451, 2.877075, 2.620255, 2.312378, 2.132935, 2.045898, 2.084381, 
    2.083649, 2.111465, 2.155411, 2.173767, 2.194397, 2.250381, 2.233261, 
    2.191147, 2.138809, 2.156448, 2.225784, 2.3517, 2.52005, 2.695831, 
    2.875641, 3.004684, 3.010223, 2.730728, 2.779297, 2.671356, 2.614777, 
    2.545761, 2.454041, 2.475662, 2.417633, 2.335678, 1.660675, 1.364914, 
    1.264908, 1.305588, 1.350525, 1.422333, 1.518997,
  1.725006, 1.696228, 1.72937, 1.830795, 1.965103, 2.132935, 2.273636, 
    2.334442, 2.336395, 2.289719, 2.275131, 2.263611, 2.309692, 2.367325, 
    2.45105, 2.248825, 2.123901, 2.003448, 1.985809, 2.083328, 1.897079, 
    1.597916, 1.404022, 1.436203, 1.658325, 1.747528, 1.620758, 1.626572, 
    1.684036, 1.842575, 1.998901, 2.00383, 1.943802, 1.952667, 1.976364, 
    2.002472, 2.018814, 1.90274, 1.589981, 1.323441, 1.21022, 1.306244, 
    1.41777, 1.520828, 1.59343, 1.740692, 1.212234, 1.328125, 1.333725, 
    1.3759, 1.519989, 1.738541, 1.844925, 1.941864, 2.003845, 1.997406, 
    1.917252, 1.734238, 1.78241, 1.840958, 1.994797, 2.056061, 2.044006, 
    2.109894, 2.107819, 2.116989, 2.143616, 2.173645, 2.144852, 1.931244, 
    2.604813, 2.667908, 2.636658, 2.705139, 2.737701, 2.638412, 3.0336, 
    3.228058, 3.385605, 3.301575, 3.148636, 2.885147, 2.638016, 2.432159, 
    2.442383, 2.469009, 2.500717, 2.58223, 2.681519, 2.726242, 2.892441, 
    2.835876, 2.336533, 2.060608, 1.976379, 1.822983,
  3.554626, 2.984772, 2.675064, 2.221741, 2.025131, 2.008865, 2.202347, 
    2.585739, 2.699478, 2.783325, 2.874863, 2.659576, 2.330734, 2.154297, 
    2.055405, 1.909775, 1.803253, 1.815826, 1.797134, 1.714844, 1.619598, 
    1.412247, 1.118362, 1.019455, 1.06218, 1.034698, 1.058533, 1.085159, 
    1.126755, 1.158401, 1.207489, 1.19342, 1.199295, 1.254166, 1.306961, 
    1.242767, 1.179886, 1.103851, 1.060944, 1.040756, 1.118942, 1.228577, 
    1.205734, 1.177994, 1.251114, 1.283066, 1.287766, 1.341873, 1.40332, 
    1.497131, 1.688156, 1.909897, 2.018494, 2.115158, 2.186523, 2.232559, 
    2.215164, 2.147278, 2.146103, 2.218887, 2.330658, 2.411789, 2.495316, 
    2.491867, 2.488281, 2.384445, 2.346161, 2.37442, 2.504166, 2.725266, 
    3.074417, 3.417053, 3.605209, 3.681976, 3.480728, 3.200195, 2.871994, 
    2.673752, 3.093491, 3.039444, 2.956863, 2.75769, 2.54039, 2.402222, 
    2.45578, 2.568222, 2.771881, 2.908981, 2.923248, 2.882874, 2.990097, 
    3.120895, 3.248627, 3.406372, 3.436722, 3.574081,
  3.457626, 3.594604, 3.558273, 3.572388, 3.402939, 3.147797, 2.985687, 
    2.877808, 2.793427, 2.842972, 3.000183, 3.100128, 3.245651, 3.332611, 
    3.106186, 2.924484, 2.750061, 2.559769, 2.500458, 2.568741, 2.65892, 
    2.627075, 2.482742, 2.287231, 1.945892, 1.838928, 1.83255, 1.714645, 
    1.313858, 0.8141327, 0.3233795, 0.06718445, -0.0145874, 0.87883, 
    1.267838, 1.704041, 2.089264, 2.376175, 2.577545, 2.661911, 2.672073, 
    2.610764, 2.50795, 2.496674, 2.469711, 2.356537, 2.313873, 2.065674, 
    1.603119, 1.093567, 0.9540405, 0.8360596, 0.8547974, 1.056122, 1.375397, 
    1.657379, 1.812256, 1.865326, 1.967316, 2.104828, 2.353729, 2.605103, 
    2.876434, 3.131409, 3.329453, 3.618195, 3.805359, 4.014526, 4.358673, 
    4.558167, 4.887146, 5.54657, 5.552795, 5.828583, 5.223511, 4.892639, 
    4.338013, 3.706055, 3.268951, 3.157776, 3.124542, 3.113434, 3.180481, 
    3.157104, 3.150192, 3.204239, 3.368103, 3.473953, 3.515808, 3.526047, 
    3.476822, 3.446411, 3.37291, 3.375137, 3.377014, 3.378326,
  3.594421, 3.629501, 3.754547, 3.992844, 4.210037, 4.057358, 3.920837, 
    3.742584, 3.617966, 3.583557, 3.760818, 3.867996, 4.279449, 4.555618, 
    4.885818, 4.749222, 4.226593, 4.312424, 4.433075, 4.358917, 4.470764, 
    4.270828, 3.94075, 3.509903, 3.037506, 2.613098, 2.540314, 2.463547, 
    2.134964, 1.397705, 0.2570496, 0.560791, 0.8311157, 0.934906, 1.233398, 
    2.428009, 3.017181, 2.805725, 2.993988, 2.507355, 2.525574, 2.414734, 
    2.26178, 2.509705, 2.719055, 2.814056, 2.475769, 1.383789, 0.05697632, 
    -1.132355, -1.661591, -1.634033, -1.624023, -1.570099, -1.321106, 
    -0.903595, -0.4160156, -0.2520142, 0.1360779, 0.8233032, 1.672974, 
    2.511993, 3.040955, 3.406311, 3.955963, 4.578857, 4.646698, 4.476227, 
    4.344543, 4.140442, 4.104034, 4.15686, 4.24707, 4.697601, 5.026123, 
    4.955078, 4.446808, 4.093414, 3.757874, 3.253326, 3.23175, 3.705078, 
    3.870636, 3.804749, 3.586853, 3.482239, 3.536346, 3.717651, 3.928894, 
    4.056519, 4.212036, 4.134186, 3.95816, 3.774811, 3.634171, 3.604156,
  4.607361, 4.829956, 4.839935, 5.059174, 5.314514, 5.436401, 5.131561, 
    4.591461, 4.495636, 4.461914, 3.831635, 3.739594, 4.058533, 4.803528, 
    5.323425, 5.630524, 5.880402, 6.322479, 6.61972, 6.795898, 6.482544, 
    5.906067, 5.06015, 4.123291, 3.263947, 2.705536, 2.613464, 2.548218, 
    2.525116, 2.163361, 1.901001, 1.466705, 1.123169, 1.005585, 0.9934998, 
    1.177612, 1.565704, 1.77832, 1.800507, 1.791534, 2.0336, 2.419312, 
    2.818604, 2.886261, 2.58847, 2.375854, 2.204498, 1.855072, 0.8613892, 
    0.09338379, -0.07168579, -0.0859375, -0.1645203, -0.3336487, -0.4947205, 
    -0.5990295, -0.6495972, -0.4470825, 0.04830933, 0.5502014, 0.9768066, 
    1.254486, 1.441711, 1.692841, 1.850586, 1.972534, 2.187439, 2.304871, 
    2.278656, 2.385376, 2.472595, 2.386261, 2.364319, 2.378143, 2.319397, 
    2.09668, 1.691528, 1.573608, 1.595428, 1.603271, 1.643341, 1.743073, 
    1.954437, 2.145355, 2.417053, 2.81131, 3.148163, 3.59082, 3.832031, 
    4.017853, 4.2146, 4.450592, 4.640442, 4.600769, 4.559235, 4.55307,
  3.295837, 3.429688, 3.655273, 3.557709, 3.219391, 3.115112, 3.096802, 
    3.055481, 2.947723, 2.671448, 2.551941, 2.508087, 2.530884, 2.691223, 
    3.003784, 3.401001, 3.720123, 4.071503, 4.424286, 4.514709, 4.483337, 
    4.092499, 3.709778, 2.905792, 2.343628, 2.224854, 2.321991, 2.401947, 
    2.366669, 2.235809, 1.993439, 1.642181, 1.395203, 1.31308, 1.396881, 
    1.603638, 1.901031, 2.119324, 2.162628, 2.036652, 2.099609, 2.455078, 
    2.688751, 2.5177, 2.096619, 1.977997, 1.992126, 1.960419, 1.572601, 
    1.140106, 0.8806152, 0.6891174, 0.5393372, 0.4085388, 0.3113708, 
    0.2590332, 0.2894592, 0.4266357, 0.6394653, 0.8527527, 1.016174, 
    1.119812, 1.208984, 1.280151, 1.324677, 1.37973, 1.473511, 1.612244, 
    1.69751, 1.767334, 1.8349, 1.847778, 1.785675, 1.669189, 1.418549, 
    1.126617, 1.250793, 2.034698, 2.087952, 1.404053, 1.335419, 1.423828, 
    1.795013, 1.696991, 1.674469, 1.959381, 2.518005, 3.009888, 3.371155, 
    3.728119, 3.987946, 4.110413, 3.943451, 3.68042, 3.250702, 3.131775,
  2.15274, 2.303711, 2.404938, 2.419922, 2.413544, 2.432343, 2.508179, 
    2.589447, 2.628174, 2.589386, 2.608551, 2.70874, 2.748566, 2.724884, 
    2.756958, 2.855225, 3.09024, 3.452942, 3.672577, 3.519348, 3.309387, 
    3.316528, 3.263306, 2.997986, 2.76355, 2.711395, 2.753387, 2.763458, 
    2.751678, 2.65567, 2.424927, 2.079102, 1.790497, 1.719208, 1.819092, 
    1.923889, 1.948334, 1.861572, 1.743622, 1.788422, 2.091278, 2.435547, 
    2.488831, 2.193909, 2.140076, 2.13382, 2.040192, 1.973511, 1.831818, 
    1.477722, 1.150208, 0.9937439, 0.9768372, 0.9889832, 0.9595032, 
    0.9195251, 0.9360962, 1.039734, 1.202545, 1.295959, 1.303101, 1.314392, 
    1.342834, 1.342438, 1.31958, 1.29361, 1.331299, 1.370361, 1.365692, 
    1.362488, 1.373291, 1.334229, 1.254669, 1.138214, 1.010345, 1.140961, 
    1.80603, 2.22702, 1.911652, 1.633636, 1.339447, 1.355469, 1.755859, 
    1.870514, 1.712311, 1.743164, 1.956604, 2.195984, 2.370422, 2.50061, 
    2.505707, 2.40976, 2.334198, 2.290894, 2.212769, 2.116669,
  2.14917, 2.301422, 2.42688, 2.507385, 2.568298, 2.677155, 2.882813, 
    3.081879, 3.142181, 3.236603, 3.443817, 3.545837, 3.490875, 3.368958, 
    3.239777, 3.084961, 3.016479, 3.238403, 3.477753, 3.725403, 4.168518, 
    4.415466, 4.102051, 3.53363, 3.168793, 2.998596, 2.845459, 2.709625, 
    2.604675, 2.41626, 2.134216, 1.894379, 1.787933, 1.786621, 1.793274, 
    1.703064, 1.515076, 1.323547, 1.240021, 1.388824, 1.947174, 2.39444, 
    2.445679, 2.249847, 2.502686, 2.43573, 2.207306, 2.044617, 1.969818, 
    1.847809, 1.735901, 1.710114, 1.692078, 1.630371, 1.591888, 1.586426, 
    1.543518, 1.510651, 1.548401, 1.594116, 1.583679, 1.536407, 1.452728, 
    1.389191, 1.346466, 1.284576, 1.243683, 1.21756, 1.179291, 1.128967, 
    1.116364, 1.104767, 1.079102, 1.060822, 1.031616, 1.096863, 1.518311, 
    1.955017, 1.839935, 1.626373, 1.455688, 1.438049, 1.721161, 1.7117, 
    1.544006, 1.551483, 1.690887, 1.90274, 2.090302, 2.145844, 2.106842, 
    2.063416, 2.023621, 1.983093, 1.976318, 2.032349,
  2.415955, 2.547882, 2.626068, 2.593781, 2.579315, 2.932373, 3.643066, 
    4.136902, 4.262451, 4.389862, 4.54776, 4.434479, 3.970673, 3.560638, 
    3.272705, 3.036041, 2.923645, 2.993347, 3.183411, 3.384369, 3.480591, 
    3.318054, 2.87738, 2.386353, 2.12146, 1.999756, 1.906403, 1.792938, 
    1.67868, 1.585907, 1.543457, 1.576141, 1.533752, 1.347168, 1.131653, 
    1.04071, 1.090668, 1.22348, 1.435974, 1.607178, 2.049652, 2.481476, 
    2.453491, 2.31958, 2.602173, 2.825226, 2.354279, 2.214355, 2.264496, 
    2.377777, 2.548584, 2.492279, 2.265533, 2.016052, 1.861664, 1.798096, 
    1.67926, 1.577698, 1.611084, 1.663849, 1.642151, 1.538574, 1.444427, 
    1.418121, 1.370148, 1.292206, 1.283234, 1.263763, 1.247894, 1.299835, 
    1.320221, 1.315796, 1.33136, 1.307648, 1.209473, 1.091827, 1.148804, 
    1.281525, 1.402405, 1.593201, 1.518524, 1.505402, 1.678162, 1.832001, 
    1.871948, 1.92627, 2.042419, 2.177063, 2.349701, 2.367737, 2.249268, 
    2.198853, 2.165771, 2.117798, 2.163116, 2.274384,
  2.350037, 2.29892, 2.211517, 2.210297, 2.489288, 3.148529, 3.457825, 
    3.545105, 3.628082, 3.440399, 2.977051, 2.591675, 2.243134, 2.019104, 
    1.908905, 1.894623, 1.887878, 1.890869, 1.920868, 1.851929, 1.695404, 
    1.470795, 1.209869, 1.058563, 0.9987793, 0.9903259, 1.014557, 1.008057, 
    1.167664, 1.740204, 2.02417, 1.755554, 1.424103, 1.009216, 0.8463135, 
    1.190308, 1.501587, 1.542297, 1.696655, 1.839752, 2.0495, 2.562927, 
    2.824646, 2.574768, 2.597534, 2.771759, 2.674316, 2.315277, 2.397369, 
    2.280823, 2.093414, 1.95752, 1.862335, 1.718781, 1.618439, 1.559296, 
    1.475494, 1.43689, 1.528656, 1.611237, 1.601776, 1.578033, 1.584076, 
    1.6008, 1.583557, 1.548279, 1.552643, 1.536438, 1.586731, 1.632965, 
    1.597931, 1.580109, 1.5495, 1.446198, 1.326782, 1.189545, 1.136566, 
    1.379364, 1.693451, 1.573944, 1.578339, 1.684204, 2.141876, 2.488068, 
    2.699188, 2.713776, 2.632843, 2.582123, 2.520599, 2.361145, 2.270599, 
    2.272217, 2.294098, 2.285004, 2.268585, 2.304199,
  1.963043, 1.935699, 1.964539, 2.118927, 2.366364, 2.456299, 2.398651, 
    2.353882, 2.718201, 2.344604, 1.546692, 1.414093, 1.473541, 1.473511, 
    1.37085, 1.325897, 1.315308, 1.233307, 1.080505, 0.8228455, 0.6294556, 
    0.6255493, 0.7017212, 0.8544006, 1.039154, 1.212158, 1.422882, 1.737976, 
    2.305542, 2.515961, 1.785309, 1.692627, 1.652313, 1.520599, 1.512665, 
    1.575806, 1.559357, 1.564606, 1.744232, 1.745453, 1.183838, 2.703308, 
    3.455627, 3.233887, 2.970856, 2.966248, 2.659668, 2.223755, 1.928101, 
    1.462524, 1.190521, 1.184418, 1.206635, 1.229797, 1.299561, 1.378082, 
    1.442535, 1.523346, 1.639282, 1.740784, 1.770874, 1.780548, 1.802307, 
    1.83844, 1.833557, 1.797546, 1.771973, 1.767609, 1.775085, 1.717529, 
    1.631042, 1.568512, 1.456543, 1.337921, 1.275543, 1.086365, 1.078278, 
    1.954437, 2.326752, 1.838104, 1.903076, 2.212463, 2.640686, 2.948669, 
    2.507385, 2.335907, 2.332642, 2.271515, 2.096771, 1.978668, 1.999847, 
    2.047363, 1.980103, 1.93335, 1.922241, 1.930542,
  1.799561, 1.757507, 1.765289, 1.798096, 1.937134, 3.210968, 3.809784, 
    4.096832, 3.880585, 2.350891, 2.047852, 2.027679, 1.947144, 1.86145, 
    1.807281, 1.787872, 1.783752, 1.706024, 1.631165, 1.625732, 1.741486, 
    1.886108, 1.991119, 2.089233, 2.19812, 2.311615, 2.491913, 2.648743, 
    2.582397, 2.015503, 1.753723, 3.199646, 2.349701, 1.716705, 1.868378, 
    1.529205, 1.595032, 1.530029, 1.27301, 1.455627, 1.226868, 2.267365, 
    2.289063, 2.468719, 2.558838, 2.537292, 2.146393, 1.565918, 1.264679, 
    1.092468, 1.135345, 1.352173, 1.532257, 1.607056, 1.67218, 1.686371, 
    1.692932, 1.735138, 1.762665, 1.814484, 1.845276, 1.856873, 1.823334, 
    1.823029, 1.822449, 1.787537, 1.72049, 1.639099, 1.539368, 1.438354, 
    1.339905, 1.258057, 1.169159, 1.143372, 1.089294, 0.9008789, 1.155579, 
    2.684296, 3.206787, 2.3508, 2.095367, 2.625549, 2.867035, 2.641388, 
    2.345428, 2.055389, 2.011841, 1.924957, 1.971741, 1.974823, 1.868317, 
    1.833923, 1.803741, 1.802765, 1.801788, 1.796753,
  1.620087, 1.608185, 1.720734, 1.939087, 2.404602, 3.809814, 4.504791, 
    4.655426, 3.941284, 2.455933, 2.175323, 2.33606, 2.39447, 2.293365, 
    2.470642, 2.549927, 2.606812, 2.581299, 2.519409, 2.521423, 2.484497, 
    2.473633, 2.45813, 2.456726, 2.453522, 2.383667, 2.347046, 2.169983, 
    1.999664, 1.878174, 1.928894, 3.27124, 2.580383, 2.256165, 2.240021, 
    1.840149, 1.817871, 1.602386, 1.210693, 1.248444, 1.076721, 1.623505, 
    1.500397, 1.592773, 1.74881, 1.735138, 1.682343, 1.722382, 1.745239, 
    1.85202, 1.914063, 1.911591, 1.872589, 1.80545, 1.748169, 1.669586, 
    1.627136, 1.617279, 1.614502, 1.649353, 1.641327, 1.610016, 1.570953, 
    1.573944, 1.578644, 1.529144, 1.471161, 1.383026, 1.299957, 1.238953, 
    1.149384, 1.119904, 1.094238, 0.9893799, 0.8319397, 0.9347229, 1.657135, 
    3.484863, 4.313873, 2.932129, 2.808563, 3.379395, 3.564545, 3.52066, 
    2.577545, 1.985748, 1.885132, 1.988861, 1.961243, 1.882477, 1.799652, 
    1.777985, 1.773376, 1.733215, 1.642609, 1.634979,
  1.65387, 1.848419, 2.10141, 2.576416, 4.153137, 4.258667, 4.464539, 
    4.794281, 4.611481, 4.190277, 2.281372, 2.470428, 4.015503, 2.433411, 
    2.405731, 2.547516, 2.452698, 2.452423, 2.339264, 2.249023, 2.166748, 
    2.135864, 2.079803, 2.068756, 2.075287, 2.046875, 2.02475, 1.948578, 
    1.923615, 1.999908, 2.098877, 3.317291, 3.148834, 2.992035, 2.72052, 
    1.907043, 1.559937, 1.315308, 1.452484, 1.371796, 1.191162, 1.652924, 
    1.825073, 1.977081, 2.060211, 2.040833, 2.016144, 2.068665, 2.024994, 
    1.947601, 1.86908, 1.791016, 1.724243, 1.646027, 1.568634, 1.551514, 
    1.520386, 1.496613, 1.523895, 1.548889, 1.548889, 1.542969, 1.544525, 
    1.546692, 1.528107, 1.399872, 1.349152, 1.285492, 1.235291, 1.142487, 
    1.115112, 1.108856, 1.011047, 0.8818054, 0.9941101, 1.433502, 2.337891, 
    4.277191, 4.750793, 3.486206, 4.559753, 5.236572, 5.329803, 4.335022, 
    4.349762, 2.1828, 1.723053, 1.819031, 1.779633, 1.684784, 1.636871, 
    1.559845, 1.518402, 1.486084, 1.455933, 1.539398,
  2.008667, 2.225128, 2.353302, 2.715393, 4.757172, 4.838074, 4.746216, 
    4.66861, 4.503967, 4.546082, 2.378143, 2.419769, 3.921143, 3.230469, 
    2.220703, 2.293762, 2.223816, 2.18457, 2.087891, 2.02832, 1.999878, 
    2.00943, 2.037964, 2.082886, 2.14447, 2.131134, 2.090759, 2.039856, 
    2.054352, 2.18866, 2.257111, 2.333862, 3.332031, 3.084839, 2.314575, 
    1.97467, 1.828583, 1.963348, 2.160217, 1.878784, 1.944916, 2.107819, 
    2.2901, 2.354553, 2.267883, 2.182159, 2.081909, 1.978302, 1.897064, 
    1.820648, 1.803528, 1.754272, 1.700562, 1.673828, 1.677795, 1.686127, 
    1.6633, 1.714996, 1.78006, 1.829437, 1.889191, 1.921295, 1.860718, 
    1.797272, 1.707123, 1.598114, 1.499725, 1.408325, 1.323059, 1.259888, 
    1.212372, 1.169495, 1.174072, 1.369995, 1.57074, 1.68512, 2.585754, 
    4.414459, 4.315063, 4.164917, 5.462891, 5.808533, 5.572388, 5.551941, 
    5.387238, 4.105988, 1.773224, 1.790222, 1.774109, 1.67865, 1.636597, 
    1.559448, 1.544464, 1.537109, 1.613037, 1.821136,
  2.430664, 2.44693, 2.454102, 2.541931, 4.414764, 4.781189, 4.363739, 
    4.105988, 3.979248, 4.557953, 3.573883, 2.44278, 3.522217, 3.210693, 
    2.159821, 2.14267, 2.12207, 2.119141, 2.088867, 2.084229, 2.115692, 
    2.155212, 2.225891, 2.247986, 2.214722, 2.220703, 2.186188, 2.242554, 
    2.347656, 2.440369, 2.43515, 2.421112, 2.630157, 3.904572, 3.156586, 
    2.855865, 2.924042, 2.431122, 2.89389, 2.278076, 2.37027, 2.537933, 
    2.531952, 2.507141, 2.291718, 2.159454, 2.084045, 1.985535, 1.950073, 
    1.944763, 1.919556, 1.914856, 1.918365, 1.985199, 2.036011, 2.120453, 
    2.190887, 2.240753, 2.281982, 2.317505, 2.342133, 2.306, 2.262756, 
    2.146149, 2.075836, 2.031372, 1.944794, 1.884094, 1.790955, 1.710876, 
    1.685333, 1.756195, 1.908966, 1.971313, 2.009186, 2.248444, 4.012054, 
    4.256714, 3.661621, 4.916077, 5.402466, 5.064362, 4.997772, 4.352753, 
    5.013733, 3.675018, 1.837036, 1.87439, 1.849396, 1.855469, 1.897339, 
    1.93573, 1.996155, 2.06778, 2.161194, 2.299683,
  2.551605, 2.524414, 2.477539, 2.515747, 3.967621, 4.434174, 4.382233, 
    4.079926, 4.247162, 4.146667, 3.774078, 2.270844, 2.166077, 2.118347, 
    2.104614, 2.19342, 2.199799, 2.225952, 2.212646, 2.254364, 2.279907, 
    2.331512, 2.300476, 2.300598, 2.281464, 2.329102, 2.372131, 2.436523, 
    2.554413, 2.637939, 2.656921, 2.653198, 2.693481, 2.721466, 2.661072, 
    3.439758, 3.238617, 2.680206, 3.047272, 2.457092, 2.493103, 2.61142, 
    2.532745, 2.43045, 2.307739, 2.229156, 2.146088, 2.130096, 2.125336, 
    2.133728, 2.129944, 2.170898, 2.229248, 2.318298, 2.397339, 2.468658, 
    2.514893, 2.584442, 2.581512, 2.61554, 2.603821, 2.548553, 2.467957, 
    2.38446, 2.353516, 2.280975, 2.216461, 2.199341, 2.160797, 2.165619, 
    2.232605, 2.251617, 2.249481, 2.166931, 2.583588, 3.817719, 3.621277, 
    3.48111, 4.065125, 5.015991, 4.688446, 4.52597, 4.225433, 3.802063, 
    4.192322, 3.032928, 1.930145, 2.022736, 2.06543, 2.137817, 2.175964, 
    2.244385, 2.283386, 2.413818, 2.497589, 2.595642,
  2.55423, 2.644409, 2.639954, 2.547852, 3.604492, 4.010803, 3.613403, 
    3.346375, 3.833466, 4.054901, 3.615875, 2.213074, 2.141968, 2.179016, 
    2.197083, 2.304108, 2.315704, 2.361267, 2.327545, 2.348358, 2.319519, 
    2.317688, 2.273621, 2.31665, 2.312225, 2.399017, 2.445099, 2.469971, 
    2.522217, 2.584381, 2.621155, 2.610291, 2.585724, 2.611328, 2.502594, 
    2.529877, 2.564117, 2.480865, 2.265228, 2.450134, 2.503632, 2.503845, 
    2.435944, 2.368744, 2.307465, 2.217316, 2.141785, 2.141022, 2.110016, 
    2.13559, 2.17981, 2.248566, 2.298492, 2.369934, 2.436249, 2.528564, 
    2.574554, 2.61264, 2.631989, 2.629944, 2.598755, 2.562561, 2.492065, 
    2.482147, 2.423462, 2.379822, 2.37265, 2.362122, 2.352875, 2.372406, 
    2.373199, 2.308136, 2.338867, 2.42981, 2.593048, 2.961761, 3.38736, 
    4.436768, 4.00061, 3.884003, 4.117279, 4.251617, 4.154266, 4.380737, 
    3.748291, 3.42038, 2.840942, 2.145203, 2.289001, 2.331451, 2.357086, 
    2.445526, 2.504059, 2.608704, 2.596497, 2.626038,
  2.733765, 2.846405, 2.783722, 2.789459, 3.757385, 4.12027, 3.417908, 
    3.055786, 3.280792, 3.151581, 3.304871, 2.267975, 2.134888, 2.238281, 
    2.358459, 2.425385, 2.478058, 2.479095, 2.411346, 2.390778, 2.357117, 
    2.329224, 2.317627, 2.381958, 2.417908, 2.548889, 2.536407, 2.573029, 
    2.781128, 2.56424, 2.539459, 2.567444, 2.557953, 2.65451, 2.643555, 
    2.46283, 2.322601, 2.18222, 2.404755, 2.528595, 2.5177, 2.382416, 
    2.283844, 2.234375, 2.11853, 2.057739, 2.00528, 2.006439, 2.050415, 
    2.170807, 2.30127, 2.466644, 2.550262, 2.607635, 2.641388, 2.645203, 
    2.644989, 2.616669, 2.572327, 2.564606, 2.544281, 2.5513, 2.515503, 
    2.503174, 2.454346, 2.463013, 2.447784, 2.458649, 2.4599, 2.440948, 
    2.417908, 2.473389, 2.547638, 2.650787, 2.505127, 3.022186, 4.078064, 
    3.965424, 3.335571, 2.275421, 3.287842, 4.291443, 3.967987, 4.565216, 
    4.068176, 3.475555, 3.319672, 2.304169, 2.467133, 2.544861, 2.60434, 
    2.652344, 2.684357, 2.694489, 2.70343, 2.71936,
  2.848633, 2.928375, 2.816925, 3.110931, 3.827057, 3.50943, 2.739838, 
    2.901367, 3.270844, 2.653656, 3.040283, 3.211792, 2.228271, 2.296417, 
    2.409058, 2.473175, 2.512451, 2.390167, 2.323059, 2.302734, 2.315125, 
    2.341614, 2.354492, 2.426941, 2.50415, 2.590576, 2.55899, 2.939636, 
    2.76947, 2.541595, 2.463745, 2.597534, 2.819061, 2.480347, 2.560333, 
    2.595825, 2.691101, 2.762024, 2.714783, 2.521729, 2.482239, 2.350128, 
    2.223114, 2.146332, 2.053253, 2.036316, 2.068878, 2.173828, 2.419342, 
    2.699615, 2.870453, 2.932373, 2.873688, 2.795959, 2.712311, 2.655273, 
    2.614441, 2.579803, 2.541077, 2.544983, 2.550568, 2.572723, 2.565948, 
    2.541656, 2.533661, 2.537262, 2.558014, 2.598785, 2.548767, 2.548309, 
    2.473755, 2.472717, 2.380157, 2.319, 2.223267, 3.154388, 3.667755, 
    3.378571, 2.87793, 1.386505, 2.162445, 4.401398, 4.544891, 4.222626, 
    3.454773, 2.405365, 2.370575, 2.40332, 2.563416, 2.684265, 2.735168, 
    2.72876, 2.727325, 2.731781, 2.742096, 2.764923,
  2.6698, 2.778259, 2.61615, 2.876831, 3.086456, 2.918823, 2.982086, 
    2.913483, 3.152008, 3.190704, 3.170166, 3.651978, 3.260834, 2.327881, 
    2.458649, 2.581665, 2.611359, 2.476837, 2.310455, 2.223389, 2.188782, 
    2.217377, 2.243927, 2.282684, 2.304108, 2.349884, 2.457031, 3.052002, 
    2.496307, 2.385773, 2.230865, 2.4841, 2.489777, 2.234222, 2.080963, 
    1.879578, 1.804169, 1.996094, 2.298248, 2.420776, 2.377197, 2.255066, 
    2.149811, 2.086914, 2.015991, 2.066864, 2.142456, 2.347046, 2.640442, 
    2.923645, 3.079987, 3.157928, 3.112427, 3.026825, 2.902557, 2.828186, 
    2.74585, 2.691406, 2.637115, 2.614532, 2.640808, 2.653961, 2.605011, 
    2.571564, 2.523834, 2.490875, 2.485229, 2.484222, 2.388794, 2.361908, 
    2.234253, 2.151642, 1.974091, 1.882538, 1.843109, 2.713409, 3.34375, 
    3.008636, 2.645691, 2.487946, 3.263702, 4.748138, 4.863983, 2.445313, 
    2.297333, 2.302216, 2.351868, 2.334686, 2.343414, 2.45105, 2.497131, 
    2.530487, 2.533447, 2.531036, 2.555481, 2.540039,
  2.602905, 2.734253, 2.70813, 2.948822, 2.908783, 2.819489, 2.967834, 
    2.958679, 3.190765, 3.474487, 3.38205, 4.296478, 3.57309, 2.336456, 
    2.374237, 2.52298, 2.653259, 2.767822, 2.608429, 2.47406, 2.230713, 
    2.054138, 2.082031, 2.172394, 2.346283, 2.303253, 2.99527, 2.702148, 
    2.340546, 2.259216, 2.302856, 2.544586, 1.931915, 2.1875, 2.223785, 
    2.045166, 2.055573, 2.20517, 2.379547, 2.421539, 2.344818, 2.235443, 
    2.095459, 1.992401, 1.962311, 2.019745, 1.989288, 1.950165, 2.011566, 
    2.076538, 2.154785, 2.266693, 2.312408, 2.435852, 2.492401, 2.504822, 
    2.459167, 2.50415, 2.545258, 2.565796, 2.555725, 2.536133, 2.441193, 
    2.421082, 2.376678, 2.392303, 2.253448, 2.28653, 2.326172, 2.215515, 
    2.094391, 1.923767, 1.756439, 1.867249, 2.077759, 2.638733, 2.826843, 
    2.774872, 3.37381, 3.425507, 3.584808, 3.3685, 2.780853, 2.355072, 
    2.477539, 2.549805, 2.606842, 2.521088, 2.358521, 2.237823, 2.219849, 
    2.291931, 2.333466, 2.381104, 2.679474, 2.585602,
  2.733215, 2.70639, 2.885345, 3.152924, 3.03476, 3.029999, 3.011993, 
    3.176514, 3.343872, 3.550781, 4.014648, 4.249359, 4.208832, 3.250214, 
    2.527924, 2.51825, 2.591278, 2.583588, 2.528564, 2.411072, 2.3237, 
    2.451447, 2.1539, 2.064667, 2.160339, 2.333221, 2.383545, 2.573883, 
    2.34967, 2.271088, 2.32843, 2.480408, 2.313171, 2.384644, 2.275635, 
    2.244049, 2.326263, 2.321075, 2.329926, 2.245941, 2.227234, 2.20874, 
    2.115906, 2.07782, 2.097626, 2.094666, 2.097382, 2.063263, 2.03894, 
    2.091156, 2.099091, 2.070496, 2.054962, 2.122284, 2.19165, 2.196411, 
    2.155853, 2.218292, 2.288208, 2.362427, 2.337677, 2.353058, 2.379089, 
    2.396942, 2.427399, 2.495026, 2.542725, 2.648987, 2.68573, 2.75351, 
    2.673309, 2.44577, 2.639954, 2.457153, 2.611084, 2.814789, 2.743744, 
    2.997528, 5.210632, 4.244568, 2.356323, 2.364014, 2.421234, 2.408783, 
    2.385803, 2.371033, 2.483459, 2.473694, 2.440369, 2.396393, 2.441986, 
    2.429169, 2.42337, 2.830414, 2.87381, 2.777466,
  2.703644, 2.797119, 3.000366, 3.202209, 3.691986, 4.568207, 4.307739, 
    4.009949, 3.363007, 3.62207, 5.863007, 4.698792, 3.970215, 3.854919, 
    2.758606, 2.641541, 2.677399, 2.516296, 2.500854, 2.391846, 2.695648, 
    2.579559, 2.317322, 2.270508, 2.294403, 2.364075, 2.33606, 2.570313, 
    2.285828, 2.343628, 2.278137, 2.516937, 2.563782, 2.352081, 2.24472, 
    2.28772, 2.329285, 2.268524, 2.216034, 2.16098, 2.150085, 2.155701, 
    2.129822, 2.12384, 2.166718, 2.108215, 2.04657, 2.073578, 2.086334, 
    2.153778, 2.171722, 2.206696, 2.253906, 2.312866, 2.308258, 2.318756, 
    2.334625, 2.382751, 2.408203, 2.444702, 2.427155, 2.486786, 2.45462, 
    2.439606, 2.503204, 2.654694, 2.883972, 3.021484, 2.946655, 2.977509, 
    2.824554, 2.763062, 3.811523, 3.875336, 2.039429, 2.107025, 2.246552, 
    2.236664, 2.329346, 2.344147, 2.275635, 2.269257, 2.207672, 2.195129, 
    2.158905, 2.268127, 2.2966, 2.332855, 2.384308, 2.482056, 2.510223, 
    2.329041, 3.104675, 3.182373, 3.024353, 2.745392,
  3.641174, 4.002167, 4.229401, 4.199707, 4.083862, 4.095428, 3.904205, 
    4.065063, 3.922821, 4.156891, 4.815216, 5.23642, 4.595184, 4.181519, 
    3.693848, 2.534821, 2.595764, 2.516602, 2.443756, 2.340912, 2.59967, 
    2.708344, 2.500702, 2.393494, 2.354279, 2.333649, 2.516235, 2.403107, 
    2.116394, 2.137177, 2.187897, 2.535431, 2.630554, 2.32843, 2.246704, 
    2.354645, 2.255768, 2.166779, 2.148132, 2.067963, 2.061432, 2.122406, 
    2.136963, 2.087769, 2.090424, 2.101318, 2.108459, 2.117584, 2.13092, 
    2.131409, 2.136139, 2.211975, 2.256775, 2.298035, 2.331268, 2.361847, 
    2.389313, 2.460144, 2.465698, 2.49942, 2.576752, 2.603699, 2.501617, 
    2.325348, 2.276154, 2.478699, 2.716187, 2.755035, 2.763184, 2.643829, 
    2.995453, 3.932861, 4.185364, 2.042328, 2.210999, 2.280731, 2.257111, 
    2.240631, 2.180084, 2.208466, 2.174622, 2.120911, 2.103394, 2.118408, 
    2.082794, 2.083832, 2.047058, 2.148773, 2.198975, 2.376831, 2.314453, 
    2.237122, 4.856476, 4.686768, 3.728851, 3.599457,
  4.064209, 3.822235, 3.702942, 3.472687, 3.304504, 2.893494, 2.766907, 
    2.945404, 3.539948, 3.342407, 2.520538, 4.409363, 5.188965, 4.502441, 
    3.939056, 2.061615, 2.21756, 2.40451, 2.4487, 2.341461, 2.520691, 
    2.801819, 2.786438, 2.631317, 2.379944, 2.575073, 2.541931, 2.799133, 
    2.801178, 2.690002, 2.2276, 2.381042, 2.514893, 2.416962, 2.379852, 
    2.357452, 2.290863, 2.202393, 2.101471, 2.054871, 2.073456, 2.117096, 
    2.096924, 2.080658, 2.076172, 2.097473, 2.153503, 2.195251, 2.228821, 
    2.208191, 2.217316, 2.291534, 2.292969, 2.297333, 2.292511, 2.288605, 
    2.28952, 2.31543, 2.34082, 2.370514, 2.443604, 2.454498, 2.318939, 
    2.046753, 1.769989, 1.703705, 2.074219, 2.448059, 2.52948, 2.519653, 
    3.75061, 5.198334, 4.55719, 2.073944, 2.285675, 2.296875, 2.202393, 
    2.197693, 2.169525, 2.137634, 2.11145, 2.132996, 2.103912, 2.078461, 
    2.034821, 2.003662, 1.975769, 1.994141, 1.952209, 2.09433, 2.13855, 
    2.507111, 4.725037, 4.537018, 4.16098, 4.312988,
  4.508484, 4.02829, 3.399292, 2.911133, 2.671936, 2.264252, 2.609894, 
    2.564056, 3.066437, 3.577393, 2.678925, 4.642853, 5.208038, 4.612488, 
    4.350281, 3.190765, 2.23233, 2.195221, 1.299408, 1.851105, 2.482941, 
    2.716919, 2.510284, 2.662048, 2.584442, 2.817963, 3.163147, 2.791412, 
    2.772644, 3.034515, 2.910156, 2.779541, 2.462311, 2.456604, 2.500671, 
    2.483215, 2.394226, 2.263275, 2.19693, 2.178986, 2.180664, 2.195251, 
    2.242249, 2.243744, 2.203247, 2.195007, 2.2276, 2.275146, 2.300659, 
    2.304321, 2.278656, 2.263885, 2.202881, 2.168671, 2.171753, 2.171234, 
    2.145508, 2.123505, 2.132874, 2.150146, 2.219269, 2.276611, 2.231567, 
    1.959961, 1.542358, 1.283661, 1.919861, 4.053131, 3.197662, 2.920441, 
    2.809937, 2.023621, 1.858704, 2.098389, 2.203064, 2.173767, 2.217682, 
    2.208984, 2.247009, 2.224091, 2.227295, 2.242584, 2.190033, 2.225647, 
    2.147858, 2.104248, 2.072388, 2.025787, 2.01004, 1.996796, 1.92157, 
    2.579437, 4.361755, 5.08078, 4.75824, 4.738251,
  4.754608, 4.206024, 3.752533, 3.276398, 2.737061, 2.204956, 2.552368, 
    2.691406, 2.846741, 3.428467, 4.113708, 4.793915, 4.605438, 4.51062, 
    4.729919, 4.415863, 4.122437, 3.456085, 2.435547, 2.094574, 2.313629, 
    2.99942, 3.09967, 3.188751, 3.046783, 2.972504, 3.025757, 2.760254, 
    2.696838, 2.955994, 3.04718, 3.163483, 3.072021, 2.592255, 2.575653, 
    2.567566, 2.5177, 2.44989, 2.399994, 2.338806, 2.300446, 2.294128, 
    2.382813, 2.395691, 2.307159, 2.269409, 2.26004, 2.265686, 2.214691, 
    2.185486, 2.222351, 2.281311, 2.243347, 2.149017, 2.127045, 2.086456, 
    2.069702, 2.057434, 2.012482, 2.055023, 2.07605, 2.086395, 2.093994, 
    1.78717, 1.45462, 1.745941, 4.221954, 4.676819, 3.595459, 2.994476, 
    2.203522, 2.120575, 2.200928, 2.286346, 1.992645, 2.021942, 2.118866, 
    2.215607, 2.342316, 2.305939, 2.262909, 2.286255, 2.248383, 2.239136, 
    2.189301, 2.18573, 2.149048, 2.123169, 2.085419, 1.981384, 1.877289, 
    1.89151, 2.464844, 4.30896, 4.945038, 4.970642,
  5.685486, 5.468079, 4.645599, 3.738129, 3.016205, 2.231384, 2.587341, 
    2.702484, 2.498962, 3.223785, 3.866089, 4.185394, 4.129639, 4.384399, 
    4.5177, 4.482849, 4.188477, 4.024811, 3.979156, 3.807739, 3.605469, 
    3.213531, 3.410034, 3.402405, 3.206726, 2.868256, 2.927399, 3.026733, 
    3.317932, 3.137604, 2.920044, 2.971161, 2.958405, 2.476501, 2.459167, 
    2.52597, 2.541565, 2.490173, 2.429047, 2.394379, 2.440613, 2.37265, 
    2.360413, 2.371674, 2.394989, 2.424866, 2.477295, 2.465698, 2.380005, 
    2.307861, 2.256561, 2.193817, 2.180603, 2.247925, 2.289978, 2.240479, 
    2.171234, 2.118927, 2.024658, 2.043243, 2.01712, 1.989258, 1.966156, 
    1.801941, 1.905792, 3.604401, 4.269043, 3.86554, 3.11145, 2.735748, 
    2.227081, 2.379242, 2.512756, 1.985413, 2.141541, 2.112061, 2.01059, 
    2.008331, 2.163788, 2.250916, 2.37207, 2.372009, 2.252808, 2.164917, 
    2.162445, 2.17395, 2.171875, 2.196564, 2.162018, 2.088959, 2.044159, 
    1.874359, 1.853302, 2.638336, 4.635925, 5.339844,
  6.068298, 5.792053, 5.266876, 3.023376, 2.482086, 2.293152, 2.223511, 
    2.505859, 2.862183, 3.036072, 3.566406, 3.94986, 4.344666, 4.506897, 
    4.438202, 4.428314, 4.067322, 4.143799, 4.421783, 4.565826, 4.17334, 
    4.192169, 4.011139, 3.600922, 3.487366, 3.296539, 3.204315, 3.533783, 
    3.740021, 3.260712, 2.946655, 2.765015, 2.440033, 2.387573, 2.920197, 
    2.622864, 2.910736, 2.934906, 2.402283, 2.325897, 2.320923, 2.341278, 
    2.361603, 2.372009, 2.465057, 2.559174, 2.611664, 2.616486, 2.571594, 
    2.52298, 2.414978, 2.331787, 2.295319, 2.283142, 2.335266, 2.425964, 
    2.360199, 2.279633, 2.217712, 2.139984, 2.066986, 1.937439, 2.048615, 
    2.370331, 3.671875, 4.27005, 4.32547, 3.576294, 3.616516, 3.293762, 
    2.16095, 2.108185, 2.312103, 2.307404, 2.405792, 2.49707, 2.315277, 
    2.120941, 2.045319, 2.178131, 2.240051, 2.191925, 2.260223, 2.221558, 
    2.083984, 1.90506, 1.824829, 2.051178, 2.263092, 2.274536, 2.166473, 
    2.023956, 1.824463, 2.065552, 2.957428, 5.38446,
  4.495239, 2.791595, 2.827667, 2.857025, 2.755524, 2.837708, 3.953705, 
    3.921875, 4.195068, 3.797638, 3.801758, 4.190155, 4.431152, 3.620575, 
    2.635742, 4.177795, 3.865967, 3.468689, 3.970367, 4.549591, 4.250061, 
    4.117889, 4.049255, 3.722229, 3.765869, 3.750793, 3.581055, 3.910431, 
    3.683716, 3.322418, 3.185394, 2.982819, 2.919556, 3.067078, 3.103485, 
    2.840302, 2.733521, 2.597473, 2.34903, 2.314209, 2.39212, 2.537689, 
    2.662109, 2.705658, 2.77655, 2.850006, 2.819, 2.753448, 2.694733, 
    2.591614, 2.474548, 2.42865, 2.426117, 2.320435, 2.227539, 2.222717, 
    2.273895, 2.34375, 2.325256, 2.242004, 2.160767, 1.974976, 2.225861, 
    3.36908, 4.357971, 4.550934, 4.976135, 4.741974, 3.960114, 3.542328, 
    2.842834, 2.561523, 2.553711, 2.511841, 2.597198, 2.746857, 2.858276, 
    2.912262, 2.619385, 2.424408, 2.255707, 2.379669, 2.577148, 2.42038, 
    2.098175, 1.669464, 1.251617, 1.278717, 1.728851, 2.087494, 2.233826, 
    2.102142, 1.876831, 2.106445, 4.033997, 4.966553,
  3.755951, 2.720245, 2.969849, 3.501709, 2.996765, 3.62439, 3.826019, 
    3.380157, 3.097137, 3.164337, 3.466003, 3.808624, 3.616699, 2.564331, 
    3.310699, 3.773438, 3.72168, 3.473175, 3.704102, 4.128113, 4.164551, 
    4.25882, 4.110107, 3.974182, 4.035309, 4.147614, 3.951904, 3.970978, 
    3.922821, 3.853302, 3.856812, 3.376068, 3.096313, 2.989807, 2.873535, 
    2.72049, 2.650879, 2.634613, 2.619354, 2.967163, 2.786041, 2.737091, 
    2.703735, 2.662537, 2.646057, 2.683624, 2.642761, 2.559784, 2.526215, 
    2.489563, 2.443115, 2.387268, 2.319641, 2.228882, 2.119629, 2.024689, 
    2.100433, 2.191284, 2.181091, 2.242218, 2.268921, 2.058258, 2.25296, 
    3.406708, 3.827057, 4.396912, 4.434601, 4.614807, 3.789886, 2.969391, 
    2.843628, 3.049805, 2.942749, 2.824158, 3.199738, 3.254852, 3.420807, 
    3.524567, 3.440155, 3.267853, 2.954712, 2.757263, 2.670746, 2.326965, 
    2.021271, 1.632233, 1.08197, 0.8517456, 1.100769, 1.482117, 1.910156, 
    2.048096, 1.892578, 2.0961, 3.580658, 4.020172,
  2.804535, 2.790527, 2.878113, 3.022949, 3.136444, 2.863647, 2.589355, 
    2.832886, 2.966827, 3.016174, 2.831329, 2.95108, 2.988434, 3.10199, 
    2.46106, 3.044708, 3.154449, 3.403473, 3.797546, 3.77475, 3.770477, 
    3.942993, 4.086151, 3.903564, 3.840149, 3.836639, 3.799988, 3.808807, 
    3.891846, 3.710968, 3.734009, 3.614594, 3.484863, 3.292236, 2.868317, 
    2.742737, 2.851349, 2.706207, 2.773071, 2.832306, 2.493317, 2.472504, 
    2.442352, 2.385834, 2.381897, 2.421326, 2.416138, 2.367096, 2.365082, 
    2.395599, 2.397034, 2.32373, 2.223602, 2.161316, 2.107391, 2.04184, 
    2.046326, 2.093018, 2.107147, 2.210388, 2.217529, 2.049774, 2.194183, 
    3.07901, 3.465546, 3.636292, 3.521423, 3.868652, 3.584595, 3.558105, 
    3.518982, 2.997559, 3.053558, 3.338684, 3.303223, 3.347107, 3.493195, 
    3.614746, 3.624817, 3.642944, 3.20047, 2.704987, 1.936737, 1.703674, 
    1.728607, 1.699585, 1.265503, 0.8856506, 0.8256836, 0.9135132, 1.290192, 
    1.766296, 1.869568, 1.874664, 2.170013, 2.881287,
  2.325806, 2.464264, 2.43454, 2.42453, 2.241364, 2.258148, 2.134918, 
    2.530762, 2.496124, 2.426147, 2.306091, 2.396118, 2.56012, 2.507538, 
    2.550354, 2.691528, 2.824982, 3.074829, 3.226654, 3.241241, 3.324585, 
    3.370605, 3.493744, 3.586731, 3.338196, 3.328369, 3.04715, 3.121002, 
    3.05072, 3.069977, 3.157349, 3.049561, 2.995117, 2.91925, 2.748779, 
    2.643555, 2.696289, 2.629944, 2.055969, 2.221191, 2.558838, 2.695923, 
    2.6073, 2.47934, 2.446716, 2.455322, 2.467804, 2.49704, 2.516693, 
    2.48114, 2.41272, 2.367157, 2.364014, 2.395752, 2.37381, 2.286438, 
    2.231415, 2.226654, 2.224121, 2.201721, 2.147491, 2.176666, 2.542542, 
    2.764862, 2.835632, 2.951965, 3.306305, 3.660004, 3.576538, 3.64444, 
    3.565308, 3.410645, 3.415466, 3.486816, 3.447174, 3.446381, 3.460602, 
    3.393982, 3.378998, 3.417084, 3.194916, 3.081543, 2.172058, 2.06424, 
    1.88623, 1.569427, 0.9880066, 0.2859192, -0.004730225, 0.1812744, 
    0.6516418, 1.194672, 1.553558, 1.698608, 1.84198, 2.016632,
  2.027649, 1.863647, 2.106415, 2.025757, 2.081024, 2.094543, 2.063965, 
    1.912537, 1.761749, 1.606262, 1.620422, 1.823517, 2.116699, 2.166626, 
    2.2966, 2.371796, 2.741119, 2.872345, 2.951538, 3.118774, 3.208313, 
    3.187012, 3.354858, 3.230713, 3.210205, 3.142273, 2.93042, 2.960205, 
    3.065552, 3.153259, 3.033539, 2.939728, 2.747253, 2.545135, 2.482361, 
    2.608398, 2.677917, 2.556854, 1.956573, 2.108612, 2.591827, 2.884613, 
    2.76828, 2.459076, 2.393524, 2.521515, 2.523132, 2.51236, 2.499939, 
    2.480164, 2.470337, 2.54306, 2.662903, 2.718719, 2.644043, 2.475342, 
    2.368988, 2.352905, 2.320129, 2.254517, 2.124939, 2.394379, 2.572601, 
    2.724091, 2.819885, 2.92337, 3.00415, 3.118896, 3.101715, 3.235199, 
    3.464294, 3.342621, 3.378204, 3.288574, 3.365906, 3.909363, 3.494202, 
    3.412231, 3.323334, 3.106689, 2.798553, 2.091217, 1.858063, 1.506531, 
    1.246399, 1.213898, 0.9726257, 0.4069824, -0.02218628, 0.06121826, 
    0.5098572, 0.9974365, 1.326324, 1.517334, 1.813202, 1.891937,
  1.309692, 1.556519, 1.385834, 1.789154, 1.814087, 2.036621, 1.862335, 
    1.869446, 1.802002, 1.697601, 1.609497, 1.720581, 1.926697, 2.163544, 
    2.340363, 2.504242, 2.697906, 2.686188, 2.819305, 2.799652, 2.909332, 
    3.164673, 3.229126, 3.157166, 3.043884, 2.930511, 2.820892, 2.712128, 
    2.835724, 2.98349, 3.167511, 3.107269, 2.798431, 2.556, 2.478638, 
    2.49527, 2.520172, 2.563995, 2.036407, 2.037567, 2.169281, 2.179291, 
    2.615295, 2.510681, 2.063416, 2.432892, 2.741119, 2.785645, 2.855103, 
    2.942871, 3.02536, 3.034027, 2.956543, 2.862793, 2.383026, 2.338776, 
    2.265961, 2.30368, 2.30188, 2.200348, 2.431274, 2.550049, 2.735687, 
    2.846069, 2.883972, 3.115601, 3.319611, 3.116791, 3.148865, 3.279236, 
    3.348816, 3.293823, 3.008209, 3.005554, 3.248566, 3.58847, 3.334961, 
    3.156708, 2.954376, 2.630005, 1.754944, 1.469788, 1.140533, 0.8253174, 
    0.8823547, 1.028046, 1.140564, 1.052429, 0.7834167, 0.7212524, 0.8999634, 
    1.13031, 1.259277, 1.278351, 1.375244, 1.656219,
  1.051605, 1.327881, 1.575836, 1.64621, 1.682037, 1.548584, 1.820526, 
    1.904114, 1.960602, 1.987244, 2.089142, 2.290222, 2.52652, 2.768097, 
    3.031647, 3.102814, 3.039154, 3.043121, 2.98996, 3.022675, 3.036896, 
    2.993835, 2.934357, 3.017456, 3.023376, 3.09198, 2.90741, 2.900055, 
    2.943542, 2.958862, 2.901123, 2.850311, 2.66391, 2.423187, 2.187622, 
    2.196503, 2.317596, 2.61145, 2.384247, 2.40567, 2.349945, 2.637695, 
    2.760284, 2.705933, 2.532349, 2.582947, 2.468079, 2.148499, 2.531036, 
    2.917908, 3.074158, 2.955658, 2.416016, 2.235046, 2.084839, 1.965759, 
    2.051056, 2.161133, 2.229767, 2.269226, 2.36972, 2.568481, 2.752808, 
    2.758728, 2.784882, 2.958771, 3.116577, 3.142639, 3.029724, 2.941681, 
    2.852844, 2.489899, 2.486481, 2.506531, 2.573792, 2.514923, 2.693115, 
    2.721252, 2.236511, 1.824097, 1.385101, 1.036591, 0.798645, 0.6626892, 
    1.105194, 0.4723816, 0.8201599, 1.11026, 1.268066, 1.334656, 1.288849, 
    1.118011, 0.8603821, 0.6860962, 0.8553772, 0.991333,
  0.4713135, 0.4273376, 0.5844727, 1.118622, 1.294098, 1.443359, 1.272095, 
    1.67807, 1.869263, 2.05423, 2.263611, 2.453003, 2.634949, 2.880005, 
    3.079437, 3.215363, 3.310883, 3.351868, 3.32724, 3.279968, 3.116425, 
    2.945251, 2.779419, 2.696411, 2.74588, 3.111115, 3.285553, 3.278137, 
    3.029053, 2.73761, 2.70697, 2.578583, 2.387115, 2.273499, 2.175079, 
    2.283264, 2.857483, 3.335632, 3.162109, 3.217468, 2.825195, 2.831787, 
    2.910797, 2.963593, 2.805084, 2.691925, 2.444, 2.382996, 2.44516, 
    2.272034, 2.373901, 2.486664, 2.182922, 2.102386, 2.088409, 2.095764, 
    2.307922, 2.626892, 2.629761, 2.574066, 2.620758, 2.611969, 2.573914, 
    2.612549, 2.637787, 2.642639, 2.699097, 2.720184, 2.757446, 2.7789, 
    2.789795, 2.892303, 3.082184, 3.090912, 2.351257, 1.971771, 1.808075, 
    2.536194, 2.582764, 2.148102, 1.227936, 1.066803, 1.682678, 2.272766, 
    2.25351, 1.807251, 1.486694, 0.7793579, 0.7599487, 0.8678894, 0.8617249, 
    1.028534, 0.6893616, 0.4220581, 0.3667908, 0.3504333,
  0.7781677, 0.7185059, 0.6593323, 0.589325, 0.3761292, 1.144135, 1.289703, 
    1.519318, 1.77774, 1.930939, 2.01236, 1.766327, 1.866486, 2.00827, 
    2.712769, 2.875244, 2.990997, 3.11087, 3.026825, 2.91217, 2.852997, 
    2.78183, 2.761963, 2.734039, 2.867706, 3.468628, 3.709778, 3.435669, 
    3.00528, 2.796722, 2.711731, 2.659515, 2.68042, 2.796539, 3.01828, 
    3.357941, 2.936981, 3.14505, 2.898956, 2.848877, 2.800507, 2.682556, 
    2.474152, 2.447632, 2.430084, 2.494141, 2.567383, 2.779419, 3.039368, 
    3.302795, 2.866394, 2.640381, 2.615112, 2.427612, 2.463165, 2.56424, 
    2.736969, 2.748169, 2.910797, 2.623444, 2.572144, 2.481201, 2.471039, 
    2.556335, 2.679352, 2.749542, 2.727539, 2.640045, 2.519714, 1.953339, 
    2.286591, 2.749664, 2.899536, 1.591919, 2.428558, 2.405792, 2.884705, 
    2.849396, 2.744843, 1.411682, 1.25, 1.212311, 2.468689, 3.155365, 
    3.180237, 3.080475, 2.889313, 2.597015, 2.211395, 2.088226, 1.387299, 
    1.220856, 0.9737549, 0.890625, 0.873291, 0.8786316,
  1.442139, 1.259186, 1.097046, 0.9261169, 0.7790833, 0.9567261, 1.39682, 
    1.793091, 1.999878, 1.988617, 1.873962, 1.810883, 1.838928, 1.949677, 
    1.975311, 3.135559, 3.171722, 3.248505, 3.163727, 3.171997, 2.859528, 
    2.642914, 2.596222, 2.521881, 2.646942, 2.703735, 2.886597, 3.089508, 
    2.939667, 2.796936, 2.883789, 2.985199, 3.003784, 3.056458, 3.01001, 
    2.240967, 2.092438, 2.067383, 2.749756, 2.969971, 3.33902, 3.473877, 
    3.4328, 3.692444, 4.009308, 4.297333, 4.591797, 4.841675, 5.157074, 
    5.129364, 5.110931, 4.824463, 4.519928, 4.323151, 4.208008, 4.123138, 
    4.107758, 4.126648, 4.050476, 3.857819, 3.630249, 3.552124, 3.458099, 
    3.571411, 3.601715, 3.628723, 3.560547, 3.451569, 3.216431, 1.944092, 
    2.851044, 3.07196, 1.666077, 3.894928, 4.288757, 4.660095, 4.713623, 
    4.323456, 3.021484, 1.929443, 1.675781, 2.765991, 3.858795, 3.642868, 
    3.748627, 3.303635, 3.064987, 3.140945, 3.00032, 3.140472, 3.93985, 
    2.545258, 2.05957, 1.697998, 1.537262, 1.517822,
  1.785522, 1.524414, 1.557739, 1.709686, 1.759033, 1.92337, 2.218811, 
    2.45932, 2.516907, 2.553314, 2.631653, 2.864777, 3.122009, 3.525238, 
    3.957367, 4.428253, 4.580414, 4.535614, 4.315613, 4.038483, 3.551636, 
    3.093964, 2.693939, 2.393372, 2.345062, 3.036591, 3.286591, 3.636139, 
    3.821594, 4.115875, 4.221558, 4.450073, 4.60318, 4.342377, 4.322784, 
    4.37619, 4.348938, 4.481171, 4.667389, 4.758118, 4.859436, 4.912048, 
    4.965027, 5.091614, 5.263672, 5.418152, 5.647736, 5.907867, 6.099213, 
    6.238159, 6.157227, 6.018494, 5.86673, 5.689789, 5.639954, 5.63855, 
    5.69043, 5.827881, 5.931427, 6.032745, 6.176239, 6.264252, 6.452911, 
    6.683777, 7.157684, 5.960541, 5.960297, 5.802948, 5.613464, 5.430939, 
    5.220367, 5.351746, 5.47937, 5.888367, 6.144012, 6.691132, 6.76947, 
    5.23407, 5.138489, 4.832214, 4.521606, 4.37027, 4.183792, 3.864716, 
    3.436005, 3.005936, 3.00769, 3.284897, 3.378784, 3.67363, 4.12207, 
    5.10907, 5.689789, 4.319275, 3.040436, 2.127594,
  5.286987, 5.1138, 4.739838, 4.41217, 4.524414, 4.680206, 4.818115, 
    5.572327, 5.630554, 5.620728, 5.683929, 5.695221, 5.844604, 5.8284, 
    5.773438, 5.634308, 5.185364, 4.796082, 4.553772, 4.36908, 4.239777, 
    4.171814, 4.021088, 3.868744, 3.683594, 4.489563, 4.585297, 4.781067, 
    5.001892, 5.208588, 5.231964, 5.32312, 5.374481, 5.329346, 5.308136, 
    5.307953, 5.31955, 5.402679, 5.496735, 5.568207, 5.625641, 5.683472, 
    5.743835, 5.780396, 5.862823, 5.948242, 6.073547, 6.184113, 6.255341, 
    6.313721, 6.363342, 6.380615, 6.315948, 6.200867, 6.130981, 6.069397, 
    6.0737, 6.141144, 6.258911, 6.338104, 6.398102, 6.450378, 6.572205, 
    6.716919, 6.807159, 6.855682, 6.773285, 6.758453, 6.745819, 6.735413, 
    6.677551, 7.052795, 6.222473, 6.060104, 5.783279, 5.457825, 5.239319, 
    5.083588, 4.943085, 4.728058, 4.510147, 4.362503, 4.214706, 4.007492, 
    3.787567, 3.675323, 3.641998, 3.77507, 4.116211, 4.524353, 4.926605, 
    5.264618, 7.260223, 6.871277, 6.151642, 5.706329,
  7.044586, 6.638977, 6.409576, 6.18457, 6.053833, 5.856384, 5.646332, 
    5.619934, 5.653595, 5.647644, 5.688538, 5.722351, 5.753082, 5.780975, 
    5.785553, 5.785919, 5.74823, 5.746155, 5.731262, 5.703979, 5.667297, 
    5.671326, 5.64856, 5.64505, 5.634705, 5.688416, 5.624023, 5.607758, 
    5.624023, 5.597931, 5.501526, 5.389526, 5.280518, 5.226166, 5.174042, 
    5.149689, 5.151947, 5.158661, 5.167969, 5.22818, 5.275269, 5.315277, 
    5.33374, 5.355591, 5.408386, 5.459198, 5.488953, 5.539734, 5.619202, 
    5.722198, 5.794342, 5.855682, 5.900726, 5.888031, 5.916473, 5.919037, 
    5.993866, 6.076447, 6.177734, 6.329834, 6.509766, 6.672058, 6.851318, 
    7.051758, 7.249481, 7.394592, 7.53894, 7.667145, 7.800201, 7.954224, 
    8.104279, 8.286987, 8.394409, 8.456512, 8.479889, 8.47525, 8.487701, 
    8.568314, 8.702454, 8.816422, 9.0634, 9.177292, 9.267319, 9.251938, 
    9.3517, 9.437744, 9.659561, 9.733185, 9.83519, 9.600937, 9.317566, 
    8.822723, 8.545105, 8.288788, 7.875458, 7.472809,
  6.62619, 6.458008, 6.395111, 6.334167, 6.25766, 6.166687, 6.080994, 
    5.984955, 5.927917, 5.899994, 5.841858, 5.786865, 5.756195, 5.768036, 
    5.748322, 5.74469, 5.75885, 5.783905, 5.818726, 5.82193, 5.817139, 
    5.799652, 5.813416, 5.819794, 5.812347, 5.79129, 5.774658, 5.762634, 
    5.752075, 5.727234, 5.683594, 5.635284, 5.554565, 5.524231, 5.497192, 
    5.458496, 5.421295, 5.378143, 5.335449, 5.306793, 5.290314, 5.243591, 
    5.241608, 5.226044, 5.238892, 5.266418, 5.253601, 5.220642, 5.244141, 
    5.288635, 5.347046, 5.401306, 5.463806, 5.544159, 5.625519, 5.739014, 
    5.861298, 5.952545, 6.103973, 6.217346, 6.330811, 6.470673, 6.602295, 
    6.737854, 6.891296, 7.036346, 7.188568, 7.345001, 7.486206, 7.609711, 
    7.744232, 7.832886, 7.914032, 8.034332, 8.18634, 8.279419, 8.386719, 
    8.46579, 8.489746, 8.483093, 8.502594, 8.472168, 8.421692, 8.338898, 
    8.246979, 8.207581, 8.141785, 8.048584, 7.950806, 7.81665, 7.671051, 
    7.541748, 7.405792, 7.246765, 7.030609, 6.836517,
  1.59787, 1.598251, 1.600082, 1.602631, 1.60672, 1.614136, 1.624039, 
    1.638229, 1.659134, 1.680878, 1.706604, 1.731125, 1.757034, 1.781921, 
    1.796967, 1.802231, 1.796494, 1.779587, 1.755417, 1.718964, 1.675079, 
    1.623062, 1.564529, 1.508408, 1.454697, 1.409073, 1.375275, 1.350021, 
    1.331329, 1.318695, 1.308685, 1.302429, 1.299362, 1.300079, 1.308151, 
    1.316422, 1.330093, 1.348846, 1.370331, 1.392654, 1.417267, 1.441803, 
    1.468445, 1.494034, 1.521957, 1.547729, 1.570206, 1.597351, 1.623138, 
    1.64624, 1.663956, 1.682251, 1.689285, 1.688309, 1.687775, 1.698837, 
    1.718048, 1.715973, 1.652237, 1.667007, 1.66127, 1.668106, 1.652176, 
    1.658936, 1.658279, 1.653076, 1.653854, 1.651962, 1.651199, 1.659012, 
    1.658997, 1.660889, 1.663559, 1.724884, 1.635941, 1.596176, 1.599762, 
    1.625534, 1.522095, 1.502625, 1.493576, 1.485031, 1.482635, 1.487839, 
    1.500671, 1.508163, 1.515198, 1.524826, 1.537643, 1.549698, 1.563171, 
    1.572998, 1.581924, 1.58992, 1.59436, 1.598129,
  1.749619, 1.689148, 1.616943, 1.544998, 1.48172, 1.439392, 1.398056, 
    1.355881, 1.319229, 1.297409, 1.285889, 1.28569, 1.307053, 1.351181, 
    1.416229, 1.498001, 1.60054, 1.715118, 1.805359, 1.853333, 1.842407, 
    1.796768, 1.713303, 1.626251, 1.546951, 1.493637, 1.462585, 1.45842, 
    1.474243, 1.490784, 1.500854, 1.510757, 1.52092, 1.536026, 1.55899, 
    1.591614, 1.636795, 1.6987, 1.778931, 1.871765, 1.969482, 2.087128, 
    2.213501, 2.323273, 2.427048, 2.564285, 2.629654, 2.720795, 2.817215, 
    2.921509, 3.004654, 3.00563, 3.069962, 3.038513, 3.285904, 2.958755, 
    2.945023, 2.950424, 2.943512, 2.939407, 2.934021, 2.934799, 2.942459, 
    2.951706, 2.964081, 2.942398, 2.917068, 2.883987, 2.922211, 2.927826, 
    2.84436, 2.762833, 2.668243, 2.57164, 2.48381, 2.322144, 2.200012, 
    2.09903, 2.058029, 2.022995, 1.873062, 1.874496, 1.717468, 1.718643, 
    1.590378, 1.562576, 1.609009, 1.641876, 1.688629, 1.74025, 1.785492, 
    1.824097, 1.853729, 1.853455, 1.840775, 1.805023,
  1.444153, 1.409073, 1.394089, 1.435242, 1.440186, 1.46434, 1.588303, 
    1.831985, 2.127609, 2.376511, 2.485825, 2.476059, 2.410507, 2.33139, 
    2.276306, 2.244217, 2.19455, 2.152496, 2.150665, 2.190445, 2.288437, 
    2.417145, 2.503403, 2.43718, 2.235367, 2.04129, 1.90126, 1.860031, 
    1.859329, 1.84404, 1.809601, 1.758682, 1.727951, 1.728012, 1.74968, 
    1.771301, 1.819931, 1.883682, 1.96994, 2.077621, 2.215057, 2.443649, 
    2.679779, 3.081085, 3.507507, 3.845337, 3.962906, 3.9935, 4.008286, 
    4.023071, 4.047287, 4.019745, 3.95401, 3.87738, 3.882965, 3.914825, 
    3.85994, 3.706421, 3.528748, 3.32634, 3.179977, 3.129196, 3.163971, 
    3.177307, 3.140701, 3.139862, 3.134781, 3.128479, 3.038361, 2.907761, 
    2.752884, 2.625153, 2.480042, 2.314072, 2.157715, 2.069244, 2.019363, 
    1.961823, 1.86911, 1.782913, 1.709274, 1.671844, 1.678482, 1.670212, 
    1.603363, 1.543518, 1.582397, 1.621445, 1.702759, 1.769165, 1.855576, 
    1.893921, 1.876266, 1.789017, 1.666885, 1.535629,
  1.893372, 2.050934, 2.253922, 2.429306, 2.546631, 2.568054, 2.545532, 
    2.470261, 2.352173, 2.246307, 2.173401, 2.181915, 2.300797, 2.450806, 
    2.599228, 2.729889, 2.835358, 2.911667, 2.937973, 2.740051, 2.424698, 
    2.152756, 1.954636, 1.901184, 2.079315, 2.350861, 2.496948, 2.505356, 
    2.492264, 2.554962, 2.622284, 2.652374, 2.655411, 2.609726, 2.507828, 
    2.37001, 2.335495, 2.334656, 2.304626, 2.249176, 2.226837, 2.24826, 
    2.325943, 2.515854, 2.973267, 3.636627, 2.204269, 2.444626, 2.456207, 
    2.631668, 2.789215, 2.939163, 3.05336, 3.166763, 3.33812, 3.560379, 
    3.748993, 3.697296, 3.615982, 3.392532, 3.265198, 3.153748, 3.138184, 
    3.043381, 2.92366, 2.890594, 2.874252, 2.793655, 2.652832, 2.580566, 
    2.594833, 2.618332, 2.64418, 2.667557, 2.619232, 2.532837, 2.468582, 
    2.435394, 2.431808, 2.317612, 2.247223, 2.19072, 2.286179, 2.327957, 
    2.393524, 2.346588, 2.298859, 2.254974, 2.212723, 1.811111, 1.823669, 
    1.85466, 1.777771, 1.768692, 1.757446, 1.802689,
  1.682709, 1.628937, 1.614471, 1.674362, 1.759262, 1.759323, 1.746048, 
    1.753342, 1.886795, 1.918182, 1.999573, 2.015961, 2.023514, 2.13269, 
    2.374557, 2.394943, 2.157883, 2.024353, 2.092346, 2.254761, 2.13179, 
    1.988434, 1.93927, 1.996704, 2.241562, 2.412766, 2.325989, 2.302628, 
    2.383469, 2.593185, 2.873657, 3.033142, 3.073975, 3.035187, 2.984787, 
    2.942856, 2.900543, 2.937195, 2.876511, 2.735306, 2.567993, 2.379181, 
    2.334473, 2.446976, 2.72789, 3.12796, 2.319107, 2.459671, 2.506348, 
    2.487915, 2.469299, 2.348267, 2.322952, 2.379135, 2.537857, 2.702637, 
    2.763184, 2.674179, 2.54776, 2.432648, 2.294174, 2.127243, 2.115982, 
    2.220993, 2.397232, 2.538895, 2.698257, 2.803268, 2.864273, 2.832916, 
    3.520599, 3.101074, 3.184143, 3.149109, 3.130066, 3.038116, 3.490387, 
    3.33226, 3.130432, 2.985001, 2.719162, 2.574646, 2.588898, 2.52243, 
    2.578552, 2.682785, 2.732651, 2.823792, 2.797363, 2.594238, 2.263962, 
    2.015259, 1.736954, 1.617538, 1.720337, 1.757523,
  2.06871, 1.795395, 2.008362, 1.871063, 1.802704, 1.81279, 1.867935, 
    2.07373, 2.165192, 2.215469, 2.233826, 2.133041, 1.972092, 1.914734, 
    1.948151, 1.918381, 1.769501, 1.698151, 1.77919, 2.029068, 2.161682, 
    1.986023, 1.740067, 1.678162, 1.757126, 1.745789, 1.762283, 1.75856, 
    1.786163, 1.831879, 1.889679, 1.959671, 2.029968, 2.040527, 2.03421, 
    2.015518, 1.911942, 1.808365, 1.748795, 1.744629, 1.793015, 1.882004, 
    1.945084, 1.997238, 1.875809, 1.890732, 1.830688, 1.781937, 1.690521, 
    1.593643, 1.499893, 1.444992, 1.414673, 1.411804, 1.533081, 1.764862, 
    2.04599, 2.275208, 2.436279, 2.513885, 2.500397, 2.581146, 2.634583, 
    2.708557, 2.827026, 2.96167, 3.153198, 3.327881, 3.485962, 3.576202, 
    3.645782, 3.901184, 4.086975, 4.107574, 4.108795, 3.948059, 3.750153, 
    3.62912, 3.912842, 3.771515, 3.450165, 3.381912, 3.319031, 3.212311, 
    3.112396, 3.065704, 3.097412, 3.138947, 3.097549, 2.997345, 2.893951, 
    2.787842, 2.742599, 2.583923, 2.455704, 2.340607,
  2.592529, 2.571899, 2.637115, 2.53653, 2.531662, 2.502563, 2.526382, 
    2.542267, 2.557358, 2.612061, 2.757782, 2.752548, 2.802872, 2.829163, 
    2.76358, 2.664734, 2.443634, 2.378021, 2.489853, 2.681, 2.782242, 
    2.740173, 2.584717, 2.329773, 2.041153, 1.917984, 1.860428, 1.705505, 
    1.456268, 1.138184, 0.9685059, 0.9178772, 0.9830933, 1.956299, 2.283234, 
    2.475876, 2.212662, 2.134827, 2.077423, 2.130676, 2.21701, 2.173767, 
    2.118713, 1.996613, 1.834778, 1.59845, 1.440369, 1.245056, 0.7352905, 
    0.2807007, -0.07406616, -0.1816101, -0.1374207, -0.1192017, 0.2745056, 
    0.6603088, 1.038483, 1.323883, 1.59436, 1.832123, 2.133179, 2.375732, 
    2.553619, 2.707642, 2.863281, 2.947144, 3.07782, 3.298248, 3.366669, 
    3.832031, 4.021759, 4.392853, 4.573395, 4.804565, 4.747345, 4.692657, 
    4.513123, 4.287781, 4.01825, 3.923065, 3.858093, 3.839355, 3.857574, 
    3.881927, 3.86734, 3.770325, 3.670197, 3.602875, 3.446686, 3.267334, 
    3.224304, 3.181335, 3.07666, 2.925476, 2.823853, 2.729523,
  3.017456, 2.971252, 2.839417, 2.778198, 2.817474, 2.885742, 2.918488, 
    2.921478, 2.872437, 2.934906, 3.009247, 3.13147, 3.306976, 3.311737, 
    3.3927, 3.200348, 3.187042, 3.30072, 3.212708, 3.287659, 3.315002, 
    3.303619, 3.187653, 2.868134, 2.468201, 2.035156, 1.677368, 1.390594, 
    1.089264, 0.7659912, 0.3903809, 0.1237793, 0.4679871, 0.7475586, 
    1.191315, 1.950623, 2.318176, 2.351501, 2.186554, 2.065979, 1.868988, 
    1.85495, 1.814728, 1.870667, 1.846039, 1.755096, 1.702759, 1.393768, 
    0.4472961, -0.3634644, -0.7579956, -0.9232788, -1.015198, -1.017761, 
    -0.7554016, -0.4820862, -0.2898254, -0.06164551, 0.06750488, 0.4587402, 
    0.9060669, 1.444794, 1.894501, 2.24942, 2.622162, 2.987976, 3.082062, 
    3.368835, 3.704163, 3.926239, 3.96402, 3.901306, 4.051697, 4.085358, 
    4.270447, 4.303558, 4.1539, 3.878662, 3.652649, 3.175659, 3.045929, 
    3.402771, 3.732391, 3.779755, 3.684479, 3.603424, 3.563416, 3.582611, 
    3.493469, 3.4534, 3.51413, 3.556854, 3.476837, 3.3013, 3.117279, 3.046753,
  3.04541, 2.977234, 2.802368, 2.769104, 3.053467, 3.092194, 2.931732, 
    2.851379, 2.77652, 2.82782, 2.656403, 2.752991, 2.93042, 2.934998, 
    3.410065, 3.905823, 4.108429, 4.225281, 4.404633, 4.852295, 4.81369, 
    4.636017, 4.279175, 3.790894, 3.031616, 2.298004, 1.820526, 1.393463, 
    1.277161, 1.131989, 1.043457, 0.9512024, 0.8751831, 0.7142944, 0.6469421, 
    0.7671204, 1.185333, 1.509186, 1.611389, 1.587433, 1.706207, 2.040619, 
    2.4245, 2.532898, 2.329559, 2.145264, 1.914856, 1.621613, 0.9135437, 
    0.06530762, -0.2121277, -0.1954956, -0.1954346, -0.3062439, -0.4839172, 
    -0.5982361, -0.7149048, -0.7088623, -0.3013916, 0.1882019, 0.6443481, 
    1.010468, 1.260803, 1.57428, 1.832947, 2.089722, 2.248322, 2.403717, 
    2.522308, 2.64682, 2.719421, 2.697632, 2.683716, 2.686981, 2.632813, 
    2.352448, 1.895905, 1.754608, 1.764648, 1.759949, 1.741486, 1.762634, 
    1.718964, 1.710022, 1.890259, 2.246368, 2.714386, 3.016632, 3.123566, 
    3.1875, 3.273315, 3.369019, 3.49411, 3.394012, 3.20874, 3.038574,
  2.242798, 2.199554, 2.406708, 2.615814, 2.509247, 2.535492, 2.589661, 
    2.570496, 2.641602, 2.604889, 2.479095, 2.43985, 2.446869, 2.51651, 
    2.714569, 2.899353, 3.095947, 3.292725, 3.322266, 2.912415, 2.661896, 
    2.513885, 2.345093, 2.339661, 2.179169, 1.939697, 1.96817, 2.056976, 
    2.087616, 2.044922, 1.84552, 1.557617, 1.301636, 1.142853, 1.130402, 
    1.284485, 1.576172, 1.887299, 2.019531, 1.972382, 2.003967, 2.204163, 
    2.417236, 2.295288, 1.983734, 1.911987, 1.959381, 1.941528, 1.607361, 
    1.090179, 0.8540344, 0.7464294, 0.6383362, 0.4926147, 0.3400269, 
    0.2185669, 0.1871948, 0.2687378, 0.4443359, 0.6441345, 0.8370972, 
    0.9916077, 1.114014, 1.230011, 1.31427, 1.398773, 1.529297, 1.691711, 
    1.804932, 1.890564, 1.97702, 1.991028, 1.96582, 1.906708, 1.668945, 
    1.275452, 1.389709, 2.595703, 2.758118, 1.705231, 1.499634, 1.455231, 
    1.602356, 1.510284, 1.310028, 1.413818, 1.746796, 2.028046, 2.303497, 
    2.3078, 2.42215, 2.613464, 2.664581, 2.64859, 2.518829, 2.321564,
  2.121674, 2.253845, 2.356628, 2.389709, 2.4198, 2.436523, 2.513916, 
    2.614014, 2.699615, 2.772919, 2.845245, 2.948334, 3.009766, 3.019653, 
    3.025391, 3.075134, 3.225128, 3.523834, 3.681519, 3.469147, 3.145111, 
    3.005005, 2.869934, 2.661438, 2.477997, 2.43631, 2.466339, 2.462952, 
    2.477539, 2.463928, 2.307343, 1.979034, 1.637878, 1.483856, 1.535736, 
    1.648773, 1.709778, 1.703003, 1.65686, 1.736023, 2.014923, 2.296906, 
    2.344391, 2.144714, 2.144501, 2.194366, 2.16925, 2.117188, 1.953644, 
    1.709564, 1.431641, 1.207275, 1.135223, 1.11792, 1.03775, 0.9483337, 
    0.9266357, 0.9880981, 1.106323, 1.204742, 1.231262, 1.235535, 1.241119, 
    1.269318, 1.313416, 1.339111, 1.365234, 1.41922, 1.448425, 1.455536, 
    1.455475, 1.436462, 1.36615, 1.239197, 1.067261, 1.130005, 1.855865, 
    2.255524, 1.936523, 1.700439, 1.441223, 1.378967, 1.519073, 1.565948, 
    1.502655, 1.597046, 1.763672, 1.972595, 2.156647, 2.289764, 2.315643, 
    2.268036, 2.225189, 2.189667, 2.153961, 2.093048,
  2.098053, 2.259308, 2.407745, 2.511108, 2.570038, 2.674683, 2.901154, 
    3.13443, 3.24173, 3.351044, 3.539459, 3.630981, 3.629425, 3.577209, 
    3.469147, 3.297852, 3.189789, 3.300842, 3.484711, 3.664124, 4.020996, 
    4.256012, 3.97113, 3.438354, 3.075623, 2.853882, 2.649231, 2.46405, 
    2.345428, 2.21814, 1.991699, 1.740387, 1.616699, 1.611877, 1.614685, 
    1.564026, 1.440338, 1.299652, 1.226868, 1.406921, 1.927826, 2.313324, 
    2.425293, 2.317627, 2.555634, 2.588959, 2.429138, 2.312286, 2.223663, 
    2.114014, 1.970154, 1.850708, 1.773712, 1.709747, 1.608307, 1.53595, 
    1.516449, 1.515015, 1.509155, 1.497375, 1.505219, 1.46814, 1.387939, 
    1.322418, 1.291168, 1.24527, 1.220856, 1.215973, 1.209015, 1.167419, 
    1.127014, 1.13913, 1.144928, 1.117798, 1.079193, 1.145416, 1.632111, 
    1.948364, 1.823792, 1.54715, 1.388214, 1.350769, 1.524292, 1.557922, 
    1.444, 1.414001, 1.473236, 1.652466, 1.83432, 1.893799, 1.904694, 
    1.937653, 1.947144, 1.898254, 1.879028, 1.953979,
  2.341248, 2.431488, 2.52182, 2.539795, 2.539917, 2.852509, 3.505096, 
    3.99646, 4.175354, 4.329834, 4.521606, 4.456604, 4.065216, 3.727905, 
    3.505676, 3.27536, 3.118652, 3.090332, 3.187683, 3.331085, 3.44516, 
    3.326324, 2.906311, 2.432526, 2.159027, 2.026459, 1.916626, 1.788361, 
    1.679657, 1.598206, 1.537842, 1.544769, 1.504303, 1.340851, 1.129913, 
    1.063873, 1.141571, 1.246368, 1.454651, 1.668579, 2.114624, 2.500427, 
    2.593109, 2.494171, 2.694824, 2.874573, 2.817749, 2.554718, 2.555878, 
    2.614441, 2.698212, 2.569183, 2.355103, 2.08844, 1.881592, 1.793213, 
    1.717377, 1.6026, 1.52771, 1.51001, 1.503235, 1.464996, 1.368408, 
    1.340454, 1.332062, 1.286041, 1.27594, 1.247711, 1.231476, 1.265961, 
    1.285889, 1.314026, 1.346191, 1.303101, 1.191711, 1.074951, 1.237518, 
    1.632019, 1.771881, 1.554779, 1.399658, 1.309082, 1.500885, 1.701843, 
    1.69281, 1.635773, 1.634277, 1.732971, 1.888885, 1.943848, 1.887543, 
    1.903809, 1.928802, 1.940765, 2.051666, 2.213531,
  2.247559, 2.179657, 2.110565, 2.123749, 2.39801, 2.991516, 3.28537, 
    3.511505, 3.722321, 3.544434, 3.083252, 2.701874, 2.392487, 2.180054, 
    2.061676, 2.037659, 2.004028, 1.944885, 1.940582, 1.86795, 1.743988, 
    1.59198, 1.374176, 1.215271, 1.128296, 1.133087, 1.17688, 1.179321, 
    1.319763, 1.718384, 1.968842, 1.776031, 1.466919, 1.080902, 0.9270325, 
    1.213837, 1.528595, 1.619446, 1.821869, 2.155487, 2.207062, 2.73468, 
    2.993011, 2.781921, 2.743286, 2.831543, 2.778748, 2.650238, 2.575287, 
    2.375397, 2.147186, 1.995667, 1.921509, 1.776276, 1.664948, 1.623718, 
    1.559601, 1.482269, 1.4758, 1.516907, 1.525818, 1.499054, 1.480103, 
    1.520538, 1.537476, 1.513458, 1.521393, 1.48114, 1.504272, 1.558167, 
    1.532898, 1.544128, 1.503235, 1.409393, 1.30777, 1.145752, 1.251068, 
    1.808594, 1.893951, 1.699646, 1.441101, 1.506622, 1.95459, 2.184875, 
    2.149963, 2.068481, 2.004211, 1.954834, 1.983795, 1.941376, 1.910797, 
    1.936249, 2.003693, 2.11734, 2.180176, 2.230499,
  1.850861, 1.799316, 1.830231, 1.994568, 2.334015, 2.459015, 2.404205, 
    2.498657, 2.922272, 2.416473, 1.643707, 1.474335, 1.556274, 1.565735, 
    1.418549, 1.319946, 1.303558, 1.256683, 1.167023, 0.991333, 0.8661194, 
    0.8416138, 0.8722229, 1.003357, 1.111298, 1.23233, 1.437714, 1.709656, 
    2.180634, 2.419617, 1.775299, 1.722229, 1.663849, 1.525513, 1.597015, 
    1.70639, 1.743469, 2.067993, 2.298553, 2.185516, 1.674255, 2.884064, 
    3.474548, 3.212219, 2.995026, 2.985168, 2.801056, 2.457062, 2.08429, 
    1.540771, 1.246155, 1.259644, 1.324707, 1.366241, 1.414734, 1.484192, 
    1.536804, 1.559601, 1.603088, 1.672546, 1.698364, 1.685974, 1.680634, 
    1.721039, 1.737854, 1.723938, 1.718597, 1.687988, 1.648346, 1.626282, 
    1.561035, 1.508759, 1.398285, 1.30896, 1.262268, 1.103638, 1.221313, 
    2.747284, 2.384552, 1.564819, 1.363159, 1.587158, 2.179413, 2.690521, 
    2.191742, 1.966064, 1.981598, 1.969696, 1.886627, 1.77124, 1.782318, 
    1.856934, 1.857666, 1.876923, 1.873077, 1.865845,
  1.738892, 1.675507, 1.690643, 1.762756, 1.871979, 2.823486, 3.609894, 
    4.025543, 3.329895, 2.231964, 2.035217, 2.129639, 2.095001, 2.020416, 
    1.911316, 1.816284, 1.81842, 1.76416, 1.66983, 1.685242, 1.828552, 
    1.939209, 2.01416, 2.089935, 2.158356, 2.228027, 2.397369, 2.517029, 
    2.46286, 1.943329, 1.786804, 3.705933, 3.011536, 2.453888, 2.601105, 
    2.578918, 2.742462, 2.5513, 2.294647, 1.980316, 1.274658, 2.129883, 
    2.150635, 2.30246, 2.513641, 2.581909, 2.288452, 1.701263, 1.38382, 
    1.246063, 1.24942, 1.440796, 1.5784, 1.630371, 1.66272, 1.691162, 
    1.704926, 1.714996, 1.667145, 1.683868, 1.685242, 1.686493, 1.681946, 
    1.688049, 1.702362, 1.675995, 1.591431, 1.506592, 1.43338, 1.382843, 
    1.310059, 1.253204, 1.202759, 1.176483, 1.13974, 1.001343, 1.214661, 
    2.432831, 2.844116, 2.15686, 1.805359, 2.150146, 2.140137, 2.222198, 
    2.040802, 1.854095, 1.847961, 1.797394, 1.883392, 1.926483, 1.842682, 
    1.827576, 1.76709, 1.790466, 1.764801, 1.747803,
  1.563202, 1.551331, 1.656433, 1.800873, 2.158173, 3.284698, 4.588135, 
    4.425568, 3.199402, 2.334839, 2.215485, 2.427429, 2.495117, 2.302277, 
    2.501373, 2.527405, 2.553986, 2.529694, 2.436188, 2.471497, 2.425507, 
    2.442963, 2.429993, 2.401031, 2.394745, 2.292328, 2.225159, 2.059357, 
    1.921814, 1.821167, 1.983398, 3.954742, 3.87973, 3.177734, 3.128723, 
    2.765411, 2.914856, 3.03653, 2.824982, 2.494324, 1.429749, 1.520752, 
    1.392761, 1.548828, 1.805145, 1.883087, 1.861328, 1.873779, 1.876038, 
    1.901703, 1.930328, 1.917053, 1.856079, 1.770966, 1.674988, 1.586914, 
    1.536591, 1.471344, 1.449951, 1.48172, 1.470581, 1.429291, 1.38327, 
    1.36496, 1.402405, 1.352081, 1.321808, 1.291656, 1.25058, 1.229156, 
    1.176605, 1.184662, 1.16684, 1.091766, 0.9390869, 1.047302, 1.614624, 
    2.897156, 3.894806, 2.691254, 2.117462, 2.616394, 2.639069, 2.710938, 
    2.351471, 1.903717, 1.869781, 1.955017, 1.938202, 1.868408, 1.835541, 
    1.817993, 1.812042, 1.751892, 1.623627, 1.562256,
  1.645569, 1.808319, 2.014526, 2.319, 3.32785, 3.884644, 4.588989, 4.111786, 
    3.637573, 3.845184, 2.396759, 2.559753, 4.14447, 2.429688, 2.314117, 
    2.480011, 2.350403, 2.343048, 2.231323, 2.213165, 2.170227, 2.149872, 
    2.142181, 2.105347, 2.085144, 2.017517, 1.994019, 1.922668, 1.932526, 
    2.021942, 2.172516, 3.984833, 4.181915, 3.802795, 3.73822, 3.092712, 
    2.863678, 2.918549, 2.914856, 2.3284, 1.434753, 1.632538, 1.782288, 
    1.961212, 2.027649, 2.050049, 2.04837, 2.093292, 2.032227, 1.925903, 
    1.844421, 1.725983, 1.627472, 1.471924, 1.364502, 1.348022, 1.325958, 
    1.307953, 1.344788, 1.343903, 1.335236, 1.372986, 1.397461, 1.430664, 
    1.463196, 1.391083, 1.334961, 1.312622, 1.288544, 1.206787, 1.199524, 
    1.215942, 1.091827, 1.014587, 1.069305, 1.497955, 2.387573, 3.971741, 
    4.459808, 3.129791, 2.740814, 3.497406, 3.956848, 4.086639, 4.090302, 
    2.296997, 1.806091, 1.860138, 1.824982, 1.718933, 1.682281, 1.607544, 
    1.532684, 1.501617, 1.473724, 1.532745,
  2.008148, 2.178009, 2.307373, 2.464111, 3.838348, 4.637939, 4.390106, 
    4.228516, 4.419525, 4.416901, 2.471893, 2.462891, 3.961639, 3.390839, 
    2.138733, 2.178406, 2.083649, 2.082764, 2.062622, 2.05545, 2.083405, 
    2.092041, 2.169281, 2.194397, 2.188477, 2.133942, 2.084045, 2.057831, 
    2.139069, 2.273071, 2.368622, 2.680389, 3.978333, 3.922913, 3.564728, 
    3.188782, 3.060028, 3.116364, 2.775726, 1.967987, 1.825653, 2.057709, 
    2.229309, 2.26413, 2.198761, 2.165741, 2.095367, 2.036469, 1.962952, 
    1.881104, 1.826263, 1.689789, 1.592834, 1.518036, 1.497528, 1.540833, 
    1.555084, 1.59668, 1.699982, 1.761505, 1.83905, 1.878174, 1.868561, 
    1.847656, 1.768829, 1.65506, 1.577026, 1.49881, 1.414459, 1.372894, 
    1.339478, 1.334839, 1.35202, 1.535614, 1.623566, 1.683502, 2.628693, 
    4.357941, 4.020264, 3.685089, 3.463593, 4.102844, 4.667969, 5.418884, 
    5.808655, 4.863983, 1.858215, 1.812866, 1.816284, 1.681183, 1.641296, 
    1.589172, 1.601349, 1.595581, 1.671051, 1.853455,
  2.358215, 2.375519, 2.418427, 2.418121, 4.132629, 4.976379, 4.249176, 
    4.066101, 4.140869, 4.451172, 3.736633, 2.433441, 3.154816, 3.303589, 
    2.097015, 2.070435, 2.09082, 2.107819, 2.160156, 2.22876, 2.288544, 
    2.314819, 2.335999, 2.312836, 2.272186, 2.304291, 2.289856, 2.375916, 
    2.47345, 2.550079, 2.57547, 2.600067, 2.913422, 3.855225, 3.514038, 
    3.4729, 3.381256, 2.427429, 2.810364, 2.087158, 2.244019, 2.403473, 
    2.394806, 2.372314, 2.235809, 2.171417, 2.11203, 2.087555, 2.05658, 
    2.025116, 1.962372, 1.878906, 1.848755, 1.909241, 1.957733, 2.034637, 
    2.123322, 2.192108, 2.294159, 2.353516, 2.388336, 2.349548, 2.282867, 
    2.2099, 2.134644, 2.070831, 1.975037, 1.927734, 1.851196, 1.836182, 
    1.843231, 1.917511, 2.008026, 2.028503, 2.048309, 2.236084, 3.919922, 
    4.177307, 3.831207, 4.404022, 3.944061, 3.958252, 4.464783, 4.562683, 
    6.308716, 4.961731, 1.811981, 1.894989, 1.870636, 1.839325, 1.922729, 
    1.915497, 2.038483, 2.108398, 2.217529, 2.30838,
  2.490021, 2.473511, 2.52948, 2.539398, 3.912689, 4.91394, 4.033325, 
    3.712891, 4.258911, 4.203522, 3.654541, 2.201508, 2.09726, 2.095764, 
    2.085114, 2.182373, 2.225861, 2.263275, 2.30545, 2.366608, 2.385529, 
    2.37915, 2.372528, 2.381897, 2.422272, 2.453247, 2.477661, 2.568115, 
    2.622131, 2.66217, 2.69101, 2.686584, 2.770966, 2.762238, 2.66864, 
    3.448578, 3.189636, 2.503754, 2.765839, 2.33429, 2.387939, 2.443024, 
    2.421021, 2.377014, 2.296295, 2.254272, 2.241852, 2.251495, 2.220093, 
    2.182953, 2.131989, 2.157745, 2.223633, 2.313416, 2.391418, 2.464325, 
    2.531372, 2.609558, 2.642517, 2.618408, 2.5737, 2.49585, 2.423431, 
    2.363861, 2.306122, 2.266022, 2.192902, 2.178986, 2.175964, 2.212372, 
    2.269684, 2.2724, 2.31723, 2.317261, 2.728973, 3.878113, 3.942047, 
    3.597046, 3.823517, 3.851288, 3.502197, 3.901703, 4.14975, 4.2966, 
    5.63559, 4.176697, 1.965881, 2.045441, 2.113922, 2.141663, 2.180511, 
    2.21817, 2.299042, 2.393097, 2.468811, 2.527863,
  2.556122, 2.598236, 2.68515, 2.496307, 4.039276, 4.761383, 3.109833, 
    2.847443, 3.361115, 3.640686, 3.116455, 2.175262, 2.200073, 2.194275, 
    2.279877, 2.354584, 2.316925, 2.385132, 2.370392, 2.373047, 2.359131, 
    2.356659, 2.382111, 2.415405, 2.448639, 2.518555, 2.568298, 2.577606, 
    2.525543, 2.563416, 2.568512, 2.577942, 2.568817, 2.601685, 2.551575, 
    2.530457, 2.524353, 2.522064, 2.546082, 2.341858, 2.372406, 2.364777, 
    2.38562, 2.357025, 2.299103, 2.255981, 2.22049, 2.187561, 2.136719, 
    2.15625, 2.184631, 2.269409, 2.352478, 2.443573, 2.510193, 2.597717, 
    2.62851, 2.649353, 2.660156, 2.62735, 2.584381, 2.535065, 2.485138, 
    2.438721, 2.404633, 2.378723, 2.365295, 2.356049, 2.36322, 2.40683, 
    2.41803, 2.398132, 2.503784, 2.619446, 2.715027, 3.439911, 3.614868, 
    3.898041, 3.399475, 3.294861, 2.969788, 3.054169, 3.51355, 4.567444, 
    4.262573, 4.210236, 3.62912, 2.21402, 2.40564, 2.419342, 2.406097, 
    2.492981, 2.523743, 2.581757, 2.572968, 2.575592,
  2.732544, 2.804443, 2.782959, 2.658325, 4.162354, 4.562439, 2.939056, 
    2.808533, 2.898773, 2.700104, 3.343628, 2.237427, 2.178925, 2.2948, 
    2.428772, 2.466919, 2.475983, 2.442657, 2.425659, 2.416992, 2.408844, 
    2.423126, 2.412323, 2.477081, 2.545715, 2.675385, 2.733063, 2.709625, 
    2.658478, 2.567902, 2.532623, 2.561676, 2.563019, 2.593414, 2.626434, 
    2.488739, 2.312622, 2.335236, 2.438538, 2.58139, 2.421875, 2.284454, 
    2.231659, 2.228302, 2.163696, 2.108765, 2.088593, 2.161194, 2.291809, 
    2.400391, 2.544403, 2.629822, 2.692596, 2.725067, 2.763855, 2.772461, 
    2.737885, 2.721039, 2.709869, 2.693481, 2.647339, 2.628326, 2.604126, 
    2.56543, 2.572906, 2.572052, 2.567505, 2.549225, 2.548553, 2.567078, 
    2.579498, 2.644623, 2.7052, 2.776245, 2.589386, 3.053436, 3.632477, 
    2.876617, 3.513062, 3.138428, 2.769135, 2.826813, 3.408905, 4.313141, 
    3.94278, 3.8284, 3.879883, 2.420319, 2.637115, 2.598907, 2.602936, 
    2.623901, 2.637695, 2.661591, 2.671875, 2.69455,
  2.790192, 2.848236, 2.7211, 3.067963, 3.588531, 3.297577, 2.901154, 
    2.912292, 2.757446, 2.004486, 3.140472, 3.194916, 2.295563, 2.351044, 
    2.449524, 2.396332, 2.363037, 2.279816, 2.31665, 2.334381, 2.364136, 
    2.413483, 2.414246, 2.492035, 2.596405, 2.736176, 2.701263, 2.504547, 
    2.476868, 2.561584, 2.455139, 2.65976, 2.661987, 2.382721, 2.51059, 
    2.648254, 2.63266, 2.594391, 2.68985, 2.421143, 2.39682, 2.29718, 
    2.175629, 2.09967, 2.107605, 2.176239, 2.357422, 2.65918, 2.977539, 
    3.103577, 3.156708, 3.133118, 3.096802, 3.079468, 3.094421, 3.093292, 
    3.074219, 3.046692, 3.037231, 3.014069, 2.937378, 2.85611, 2.823761, 
    2.810272, 2.842651, 2.824493, 2.790741, 2.758118, 2.699554, 2.67038, 
    2.593689, 2.578064, 2.439331, 2.338348, 2.235931, 3.004608, 3.432617, 
    3.101898, 3.461456, 3.267334, 2.955994, 3.87085, 3.805267, 3.614777, 
    3.244598, 2.46344, 2.504181, 2.517914, 2.651428, 2.663849, 2.709503, 
    2.680511, 2.723389, 2.738678, 2.732178, 2.748688,
  2.531006, 2.700348, 2.585724, 3.015533, 3.172852, 3.091278, 3.291992, 
    3.24585, 2.790802, 2.700073, 2.687897, 3.798035, 3.577759, 2.394897, 
    2.451477, 2.54422, 2.518738, 2.364166, 2.292969, 2.256836, 2.222992, 
    2.281708, 2.262024, 2.278259, 2.320984, 2.453857, 2.561188, 2.518616, 
    2.397797, 2.394745, 2.479095, 2.573975, 2.486328, 2.232422, 2.142456, 
    1.946503, 1.818939, 2.016907, 2.298065, 2.376099, 2.343933, 2.272186, 
    2.149811, 2.088806, 2.147064, 2.316864, 2.590057, 2.943176, 3.269073, 
    3.461639, 3.544342, 3.535828, 3.478058, 3.443939, 3.420044, 3.38327, 
    3.334442, 3.244873, 3.177399, 3.097839, 3.036194, 2.944855, 2.881531, 
    2.844147, 2.782745, 2.728699, 2.654694, 2.621948, 2.543945, 2.477844, 
    2.357025, 2.21991, 2.026489, 1.888458, 1.835083, 2.793304, 3.658325, 
    3.348511, 3.266602, 3.448059, 3.679291, 4.1474, 4.106262, 2.358734, 
    2.380585, 2.311615, 2.37381, 2.389648, 2.414246, 2.4375, 2.479645, 
    2.468933, 2.492432, 2.503967, 2.509369, 2.441193,
  2.816162, 2.788727, 2.866119, 3.138916, 3.194397, 3.227386, 3.278168, 
    3.1763, 3.050598, 3.081757, 2.985199, 3.278961, 3.570648, 2.424561, 
    2.377075, 2.532349, 2.671448, 2.731445, 2.621155, 2.556, 2.404388, 
    2.320313, 2.28595, 2.27124, 2.356262, 2.31543, 2.976776, 2.735046, 
    2.375732, 2.26239, 2.309845, 2.654999, 2.036072, 2.255341, 2.295044, 
    2.125397, 2.10437, 2.217072, 2.364929, 2.423431, 2.391876, 2.332489, 
    2.190826, 2.066925, 2.048767, 2.0495, 2.092316, 2.136139, 2.297424, 
    2.481262, 2.60025, 2.682312, 2.733551, 2.827789, 2.856964, 2.829102, 
    2.777008, 2.715179, 2.69635, 2.677948, 2.649628, 2.55481, 2.469391, 
    2.448029, 2.377533, 2.428986, 2.342316, 2.362488, 2.450134, 2.447723, 
    2.376556, 2.181946, 2.029694, 2.016998, 2.075378, 2.81601, 3.05014, 
    3.056122, 3.66745, 4.187225, 3.496307, 3.172791, 2.666779, 2.360474, 
    2.437134, 2.478455, 2.495361, 2.478394, 2.459839, 2.327148, 2.320313, 
    2.330383, 2.334625, 2.350464, 2.700775, 2.810944,
  3.027344, 2.931183, 3.154572, 3.580933, 3.718384, 3.471741, 3.381256, 
    3.358795, 3.382935, 3.222839, 3.269226, 3.471436, 3.333069, 2.814575, 
    2.444977, 2.470886, 2.656586, 2.595123, 2.502014, 2.412506, 2.336151, 
    2.468109, 2.424225, 2.233063, 2.298828, 2.304688, 2.324219, 2.782867, 
    2.345398, 2.262573, 2.279297, 2.380859, 2.363007, 2.459198, 2.283661, 
    2.293549, 2.367126, 2.312775, 2.329224, 2.2453, 2.257172, 2.25351, 
    2.211975, 2.170166, 2.165924, 2.186066, 2.160736, 2.073303, 2.109436, 
    2.204041, 2.215546, 2.166718, 2.154175, 2.187958, 2.202789, 2.231964, 
    2.180206, 2.168488, 2.224945, 2.346527, 2.368958, 2.352203, 2.397186, 
    2.447388, 2.465759, 2.551575, 2.627289, 2.720947, 2.741547, 2.78775, 
    2.76004, 2.612579, 2.706726, 2.597137, 2.983337, 3.058594, 2.91275, 
    3.362518, 5.156067, 4.487, 2.342957, 2.388, 2.420441, 2.342041, 2.337311, 
    2.351929, 2.437347, 2.54538, 2.555847, 2.492249, 2.514191, 2.433838, 
    2.474915, 2.849457, 2.963867, 2.993958,
  3.22937, 3.364319, 3.367706, 3.671692, 4.34491, 4.627289, 4.928253, 
    4.541199, 3.631714, 4.515564, 4.554688, 4.580139, 3.568939, 3.221405, 
    2.568542, 2.559265, 2.623688, 2.466614, 2.437897, 2.317261, 2.650848, 
    2.786987, 2.42807, 2.387177, 2.3526, 2.244202, 2.153503, 2.754181, 
    2.549652, 2.548828, 2.283386, 2.461395, 2.507996, 2.486786, 2.233398, 
    2.269196, 2.294861, 2.249725, 2.217834, 2.171814, 2.185944, 2.205933, 
    2.187134, 2.187683, 2.202972, 2.189453, 2.160919, 2.192383, 2.281128, 
    2.330872, 2.360229, 2.339447, 2.329559, 2.355927, 2.355469, 2.376251, 
    2.376495, 2.396606, 2.423248, 2.475739, 2.443604, 2.461304, 2.453064, 
    2.484894, 2.557037, 2.695496, 2.931366, 3.055603, 2.935272, 2.923218, 
    2.789703, 2.800049, 3.269012, 3.054932, 2.169922, 2.176056, 2.178711, 
    2.187164, 2.240692, 2.287567, 2.228851, 2.273254, 2.243347, 2.228638, 
    2.14563, 2.248566, 2.262177, 2.349548, 2.384369, 2.522034, 2.517517, 
    2.363922, 3.994202, 4.227814, 4.043732, 3.216217,
  3.598053, 3.749939, 3.74942, 3.766663, 3.744904, 3.561523, 3.517059, 
    3.391296, 3.237762, 3.718292, 4.299194, 4.69928, 3.952728, 3.917236, 
    3.379761, 2.458527, 2.530975, 2.393372, 2.310425, 2.228119, 3.029877, 
    3.284576, 2.497131, 2.497009, 2.315491, 2.196167, 2.898102, 3.240936, 
    2.68869, 2.164673, 2.270569, 2.579437, 2.636902, 2.345123, 2.282623, 
    2.290649, 2.227081, 2.151703, 2.112762, 2.071136, 2.126495, 2.179169, 
    2.176422, 2.134552, 2.164642, 2.204102, 2.216675, 2.243805, 2.289581, 
    2.283722, 2.266235, 2.302673, 2.316162, 2.353241, 2.377106, 2.379608, 
    2.443298, 2.494659, 2.505737, 2.519409, 2.532867, 2.498169, 2.410736, 
    2.355774, 2.391998, 2.623566, 2.788544, 2.756378, 2.757416, 3.116211, 
    3.258087, 3.65033, 3.617462, 2.1427, 2.263733, 2.29303, 2.246399, 
    2.237305, 2.171204, 2.239014, 2.199432, 2.156128, 2.145599, 2.123871, 
    2.071625, 2.105133, 2.081177, 2.206512, 2.23703, 2.384766, 2.302277, 
    2.305542, 4.351379, 4.440735, 4.049408, 3.450531,
  3.539398, 3.500458, 3.393219, 3.401642, 3.324371, 3.133453, 3.062439, 
    3.102997, 3.26004, 2.936768, 2.525757, 4.437805, 4.552002, 4.68338, 
    4.115173, 2.718231, 2.252319, 2.283936, 2.337891, 2.269318, 3.261566, 
    3.393646, 2.949463, 2.819183, 2.322083, 2.582886, 2.792511, 2.992584, 
    3.113281, 2.617188, 2.312195, 2.411133, 2.541656, 2.493225, 2.425568, 
    2.391266, 2.284821, 2.166931, 2.072662, 2.079895, 2.154755, 2.190826, 
    2.183197, 2.175323, 2.173615, 2.203796, 2.264526, 2.300842, 2.335236, 
    2.33609, 2.333405, 2.369995, 2.370575, 2.327423, 2.294556, 2.251648, 
    2.299805, 2.357544, 2.415497, 2.453827, 2.508667, 2.444, 2.268951, 
    2.037567, 1.922211, 2.075317, 2.383057, 2.624542, 3.164459, 3.201355, 
    4.036316, 4.259308, 3.568359, 2.117188, 2.284119, 2.304993, 2.201172, 
    2.233276, 2.208588, 2.176422, 2.119049, 2.130157, 2.113037, 2.0914, 
    2.039459, 2.010742, 1.998566, 2.029236, 1.96637, 2.064362, 2.091736, 
    2.450317, 4.29129, 4.231842, 3.871338, 3.830231,
  4.033722, 3.84082, 3.426514, 3.036652, 2.970123, 2.704498, 2.933807, 
    2.967712, 3.332764, 3.370911, 2.719727, 4.402679, 4.762085, 4.933411, 
    4.610107, 3.786499, 2.292969, 2.35611, 2.298981, 2.390625, 2.82428, 
    3.216492, 2.96347, 3.078125, 2.763336, 2.840485, 2.560822, 2.633636, 
    2.877655, 2.965729, 3.196106, 2.661224, 2.382111, 2.489258, 2.46521, 
    2.445831, 2.383667, 2.279297, 2.164581, 2.163483, 2.211517, 2.206757, 
    2.230621, 2.21524, 2.239655, 2.275452, 2.313324, 2.363434, 2.384888, 
    2.428711, 2.407166, 2.359711, 2.303314, 2.231506, 2.207489, 2.171814, 
    2.119202, 2.124817, 2.187408, 2.192963, 2.263, 2.275177, 2.179108, 
    1.925598, 1.655121, 1.624695, 2.190033, 3.920898, 3.857483, 3.469177, 
    3.453064, 2.234192, 1.941864, 2.162628, 2.258453, 2.215424, 2.19162, 
    2.224091, 2.256439, 2.28418, 2.263611, 2.240967, 2.222321, 2.23111, 
    2.178772, 2.164734, 2.131836, 2.058411, 2.029938, 1.985352, 1.863007, 
    2.354828, 4.120392, 4.441345, 4.184967, 4.133911,
  4.317719, 3.998566, 3.480225, 3.37677, 3.167358, 2.732819, 3.065704, 
    2.950714, 3.029633, 3.645721, 3.895782, 4.718658, 4.896698, 5.00592, 
    4.654236, 4.197144, 4.102478, 3.740417, 3.459686, 2.742523, 2.505859, 
    3.090881, 3.603333, 3.347412, 2.865845, 3.012024, 2.981079, 2.785858, 
    2.757782, 2.663239, 2.683624, 2.581421, 2.622009, 2.463135, 2.443939, 
    2.49231, 2.48645, 2.451233, 2.34433, 2.257233, 2.221619, 2.255463, 
    2.342712, 2.37735, 2.353638, 2.337311, 2.314087, 2.337311, 2.331818, 
    2.357422, 2.411713, 2.437897, 2.424866, 2.301086, 2.21817, 2.127808, 
    2.050446, 2.037323, 2.040253, 2.093506, 2.091064, 2.051239, 1.980865, 
    1.807953, 1.622467, 1.89505, 3.716125, 4.325714, 4.408447, 4.512421, 
    3.864258, 2.480072, 2.447998, 2.49054, 2.480072, 2.1297, 2.168945, 
    2.229431, 2.294189, 2.304626, 2.305878, 2.324524, 2.315552, 2.302979, 
    2.283081, 2.300262, 2.239014, 2.220703, 2.158417, 2.008606, 1.860352, 
    1.88327, 2.386505, 3.875519, 4.131836, 4.230103,
  4.56427, 4.479431, 4.228455, 3.537506, 3.183289, 2.2789, 2.970062, 
    2.933899, 2.40152, 3.389984, 4.090668, 4.456055, 4.595001, 4.55481, 
    4.719452, 4.387085, 4.270782, 4.068573, 4.023254, 3.720642, 3.707184, 
    3.286133, 3.965546, 3.477478, 2.823425, 2.871613, 2.974823, 3.324341, 
    3.469238, 3.003052, 2.421112, 2.35791, 2.652954, 2.341522, 2.390869, 
    2.532043, 2.591095, 2.546021, 2.470825, 2.368561, 2.28894, 2.229736, 
    2.278503, 2.30307, 2.331635, 2.407684, 2.469604, 2.486084, 2.487549, 
    2.510681, 2.524689, 2.520447, 2.511414, 2.497925, 2.451538, 2.327515, 
    2.172028, 2.063141, 1.943878, 1.952148, 1.960114, 1.94989, 1.921753, 
    1.832367, 1.946014, 3.167206, 3.709381, 3.77301, 4.307312, 4.678589, 
    4.408264, 4.047516, 4.039978, 3.527069, 3.070831, 2.242249, 2.107819, 
    2.071747, 2.173981, 2.250763, 2.385742, 2.392242, 2.33606, 2.284698, 
    2.286591, 2.257813, 2.223236, 2.272919, 2.236938, 2.144287, 2.06015, 
    1.838013, 1.912567, 2.495514, 4.117035, 4.492401,
  4.52594, 4.667542, 4.741913, 2.98645, 2.581909, 2.351868, 2.092133, 
    2.24173, 2.57077, 2.874207, 3.919708, 3.934631, 3.984741, 4.027588, 
    3.809326, 3.748871, 3.722382, 3.876404, 4.180298, 4.039154, 3.453491, 
    3.746887, 3.874756, 3.573639, 3.157654, 2.609283, 2.811188, 3.879669, 
    4.431335, 3.735565, 2.828369, 2.738007, 2.656555, 2.358276, 3.143585, 
    2.505249, 3.040863, 3.095612, 2.516663, 2.455597, 2.315643, 2.220947, 
    2.244659, 2.256165, 2.27832, 2.376556, 2.473755, 2.526428, 2.561462, 
    2.610168, 2.623871, 2.640411, 2.627106, 2.5513, 2.486115, 2.416077, 
    2.263733, 2.125671, 2.040039, 2.007416, 1.974487, 1.919525, 1.981506, 
    2.061584, 2.557953, 3.07901, 3.545807, 3.640869, 3.927246, 4.203278, 
    4.068481, 4.04245, 4.012695, 3.354797, 3.23349, 3.300079, 2.474792, 
    2.260681, 2.156128, 2.209167, 2.312439, 2.250061, 2.292297, 2.296478, 
    2.203583, 2.080017, 1.939911, 2.05481, 2.246552, 2.308014, 2.225281, 
    2.036652, 1.859375, 2.015228, 2.662048, 4.046631,
  3.737549, 2.847961, 2.81427, 2.738037, 2.700134, 2.600189, 2.913116, 
    3.489288, 3.903229, 3.76059, 3.607269, 3.47052, 3.276215, 2.853882, 
    2.216156, 2.79834, 2.792755, 3.017944, 3.581268, 3.614563, 3.654358, 
    3.772919, 3.688232, 3.094269, 3.573181, 3.362488, 2.845459, 3.085999, 
    3.5513, 3.429626, 2.748627, 2.602783, 2.569733, 2.730011, 2.798767, 
    2.602448, 2.628937, 2.92157, 2.540649, 2.522064, 2.462555, 2.459442, 
    2.522064, 2.566925, 2.588165, 2.590546, 2.598816, 2.62677, 2.652283, 
    2.636627, 2.60791, 2.639893, 2.664337, 2.585266, 2.478455, 2.356262, 
    2.239777, 2.161072, 2.083862, 1.993408, 1.906647, 1.881592, 2.005676, 
    2.050568, 2.178162, 2.617615, 3.072479, 3.312256, 3.417877, 3.466095, 
    3.718506, 3.678802, 3.730316, 3.61792, 3.421631, 3.475891, 3.541382, 
    3.043243, 2.713287, 2.495239, 2.342377, 2.360291, 2.523285, 2.421692, 
    2.175842, 1.898865, 1.523773, 1.427551, 1.735596, 2.045837, 2.220642, 
    2.134369, 1.941223, 2.01413, 3.056152, 3.957001,
  3.184937, 2.786194, 2.918121, 3.259064, 2.861572, 2.716766, 2.509338, 
    2.847992, 2.963318, 2.77536, 3.024475, 2.795319, 2.625366, 2.27121, 
    2.64743, 2.753296, 2.531677, 2.567871, 2.828491, 3.153778, 3.093048, 
    2.967438, 3.063721, 2.846039, 2.976624, 3.1922, 2.912109, 2.313416, 
    2.356812, 2.402618, 2.267456, 2.22168, 2.102661, 2.133881, 1.972198, 
    1.992493, 2.573395, 2.717651, 2.802185, 3.008667, 2.830048, 2.760254, 
    2.691223, 2.682281, 2.697418, 2.718842, 2.680176, 2.592621, 2.509796, 
    2.474579, 2.485596, 2.512421, 2.50766, 2.459412, 2.365387, 2.238525, 
    2.123932, 2.02359, 1.960449, 1.959198, 1.971893, 1.935913, 2.013123, 
    1.92627, 1.833191, 1.983002, 2.375458, 2.637054, 2.639832, 2.662231, 
    2.945404, 2.992554, 3.30484, 3.5784, 3.462067, 3.842621, 3.722107, 
    3.687622, 3.322083, 3.139557, 2.843842, 2.682434, 2.645935, 2.29306, 
    1.929718, 1.661499, 1.274689, 0.9851685, 1.147339, 1.52121, 1.913605, 
    2.06134, 1.965881, 2.063843, 2.834747, 3.326721,
  2.736481, 2.980438, 3.073639, 3.107666, 2.806335, 2.603912, 2.386963, 
    2.545319, 2.622345, 2.60968, 2.698334, 2.551666, 2.324524, 2.250671, 
    2.075287, 2.212646, 2.150848, 2.170593, 2.191345, 2.171326, 2.329865, 
    2.317383, 1.993622, 1.905518, 2.163971, 1.989624, 2.09436, 2.082367, 
    1.961456, 1.988037, 2.001617, 1.983856, 1.997314, 1.958649, 1.897339, 
    1.9086, 2.128723, 2.540894, 2.611023, 2.694824, 2.506104, 2.514801, 
    2.478455, 2.399445, 2.393311, 2.431, 2.455902, 2.438965, 2.430695, 
    2.464447, 2.471313, 2.424194, 2.359741, 2.320862, 2.315918, 2.307465, 
    2.225159, 2.091827, 1.97821, 1.932983, 1.898468, 1.845581, 1.969177, 
    1.981995, 1.965698, 1.91861, 2.003387, 2.207367, 2.447021, 2.709412, 
    2.929199, 2.976105, 3.141998, 3.392609, 3.561554, 3.588196, 3.535736, 
    3.539398, 3.488037, 3.371582, 3.09079, 2.70285, 2.02179, 1.775757, 
    1.755371, 1.68219, 1.280701, 0.8269958, 0.6974487, 0.9165649, 1.336029, 
    1.732452, 1.854065, 1.944153, 2.141174, 2.565338,
  2.465393, 2.634186, 2.800323, 2.917633, 2.84375, 2.645386, 2.430939, 
    2.460571, 2.494476, 2.542145, 2.482819, 2.275848, 2.031494, 1.875122, 
    1.762115, 1.612, 1.702789, 1.830261, 1.600586, 1.561066, 1.827728, 
    1.933258, 1.977722, 2.109436, 1.897949, 1.687134, 1.550659, 2.022736, 
    1.959442, 2.004059, 2.261292, 2.221893, 2.12561, 2.164673, 2.251251, 
    2.383362, 2.319092, 2.069214, 1.997711, 2.166992, 2.409729, 2.474945, 
    2.419312, 2.294708, 2.223083, 2.273041, 2.349945, 2.429779, 2.477173, 
    2.487793, 2.46759, 2.469604, 2.513916, 2.530365, 2.50766, 2.460724, 
    2.373322, 2.244904, 2.115723, 2.003601, 1.901978, 1.935455, 2.107849, 
    2.258575, 2.330414, 2.074432, 2.0383, 2.131622, 2.327545, 2.613678, 
    2.787048, 2.897125, 3.016663, 3.190674, 3.458649, 3.657501, 3.660797, 
    3.654541, 3.57962, 3.361908, 3.135071, 2.944458, 2.17572, 1.982269, 
    1.846344, 1.535767, 1.009674, 0.2644958, -0.10849, 0.09997559, 0.6495667, 
    1.216614, 1.534729, 1.679199, 1.841949, 2.012909,
  2.349701, 1.914886, 2.231293, 2.450226, 2.750397, 2.728119, 2.598236, 
    2.344971, 2.196136, 2.083527, 1.983154, 1.774048, 1.652039, 1.741882, 
    1.620361, 1.393158, 1.31955, 1.315369, 1.213348, 1.049286, 1.154053, 
    1.390808, 1.832397, 2.244354, 2.279175, 2.039795, 2.002991, 2.180145, 
    2.257111, 2.58075, 2.665649, 3.03476, 2.811554, 2.652039, 2.779053, 
    3.087921, 3.014069, 2.329437, 1.937683, 2.043121, 2.343689, 2.509979, 
    1.915558, 2.10321, 2.051178, 2.241669, 2.33728, 2.421478, 2.485138, 
    2.516113, 2.54068, 2.632721, 2.769379, 2.82959, 2.742401, 2.608429, 
    2.509216, 2.411682, 2.27887, 2.11026, 1.907837, 1.992188, 2.098969, 
    2.328918, 2.216217, 1.984558, 1.962128, 2.019196, 2.216797, 2.539063, 
    2.789581, 3.046875, 3.234283, 3.316589, 3.486786, 3.820251, 3.873047, 
    3.919067, 3.792664, 3.549164, 3.153778, 2.253754, 1.915314, 1.570251, 
    1.411346, 1.391785, 1.118683, 0.5315552, 0.06240845, 0.07839966, 
    0.553894, 1.060059, 1.352386, 1.520264, 2.008972, 2.262726,
  1.457458, 1.70166, 1.580109, 2.169922, 2.149353, 2.113495, 1.996704, 
    2.301422, 2.289886, 2.144989, 1.875977, 1.710999, 1.626495, 1.490692, 
    1.379425, 1.355011, 1.343109, 1.33075, 1.343872, 1.314514, 1.343353, 
    1.471802, 1.687439, 1.881592, 2.05777, 2.221893, 2.371765, 2.581146, 
    3.117493, 3.352478, 3.729126, 3.832092, 3.67215, 3.674683, 3.980042, 
    3.87619, 3.235504, 2.705078, 2.075836, 2.108795, 2.236633, 2.251678, 
    2.28009, 2.305817, 2.145447, 2.506683, 2.743805, 2.736206, 2.86734, 
    2.997925, 3.085938, 3.097321, 3.042847, 2.980713, 2.938416, 2.496521, 
    2.421448, 2.403809, 2.301392, 2.104919, 2.024414, 2.316742, 2.851685, 
    2.453522, 2.027191, 1.764648, 1.731995, 1.968353, 2.441986, 2.746887, 
    2.85025, 3.046722, 2.963623, 3.098236, 3.373169, 3.733276, 4.224731, 
    3.924225, 3.652618, 3.531036, 2.063934, 1.766357, 1.430145, 1.187958, 
    1.317627, 1.381073, 1.46701, 1.301575, 1.01178, 0.9371948, 1.08316, 
    1.259277, 1.334656, 1.338959, 1.454742, 1.83194,
  1.314728, 1.608429, 2.056976, 2.138855, 2.09082, 1.790802, 2.137573, 
    2.185669, 2.163422, 2.125061, 2.032806, 1.846954, 1.709961, 1.671356, 
    1.562042, 1.447449, 1.546112, 1.65567, 1.676971, 1.828339, 1.970734, 
    2.092682, 2.2258, 2.438477, 2.724487, 3.14624, 3.469696, 3.620422, 
    3.608887, 3.731049, 4.00061, 4.74234, 5.286591, 5.578674, 5.616302, 
    5.326569, 4.601379, 4.13327, 4.236145, 3.950165, 3.731262, 3.77951, 
    3.960388, 4.637329, 4.656189, 4.181396, 3.84906, 2.761993, 3.224823, 
    3.554504, 3.538086, 3.268677, 3.177521, 3.021393, 2.825409, 2.671234, 
    2.695587, 3.09787, 3.395844, 3.366425, 3.0047, 2.758728, 2.475342, 
    2.018005, 1.780487, 1.80542, 2.150604, 2.559448, 2.853729, 2.911072, 
    2.996735, 2.673248, 2.78717, 2.876312, 3.043945, 3.141876, 4.311066, 
    4.397339, 2.897919, 2.35965, 1.807556, 1.447144, 1.208801, 1.063232, 
    2.341278, 0.9905396, 1.406128, 1.492371, 1.534851, 1.53714, 1.471771, 
    1.369629, 1.208038, 1.036041, 1.147156, 1.241455,
  0.9204712, 0.8964539, 0.9129028, 1.670135, 1.88443, 2.058197, 1.654297, 
    2.267517, 2.370331, 2.342987, 2.35318, 2.439972, 2.503967, 2.549347, 
    2.620514, 2.60611, 2.623047, 2.672211, 2.570313, 2.53244, 2.593109, 
    2.68219, 3.005737, 3.414276, 3.734955, 4.185425, 4.485504, 4.631073, 
    4.804199, 5.700104, 6.062378, 6.120972, 6.188385, 5.83551, 5.654968, 
    5.54187, 4.388565, 4.559341, 4.366867, 4.349945, 4.724548, 4.24469, 
    4.541992, 4.556183, 4.457184, 4.675476, 5.15033, 5.926239, 6.520081, 
    6.090515, 5.186646, 3.235413, 3.175262, 2.972961, 3.078156, 3.184998, 
    3.441956, 3.590363, 3.549103, 3.427765, 3.308655, 3.015991, 2.658783, 
    2.489471, 2.514465, 2.72287, 3.120087, 3.376373, 3.664215, 4.239197, 
    4.816223, 5.243103, 5.182312, 5.011017, 4.460693, 3.920319, 3.571289, 
    5.519623, 5.158295, 4.206024, 1.936371, 1.687744, 3.186218, 3.343903, 
    3.256714, 3.111298, 2.746002, 1.160156, 1.218231, 1.22052, 1.170898, 
    1.786652, 1.073639, 0.7854919, 0.765564, 0.7833252,
  1.094666, 1.113739, 1.136475, 1.151611, 1.04837, 2.094147, 2.283722, 
    2.367249, 2.391083, 2.480682, 2.429016, 1.897186, 1.950989, 2.089905, 
    3.000854, 3.442078, 3.982178, 4.393036, 4.398956, 4.07254, 3.94696, 
    3.901306, 4.045898, 4.264923, 4.651703, 4.738892, 5.09024, 5.394745, 
    5.844482, 6.491669, 6.955429, 6.883881, 6.546036, 6.019821, 4.881439, 
    4.73465, 5.557175, 4.871429, 6.514725, 6.990173, 7.770477, 7.899368, 
    7.717667, 7.792648, 5.835907, 5.793182, 6.349884, 7.654495, 8.524506, 
    10.62366, 7.739044, 5.882111, 5.362823, 5.404388, 5.407379, 5.139496, 
    5.208221, 5.264587, 4.975708, 4.494202, 4.235443, 4.561859, 4.888367, 
    5.164673, 5.427124, 5.336212, 5.162262, 5.242462, 5.395996, 3.093079, 
    5.122284, 4.758484, 5.01062, 3.259857, 5.990356, 6.638123, 7.167786, 
    6.842072, 5.585541, 2.913757, 1.985504, 1.788483, 3.669739, 4.21669, 
    4.671387, 4.620682, 4.429123, 4.075104, 3.636078, 3.559723, 2.18573, 
    2.048431, 1.79895, 1.492828, 1.22934, 1.154358,
  1.826569, 1.52533, 1.398834, 1.318359, 1.280548, 1.478882, 1.880219, 
    2.236023, 2.39447, 2.374878, 2.284821, 2.23053, 2.35144, 2.680267, 
    3.154175, 6.054749, 6.852631, 7.184845, 7.146515, 6.149902, 5.380798, 
    5.342163, 5.421631, 5.602295, 5.579376, 5.662628, 5.863083, 5.940887, 
    6.144028, 6.936813, 7.266693, 7.638214, 7.831711, 7.981201, 7.844788, 
    7.234436, 7.070709, 7.007568, 7.834778, 8.458206, 10.3217, 10.65686, 
    10.83427, 11.24352, 11.64644, 11.86284, 12.08087, 12.66571, 13.41942, 
    14.16364, 14.28999, 13.53004, 12.53444, 11.72125, 11.2596, 10.91936, 
    10.75412, 10.5838, 10.26993, 9.864777, 9.503845, 9.119476, 8.61441, 
    8.126648, 7.908081, 7.670349, 7.514801, 7.1698, 6.592072, 4.00946, 
    5.803864, 6.095734, 4.22345, 7.362213, 8.453613, 9.198273, 9.904312, 
    9.814789, 7.708801, 4.827728, 3.039551, 4.691986, 4.702164, 5.275879, 
    5.792542, 5.385361, 4.467682, 4.300613, 4.726196, 5.254852, 5.816284, 
    6.755219, 5.345856, 3.39389, 2.536224, 2.178375,
  2.707092, 2.165375, 2.015106, 2.11908, 2.156708, 2.470917, 2.955078, 
    3.639069, 4.034637, 4.643494, 5.431, 6.165833, 6.948395, 7.858368, 
    8.680023, 9.340912, 9.665131, 9.622162, 9.290131, 8.768372, 7.987671, 
    7.336823, 6.829559, 6.531677, 6.466949, 6.611359, 6.950928, 7.789474, 
    8.236481, 8.961426, 9.314529, 10.033, 10.37384, 10.39622, 10.60387, 
    10.52985, 10.22124, 9.910446, 9.822922, 9.648788, 9.730759, 9.768509, 
    9.914932, 10.10698, 10.21129, 10.23029, 10.30717, 10.44756, 10.61842, 
    10.7084, 10.74232, 10.68883, 10.63356, 10.5004, 10.41922, 10.42047, 
    10.50307, 10.52827, 10.60197, 10.67931, 10.76076, 10.7758, 10.70888, 
    10.67052, 10.27, 9.05542, 8.692719, 8.233475, 7.908157, 7.918106, 
    7.988617, 9.321762, 9.954697, 10.32437, 10.4476, 12.77716, 12.86426, 
    10.84937, 7.78804, 6.572556, 5.682312, 5.26651, 5.39241, 5.794693, 
    5.629715, 4.752518, 4.281479, 4.47464, 4.939163, 5.63942, 6.506149, 
    7.014206, 9.510941, 8.622467, 7.097198, 4.714142,
  8.062256, 7.862274, 7.394806, 6.650208, 6.610229, 6.784119, 6.942017, 
    8.292206, 8.533936, 8.525085, 8.625275, 8.737457, 8.865631, 8.948914, 
    8.915955, 8.858032, 8.737823, 8.503723, 8.397278, 8.331512, 8.283752, 
    8.215317, 8.120148, 7.885056, 7.428772, 7.797531, 7.90979, 8.547531, 
    8.800415, 9.118561, 9.456909, 9.739349, 9.878342, 9.841629, 9.748734, 
    9.58165, 9.365768, 9.179428, 8.97757, 8.850082, 8.752029, 8.563934, 
    8.46402, 8.390778, 8.350525, 8.302353, 8.283951, 8.337402, 8.420776, 
    8.504044, 8.567474, 8.661743, 8.74826, 8.835831, 8.917862, 8.903717, 
    8.924316, 8.968246, 9.125793, 9.301575, 9.478027, 9.578583, 9.669678, 
    9.828018, 9.847214, 9.688232, 9.534134, 9.308929, 9.048645, 8.858139, 
    8.468262, 7.901779, 7.575394, 7.569565, 7.089157, 6.675552, 6.078995, 
    5.617081, 5.289993, 5.064423, 4.998413, 5.037399, 5.213699, 5.33812, 
    5.323135, 5.324905, 5.36293, 5.672043, 6.045471, 6.609024, 7.114746, 
    7.484085, 9.003479, 9.060577, 8.779968, 8.44104,
  7.726135, 7.56813, 7.534393, 7.487381, 7.487793, 7.49202, 7.480484, 
    7.57254, 7.686005, 7.753998, 7.789322, 7.798569, 7.776703, 7.778397, 
    7.801117, 7.829132, 7.839844, 7.88446, 7.938309, 8.019562, 8.115707, 
    8.222656, 8.312958, 8.417145, 8.455292, 8.48407, 8.525208, 8.535385, 
    8.586411, 8.633804, 8.664871, 8.696121, 8.676773, 8.666016, 8.625488, 
    8.542938, 8.462646, 8.386734, 8.291489, 8.194992, 8.126511, 8.076462, 
    8.069626, 8.084183, 8.118103, 8.144943, 8.129044, 8.114471, 8.114151, 
    8.13002, 8.16774, 8.192276, 8.21199, 8.200989, 8.196838, 8.205994, 
    8.202103, 8.207428, 8.28862, 8.40712, 8.579773, 8.768906, 8.925858, 
    9.054962, 9.146835, 9.195313, 9.179688, 9.16713, 9.140976, 9.111664, 
    9.083023, 9.064743, 8.928497, 8.876526, 8.794312, 8.819885, 8.88974, 
    8.886108, 8.972748, 9.026077, 9.12471, 9.058304, 9.098465, 9.067352, 
    9.234726, 9.421127, 9.562531, 9.589615, 9.637146, 9.289551, 9.033615, 
    8.730835, 8.608047, 8.40625, 8.138351, 7.875931,
  7.747986, 7.622162, 7.697266, 7.781281, 7.809204, 7.800003, 7.81778, 
    7.804047, 7.791748, 7.805023, 7.800201, 7.839859, 7.88739, 7.908539, 
    7.945206, 7.95491, 7.977097, 7.99942, 8.038116, 8.045273, 8.04213, 
    8.06134, 8.094559, 8.132645, 8.144867, 8.140244, 8.135818, 8.162628, 
    8.166885, 8.132965, 8.08342, 8.059402, 8.020203, 7.979965, 7.943375, 
    7.875214, 7.837006, 7.837967, 7.815781, 7.783051, 7.73082, 7.67189, 
    7.613846, 7.574448, 7.555237, 7.548538, 7.539291, 7.512924, 7.509399, 
    7.461945, 7.42836, 7.41124, 7.426529, 7.428024, 7.426849, 7.429199, 
    7.477646, 7.544693, 7.59996, 7.634354, 7.687088, 7.76651, 7.839417, 
    7.93251, 7.99678, 8.063507, 8.183105, 8.29332, 8.396317, 8.472229, 
    8.544495, 8.608231, 8.630493, 8.63916, 8.680435, 8.667816, 8.687073, 
    8.707001, 8.711029, 8.706482, 8.678741, 8.651657, 8.606339, 8.585052, 
    8.545807, 8.524765, 8.476257, 8.433105, 8.417877, 8.400162, 8.347427, 
    8.300888, 8.242401, 8.155548, 8.007767, 7.907578,
  2.340805, 2.328171, 2.318268, 2.309021, 2.299713, 2.294708, 2.29158, 
    2.284622, 2.28273, 2.279221, 2.279022, 2.275116, 2.271729, 2.270615, 
    2.267883, 2.269257, 2.267624, 2.267288, 2.263718, 2.26091, 2.257278, 
    2.249985, 2.246399, 2.245621, 2.235138, 2.22934, 2.22049, 2.218399, 
    2.215988, 2.214432, 2.208893, 2.200958, 2.190536, 2.17485, 2.160797, 
    2.144394, 2.129288, 2.116516, 2.104538, 2.093277, 2.084351, 2.082474, 
    2.08287, 2.079346, 2.077271, 2.0755, 2.069839, 2.068405, 2.07283, 
    2.077393, 2.077652, 2.077911, 2.061905, 2.054138, 2.046936, 2.053375, 
    2.072571, 2.069199, 2.072845, 2.0634, 2.070297, 2.110992, 2.106827, 
    2.123749, 2.142426, 2.16066, 2.186508, 2.231552, 2.268539, 2.301743, 
    2.331818, 2.361252, 2.391449, 2.396667, 2.414368, 2.426483, 2.43631, 
    2.456116, 2.467377, 2.473999, 2.476089, 2.476486, 2.481354, 2.486252, 
    2.489243, 2.491913, 2.492889, 2.48912, 2.480713, 2.470428, 2.453308, 
    2.435471, 2.414703, 2.394379, 2.37413, 2.353699,
  2.257141, 2.225571, 2.21463, 2.232727, 2.269196, 2.341843, 2.423752, 
    2.509293, 2.593277, 2.667694, 2.718597, 2.757401, 2.79068, 2.814896, 
    2.833069, 2.865997, 2.897308, 2.930389, 2.944443, 2.929855, 2.896591, 
    2.854858, 2.8078, 2.7509, 2.701218, 2.660538, 2.601486, 2.527191, 
    2.447968, 2.367111, 2.294388, 2.23735, 2.203568, 2.184097, 2.168594, 
    2.161118, 2.157074, 2.161377, 2.166382, 2.184875, 2.222, 2.260345, 
    2.306763, 2.350571, 2.386246, 2.431549, 2.474396, 2.528564, 2.574524, 
    2.605988, 2.640213, 2.654724, 2.67244, 2.664627, 2.724533, 2.657013, 
    2.640091, 2.628433, 2.590942, 2.553757, 2.501358, 2.448624, 2.417175, 
    2.408447, 2.418732, 2.437744, 2.468933, 2.520874, 2.601868, 2.675369, 
    2.669312, 2.6315, 2.567108, 2.504272, 2.52504, 2.52478, 2.552795, 
    2.55336, 2.593414, 2.537033, 2.433197, 2.399658, 2.273682, 2.288986, 
    2.23735, 2.264893, 2.300705, 2.354279, 2.41156, 2.450897, 2.460663, 
    2.445816, 2.408569, 2.36145, 2.319443, 2.28775,
  2.434952, 2.447769, 2.455185, 2.475632, 2.440811, 2.354202, 2.263336, 
    2.195496, 2.193405, 2.285202, 2.427399, 2.545288, 2.61438, 2.645233, 
    2.678436, 2.709824, 2.732666, 2.719177, 2.663849, 2.588135, 2.520218, 
    2.466919, 2.418793, 2.422119, 2.515411, 2.622253, 2.70903, 2.744507, 
    2.759293, 2.730194, 2.677979, 2.596725, 2.517563, 2.467697, 2.430847, 
    2.419571, 2.42186, 2.434753, 2.452255, 2.482086, 2.514236, 2.520493, 
    2.535721, 2.573563, 2.626938, 2.624207, 2.546082, 2.50148, 2.516129, 
    2.538391, 2.529602, 2.470673, 2.413666, 2.408188, 2.483246, 2.558182, 
    2.526733, 2.421997, 2.34816, 2.252213, 2.191971, 2.153442, 2.158569, 
    2.123749, 2.035461, 1.964569, 1.956757, 2.076096, 2.184677, 2.267624, 
    2.262482, 2.218658, 2.173752, 2.159103, 2.194138, 2.216644, 2.237289, 
    2.162811, 2.085541, 1.973297, 1.910995, 1.906342, 1.917725, 1.893204, 
    1.859085, 1.86351, 1.854279, 1.87616, 1.933716, 2.025436, 2.077515, 
    2.143402, 2.174789, 2.217941, 2.286514, 2.364563,
  2.349991, 2.329407, 2.303833, 2.238983, 2.162674, 2.114899, 2.18689, 
    2.355637, 2.493408, 2.615677, 2.743286, 2.856567, 2.931366, 2.941788, 
    2.963272, 3.057602, 3.158112, 3.267563, 3.321609, 3.268799, 3.119583, 
    2.850174, 2.508514, 2.178696, 1.972061, 1.923813, 1.968475, 2.012344, 
    2.043793, 2.071274, 2.089966, 2.100449, 2.106628, 2.156815, 2.2397, 
    2.336502, 2.411957, 2.437088, 2.47023, 2.512619, 2.522766, 2.519257, 
    2.497055, 2.488663, 2.526611, 2.619202, 1.544281, 1.45639, 1.450684, 
    1.47287, 1.448486, 1.456604, 1.455566, 1.402039, 1.376801, 1.340668, 
    1.28479, 1.464355, 1.519958, 1.634827, 1.773041, 1.853424, 1.981949, 
    2.073685, 2.112274, 2.099457, 2.08696, 2.051544, 2.071854, 2.132339, 
    2.150635, 2.178497, 2.181747, 2.170837, 2.170486, 2.137787, 2.101486, 
    2.077072, 2.164337, 2.149918, 2.257446, 2.215393, 2.188965, 2.08075, 
    2.050812, 2.08252, 2.19989, 2.253998, 2.521667, 2.287552, 2.30983, 
    2.260208, 2.253815, 2.250244, 2.295044, 2.326736,
  2.247498, 2.221146, 2.191772, 2.201599, 2.192184, 2.195694, 2.245895, 
    2.207794, 2.240616, 2.296463, 2.420364, 2.452072, 2.435867, 2.486435, 
    2.614105, 2.649536, 2.548492, 2.463272, 2.406631, 2.352127, 2.380447, 
    2.287491, 2.123947, 2.020813, 2.028442, 2.087296, 2.204987, 2.261368, 
    2.292633, 2.350967, 2.408829, 2.430649, 2.431488, 2.421143, 2.487213, 
    2.560928, 2.582993, 2.532669, 2.434097, 2.298553, 2.156769, 2.105576, 
    2.108978, 2.077591, 2.045242, 2.023605, 1.347534, 1.212006, 1.074829, 
    0.9833069, 0.8661194, 0.7590637, 0.681488, 0.6644897, 0.6473083, 
    0.6036072, 0.6094666, 0.6820679, 0.7894897, 0.8997803, 1.020752, 
    1.140411, 1.234222, 1.265472, 1.289032, 1.333557, 1.456085, 1.513855, 
    1.51767, 1.354065, 2.579468, 2.491913, 2.405182, 2.214935, 2.044373, 
    1.723206, 2.249115, 2.120361, 2.096436, 2.036682, 1.824982, 1.623657, 
    1.50473, 1.464661, 1.503754, 1.617035, 1.850037, 2.016754, 2.193787, 
    2.380096, 2.559418, 2.461639, 2.444382, 2.462814, 2.483063, 2.358582,
  2.304596, 2.162476, 2.439606, 2.324585, 2.16217, 1.996002, 1.993668, 
    2.23494, 2.275818, 2.203339, 2.263367, 2.334412, 2.278381, 2.245239, 
    2.145035, 2.124725, 2.175766, 2.095428, 1.944962, 1.851746, 1.880981, 
    1.847961, 1.712021, 1.656097, 1.654602, 1.662094, 1.669189, 1.768997, 
    1.865158, 1.902328, 1.89537, 1.892761, 1.965088, 2.022705, 2.032028, 
    1.94075, 1.797119, 1.714966, 1.70871, 1.671921, 1.701355, 1.66835, 
    1.523483, 1.391205, 1.093781, 0.8378601, 0.6091003, 0.3257446, 0.1829834, 
    0.07003784, 0.04278564, -0.01293945, 0.01586914, 0.02230835, 0.08276367, 
    0.1254272, 0.2121887, 0.3093872, 0.4471741, 0.5738525, 0.7514648, 
    0.8865051, 1.09549, 1.241486, 1.398804, 1.525574, 1.638245, 1.774384, 
    1.888428, 1.979065, 2.225616, 2.506744, 2.483246, 2.36792, 2.152557, 
    1.879456, 1.644684, 1.29776, 2.077881, 2.223816, 1.976013, 1.800964, 
    1.627716, 1.523132, 1.507507, 1.613586, 1.863983, 2.02771, 2.094879, 
    2.148987, 2.184723, 2.194946, 2.314941, 2.455292, 2.51178, 2.452179,
  2.432648, 2.486084, 2.564209, 2.626862, 2.636475, 2.541748, 2.474457, 
    2.443329, 2.485199, 2.458496, 2.450226, 2.523773, 2.538727, 2.545258, 
    2.468384, 2.362915, 2.370667, 2.366516, 2.385071, 2.292694, 2.148682, 
    2.046326, 1.983368, 1.930786, 1.927765, 1.811951, 1.682129, 1.526123, 
    1.38797, 1.303314, 1.283813, 1.301605, 1.170685, 2.078674, 2.218262, 
    2.374268, 2.009888, 1.942596, 1.862213, 1.777069, 1.752319, 1.676331, 
    1.538116, 1.342987, 1.098602, 0.8243103, 0.5112305, 0.2878418, 
    0.07391357, -0.07849121, -0.1992493, -0.2601929, -0.2518005, -0.2532959, 
    -0.2540283, -0.1167908, 0.0272522, 0.1303711, 0.2420349, 0.3500366, 
    0.4710083, 0.6471252, 0.8730164, 1.121857, 1.393188, 1.679199, 1.926941, 
    2.122681, 2.25766, 2.526184, 2.739288, 2.92926, 2.995605, 2.94165, 
    2.786621, 2.593109, 2.439484, 2.338104, 2.370087, 2.459595, 2.210754, 
    1.946014, 1.76004, 1.68689, 1.739075, 1.865448, 2.026581, 2.190277, 
    2.316315, 2.328217, 2.295502, 2.255127, 2.343994, 2.484619, 2.553314, 
    2.464172,
  2.205261, 2.170776, 2.139923, 2.111694, 2.133301, 2.152771, 2.096313, 
    2.080566, 2.007599, 2.002563, 2.057709, 2.32132, 2.625427, 2.756104, 
    2.70459, 2.508881, 2.494629, 2.638428, 2.539154, 2.35556, 2.173462, 
    2.005371, 1.972412, 1.952759, 1.910065, 1.751923, 1.47699, 1.173737, 
    0.9309082, 0.8164368, 0.7448425, 0.6773071, 0.6812439, 0.7846069, 
    0.9705505, 1.392395, 1.603485, 1.593903, 1.572357, 1.428558, 1.295746, 
    1.258545, 1.291748, 1.278168, 1.152771, 0.9690552, 0.7775269, 0.5960693, 
    0.2290039, -0.2330322, -0.574707, -0.7097473, -0.721283, -0.6777954, 
    -0.4821167, -0.2687988, -0.07867432, 0.005828857, 0.03265381, 0.1315308, 
    0.3496704, 0.5439758, 0.7420349, 1.039917, 1.343933, 1.645111, 1.912231, 
    2.142303, 2.404755, 2.681824, 2.964447, 3.108643, 3.161896, 3.149963, 
    3.160614, 3.146576, 3.010864, 2.757294, 2.484467, 2.05069, 1.800751, 
    1.676208, 1.616089, 1.605377, 1.5896, 1.545074, 1.633179, 1.822601, 
    1.926392, 1.928558, 1.924255, 1.972015, 2.03421, 2.092102, 2.160583, 
    2.19458,
  1.633484, 1.609192, 1.543274, 1.556854, 1.647736, 1.656677, 1.700684, 
    1.761963, 1.754852, 1.731567, 1.685394, 1.770782, 1.944366, 2.054016, 
    2.187653, 2.307983, 2.437286, 2.503387, 2.49353, 2.521515, 2.475494, 
    2.308289, 2.169281, 2.098938, 2.008423, 1.829529, 1.478821, 1.126862, 
    0.9770508, 0.915863, 0.8292847, 0.8033142, 0.7989197, 0.7616882, 
    0.7081604, 0.7319946, 1.022156, 1.349854, 1.543518, 1.569183, 1.535522, 
    1.734741, 2.12796, 2.262787, 2.053284, 1.844757, 1.570282, 1.154205, 
    0.6148682, -0.1017761, -0.4838257, -0.4816589, -0.4316711, -0.4761963, 
    -0.5662231, -0.583252, -0.5875854, -0.605835, -0.3517761, 0.1503601, 
    0.5782166, 0.9100037, 1.225891, 1.566254, 1.849762, 2.015015, 2.19339, 
    2.379639, 2.500671, 2.614563, 2.701996, 2.753693, 2.794952, 2.774078, 
    2.654327, 2.404938, 1.950592, 1.753693, 1.712982, 1.726074, 1.715698, 
    1.681274, 1.528961, 1.256622, 1.115417, 1.137146, 1.269379, 1.496063, 
    1.598999, 1.638184, 1.77063, 1.879272, 1.883026, 1.735382, 1.599457, 
    1.616455,
  1.494904, 1.603241, 1.78833, 2.049744, 2.128632, 2.153503, 2.169006, 
    2.227875, 2.321198, 2.332184, 2.275574, 2.231476, 2.220978, 2.283386, 
    2.440186, 2.615479, 2.808563, 3.022369, 2.987549, 2.512299, 2.123199, 
    1.940552, 1.778229, 1.75351, 1.79248, 1.754852, 1.768921, 1.790649, 
    1.790527, 1.802246, 1.718903, 1.529694, 1.342224, 1.209229, 1.145813, 
    1.219574, 1.459717, 1.803497, 1.999634, 1.99704, 1.961548, 2.073608, 
    2.208374, 2.138245, 1.946381, 1.865417, 1.845215, 1.691711, 1.401947, 
    0.9627075, 0.7084961, 0.6669617, 0.5440674, 0.365509, 0.2635803, 
    0.2227478, 0.2122192, 0.2866211, 0.4537964, 0.6844788, 0.9113464, 
    1.065582, 1.226013, 1.425415, 1.574921, 1.617279, 1.721436, 1.873199, 
    1.978027, 2.05011, 2.109741, 2.133118, 2.146698, 2.08252, 1.841827, 
    1.389465, 1.436371, 2.230042, 2.408752, 1.876587, 1.682526, 1.581696, 
    1.612793, 1.497742, 1.300812, 1.353271, 1.537079, 1.662018, 1.657837, 
    1.660706, 1.662689, 1.704865, 1.715271, 1.669403, 1.609497, 1.506317,
  1.991821, 2.166504, 2.319641, 2.438629, 2.52179, 2.541656, 2.594635, 
    2.67984, 2.747681, 2.83493, 2.918396, 2.960114, 2.984589, 2.996002, 
    3.010254, 3.045074, 3.193268, 3.475342, 3.607178, 3.352905, 3.042358, 
    2.853241, 2.669373, 2.457275, 2.363129, 2.356873, 2.359283, 2.262054, 
    2.187012, 2.174377, 2.123871, 1.948486, 1.690277, 1.517151, 1.488495, 
    1.545288, 1.65094, 1.730621, 1.755249, 1.845215, 2.05603, 2.245941, 
    2.238312, 2.090454, 2.078278, 2.123291, 2.071533, 1.992249, 1.877594, 
    1.739502, 1.592072, 1.381165, 1.156494, 1.035645, 1.040802, 1.024628, 
    1.03183, 1.074829, 1.163574, 1.249695, 1.312714, 1.358307, 1.416046, 
    1.48465, 1.561554, 1.582397, 1.58728, 1.60675, 1.620026, 1.659821, 
    1.683899, 1.652771, 1.592682, 1.495056, 1.313721, 1.306244, 1.818054, 
    2.054352, 2.030701, 1.865265, 1.572754, 1.437988, 1.474426, 1.434814, 
    1.383118, 1.540009, 1.75235, 1.949707, 2.064819, 2.133301, 2.101318, 
    2.01123, 1.951965, 1.940857, 1.937073, 1.906921,
  2.062683, 2.249969, 2.407623, 2.501068, 2.538177, 2.619171, 2.845612, 
    3.064728, 3.144897, 3.253235, 3.427643, 3.492401, 3.450806, 3.377563, 
    3.298065, 3.226685, 3.200623, 3.266632, 3.362793, 3.474884, 3.775269, 
    3.992096, 3.785187, 3.293762, 2.961426, 2.751526, 2.51123, 2.277374, 
    2.110962, 1.98526, 1.873077, 1.724762, 1.596466, 1.57608, 1.593781, 
    1.612976, 1.617157, 1.527374, 1.428558, 1.600159, 2.060577, 2.354004, 
    2.425903, 2.330811, 2.500763, 2.684998, 2.547302, 2.411163, 2.292786, 
    2.275818, 2.23056, 2.079468, 1.878174, 1.728943, 1.672302, 1.638184, 
    1.591095, 1.574127, 1.570801, 1.543396, 1.562592, 1.605438, 1.568512, 
    1.54364, 1.536407, 1.489319, 1.451843, 1.417999, 1.330963, 1.289154, 
    1.306458, 1.327698, 1.329437, 1.2771, 1.196533, 1.243317, 1.755005, 
    2.121246, 2.306213, 1.716949, 1.423218, 1.337524, 1.475372, 1.549377, 
    1.516632, 1.567078, 1.579407, 1.628937, 1.770264, 1.836334, 1.81134, 
    1.789154, 1.771973, 1.779633, 1.833435, 1.921326,
  2.143524, 2.266479, 2.378998, 2.460724, 2.571136, 2.882843, 3.430634, 
    3.839691, 4.011047, 4.176727, 4.336945, 4.239868, 3.895844, 3.583038, 
    3.359344, 3.203339, 3.11084, 3.05127, 3.083954, 3.181091, 3.214569, 
    3.113129, 2.763123, 2.329956, 2.06424, 1.937286, 1.805969, 1.692352, 
    1.632446, 1.592163, 1.56781, 1.567291, 1.529999, 1.476868, 1.402252, 
    1.398163, 1.438721, 1.421295, 1.580566, 1.913177, 2.359161, 2.563049, 
    2.659607, 2.594482, 2.693848, 2.871002, 2.948181, 2.750366, 2.721893, 
    2.756134, 2.916748, 2.778931, 2.496826, 2.231415, 2.020935, 1.89859, 
    1.80304, 1.664856, 1.565582, 1.536957, 1.569305, 1.596191, 1.543243, 
    1.513489, 1.509216, 1.424896, 1.365265, 1.33902, 1.297607, 1.347015, 
    1.379395, 1.394043, 1.419647, 1.383636, 1.303986, 1.232452, 1.433167, 
    1.937988, 2.393372, 1.751526, 1.40509, 1.288055, 1.491028, 1.760254, 
    1.788391, 1.718353, 1.6297, 1.624329, 1.741638, 1.799316, 1.778229, 
    1.813446, 1.81839, 1.790833, 1.86972, 2.016174,
  2.1203, 2.137207, 2.129913, 2.166748, 2.411896, 2.888123, 3.17627, 
    3.611084, 3.785828, 3.537476, 3.065796, 2.673981, 2.357147, 2.175171, 
    2.073822, 2.062317, 2.046906, 1.992523, 1.926514, 1.845215, 1.766937, 
    1.656982, 1.503418, 1.359711, 1.24704, 1.252045, 1.295807, 1.310699, 
    1.391846, 1.5896, 1.804077, 1.726807, 1.565643, 1.339996, 1.210052, 
    1.378998, 1.635559, 1.81366, 2.153992, 3.554993, 2.605133, 2.880005, 
    3.134918, 2.973206, 2.877594, 2.941559, 2.921967, 3.03302, 2.764496, 
    2.521606, 2.343597, 2.168243, 2.056671, 1.951935, 1.781281, 1.721191, 
    1.675415, 1.542938, 1.517212, 1.570679, 1.615997, 1.621582, 1.546906, 
    1.530884, 1.560333, 1.524902, 1.52533, 1.498383, 1.491058, 1.547485, 
    1.52536, 1.558685, 1.55426, 1.437286, 1.335907, 1.175568, 1.378143, 
    2.537842, 2.550751, 1.912476, 1.417755, 1.421326, 1.843414, 2.179779, 
    2.084198, 1.884094, 1.81427, 1.743317, 1.748077, 1.768463, 1.799591, 
    1.860443, 1.84256, 1.843964, 1.891632, 1.997955,
  1.874512, 1.796204, 1.838837, 2.002716, 2.353271, 2.526978, 2.532379, 
    2.63089, 2.866943, 2.413269, 1.773651, 1.576721, 1.654266, 1.714142, 
    1.600159, 1.503143, 1.479401, 1.435486, 1.370667, 1.237061, 1.168793, 
    1.115082, 1.089691, 1.181274, 1.210571, 1.323273, 1.483429, 1.671326, 
    2.013763, 2.191162, 1.754944, 1.680176, 1.655121, 1.597321, 1.677704, 
    1.749115, 1.839417, 2.758301, 3.163574, 3.123474, 2.564728, 3.086304, 
    3.598846, 3.324036, 3.05896, 3.043121, 2.843109, 2.566711, 2.240906, 
    1.763977, 1.51358, 1.446045, 1.443451, 1.47934, 1.488068, 1.544189, 
    1.585144, 1.581665, 1.615448, 1.706238, 1.755829, 1.754791, 1.707855, 
    1.694733, 1.688446, 1.670593, 1.635834, 1.606171, 1.553223, 1.544769, 
    1.490967, 1.476807, 1.368988, 1.260468, 1.2229, 1.055054, 1.345947, 
    4.159607, 2.989197, 1.172302, 1.17334, 1.497101, 1.896759, 2.465057, 
    2.222748, 1.932129, 1.928619, 1.916046, 1.839081, 1.705414, 1.711426, 
    1.770721, 1.757904, 1.783478, 1.783112, 1.838104,
  1.744446, 1.698059, 1.768738, 1.812012, 2.115845, 3.965851, 4.133636, 
    3.609802, 3.146301, 2.29129, 2.146637, 2.230713, 2.214111, 2.160187, 
    2.013458, 1.942566, 1.956177, 1.892548, 1.798492, 1.768341, 1.829529, 
    1.897308, 1.995239, 2.082001, 2.138062, 2.225677, 2.366302, 2.432251, 
    2.291046, 1.85321, 1.811829, 3.148865, 2.94632, 2.715332, 3.058868, 
    3.116577, 3.303619, 3.599945, 3.630585, 3.401581, 3.179565, 2.305237, 
    2.026764, 2.192108, 2.410797, 2.536041, 2.249054, 1.739807, 1.546021, 
    1.470276, 1.445679, 1.526154, 1.591583, 1.623718, 1.657776, 1.679779, 
    1.70108, 1.760773, 1.767609, 1.796844, 1.771576, 1.716888, 1.681793, 
    1.601471, 1.590393, 1.528442, 1.420929, 1.332642, 1.279205, 1.259918, 
    1.188141, 1.181091, 1.119904, 1.087982, 1.032501, 0.9126892, 1.180817, 
    2.456085, 2.683441, 1.815063, 1.624969, 2.156403, 2.155121, 2.189026, 
    2.009796, 1.839539, 1.872284, 1.797424, 1.834991, 1.835327, 1.809174, 
    1.829071, 1.726532, 1.742676, 1.723206, 1.744568,
  1.562592, 1.526978, 1.676514, 1.772705, 2.357849, 3.891754, 3.886902, 
    3.715454, 3.2005, 2.370544, 2.294891, 2.514221, 2.471985, 2.335052, 
    2.467163, 2.517334, 2.545013, 2.469818, 2.412415, 2.414154, 2.341431, 
    2.341309, 2.316437, 2.286285, 2.2771, 2.200958, 2.094482, 1.950348, 
    1.86734, 1.80661, 2.063446, 3.732697, 4.009155, 3.631409, 3.575165, 
    3.11795, 3.427979, 3.988037, 4.21759, 4.075684, 3.634155, 1.64859, 
    1.333893, 1.577698, 1.828217, 1.965851, 1.951721, 1.906219, 1.900177, 
    1.928864, 1.934143, 1.857666, 1.819122, 1.765198, 1.694946, 1.604462, 
    1.550934, 1.567719, 1.57132, 1.568115, 1.539001, 1.45224, 1.36084, 
    1.240295, 1.226807, 1.221313, 1.230133, 1.190582, 1.169434, 1.171967, 
    1.101196, 1.136749, 1.124908, 1.042419, 0.8845825, 1.057068, 1.587738, 
    2.352966, 3.547485, 2.823395, 2.217804, 2.654114, 2.970856, 2.911957, 
    2.285736, 1.910065, 1.926971, 1.929657, 1.917267, 1.85318, 1.867493, 
    1.861816, 1.809631, 1.79541, 1.667999, 1.622375,
  1.633545, 1.756042, 1.96286, 2.363892, 3.807007, 3.585632, 3.24762, 
    3.386414, 3.745392, 3.443848, 2.397827, 2.548004, 3.424591, 2.357025, 
    2.262268, 2.415863, 2.268402, 2.258423, 2.171326, 2.102509, 2.062988, 
    2.045807, 2.044952, 2.041626, 2.047943, 1.985443, 1.929932, 1.890656, 
    1.964355, 2.055695, 2.27655, 4.112793, 4.276917, 3.952576, 4.045807, 
    3.484406, 3.564117, 4.005432, 3.874176, 3.503784, 2.802582, 1.690399, 
    1.845673, 2.037781, 2.07373, 2.103485, 2.051666, 2.088501, 1.992615, 
    1.901794, 1.834015, 1.692413, 1.618195, 1.501801, 1.437683, 1.441315, 
    1.442139, 1.467529, 1.459015, 1.399902, 1.348297, 1.30426, 1.329834, 
    1.287537, 1.297821, 1.298462, 1.30835, 1.277527, 1.243347, 1.200287, 
    1.18811, 1.18988, 1.014618, 1.000885, 1.036041, 1.542877, 2.400269, 
    3.357391, 4.607178, 3.475311, 2.674011, 3.160919, 3.075287, 3.185913, 
    3.454468, 2.269257, 1.95282, 1.969818, 1.916962, 1.816376, 1.768768, 
    1.69931, 1.597504, 1.53421, 1.499054, 1.56131,
  1.944244, 2.122437, 2.201782, 2.490265, 4.226685, 4.023926, 3.489624, 
    3.696136, 3.970459, 3.754272, 2.4711, 2.405212, 3.171112, 3.265076, 
    2.101074, 2.110382, 2.027527, 2.059418, 2.1008, 2.075012, 2.104584, 
    2.093262, 2.120728, 2.111237, 2.09729, 2.061432, 2.050385, 2.088318, 
    2.201935, 2.299072, 2.370544, 2.859863, 4.487915, 4.682922, 4.47464, 
    3.995667, 3.919891, 3.884155, 3.637512, 2.843475, 1.891632, 2.001801, 
    2.177917, 2.191101, 2.204987, 2.185699, 2.129578, 2.099518, 2.010376, 
    1.963013, 1.86142, 1.774963, 1.695435, 1.66037, 1.667358, 1.695862, 
    1.704895, 1.708252, 1.750671, 1.72757, 1.744751, 1.721069, 1.757904, 
    1.744843, 1.669037, 1.629578, 1.594818, 1.519348, 1.44516, 1.400177, 
    1.352905, 1.399902, 1.388885, 1.602051, 1.562988, 1.693146, 2.588806, 
    3.908173, 4.596954, 3.458801, 2.703796, 3.261871, 3.26416, 3.710602, 
    4.892548, 4.640533, 1.993469, 1.915314, 1.882019, 1.782196, 1.720398, 
    1.637604, 1.630219, 1.63147, 1.695099, 1.848145,
  2.293518, 2.388367, 2.416595, 2.528381, 4.506622, 4.425293, 3.706329, 
    3.728088, 4.128693, 4.49939, 3.729553, 2.341553, 2.968903, 3.579132, 
    2.096252, 2.100098, 2.145813, 2.192413, 2.251587, 2.28833, 2.319305, 
    2.298248, 2.277618, 2.285583, 2.304138, 2.296967, 2.317261, 2.410919, 
    2.504913, 2.52948, 2.488892, 2.548279, 2.837128, 4.146912, 4.055115, 
    3.914032, 3.754517, 2.408478, 2.937012, 2.02478, 2.060394, 2.238068, 
    2.255066, 2.247833, 2.237061, 2.207001, 2.230621, 2.237854, 2.213165, 
    2.151917, 2.060333, 1.98941, 1.978668, 2.018738, 2.055267, 2.136108, 
    2.201843, 2.230377, 2.263519, 2.255707, 2.25647, 2.21991, 2.186768, 
    2.157135, 2.082001, 2.04306, 1.945343, 1.927979, 1.888062, 1.901154, 
    1.886688, 1.953369, 1.962494, 1.995941, 1.966553, 2.330048, 3.974518, 
    4.31955, 4.08316, 3.189606, 2.721527, 3.269806, 3.556732, 3.165649, 
    4.786743, 4.708099, 1.849976, 1.93335, 1.927307, 1.867218, 1.915222, 
    1.901672, 2.024261, 2.101868, 2.190613, 2.27829,
  2.463226, 2.503998, 2.632477, 2.570953, 3.740662, 3.603546, 3.192871, 
    3.378143, 4.126343, 4.593109, 4.006866, 2.178955, 2.102356, 2.173431, 
    2.188232, 2.344574, 2.353729, 2.355286, 2.33252, 2.357788, 2.367615, 
    2.393982, 2.432922, 2.41983, 2.423401, 2.417419, 2.47879, 2.546387, 
    2.589539, 2.598083, 2.608887, 2.639984, 2.61554, 2.583679, 2.452698, 
    3.517609, 3.278687, 2.395538, 2.93811, 2.121185, 2.136871, 2.27478, 
    2.247559, 2.26709, 2.292175, 2.343384, 2.367432, 2.349731, 2.293274, 
    2.22464, 2.200104, 2.221588, 2.241425, 2.305115, 2.36911, 2.410492, 
    2.479614, 2.520538, 2.515656, 2.505676, 2.469849, 2.44455, 2.380707, 
    2.34137, 2.267456, 2.241699, 2.194427, 2.223145, 2.204041, 2.23584, 
    2.245392, 2.268921, 2.366577, 2.446136, 2.77417, 3.932526, 3.559265, 
    3.579926, 3.400818, 2.837402, 2.998718, 3.203278, 3.368378, 3.258118, 
    4.354218, 4.164124, 2.003357, 2.065521, 2.15094, 2.138824, 2.172821, 
    2.226715, 2.307709, 2.382568, 2.414429, 2.485107,
  2.564606, 2.617218, 2.70224, 2.47464, 3.937469, 3.636688, 3.002625, 
    2.929077, 3.163361, 4.209015, 3.696655, 2.207062, 2.27121, 2.370483, 
    2.462128, 2.522736, 2.504059, 2.526459, 2.41922, 2.437286, 2.423248, 
    2.421112, 2.422241, 2.459259, 2.503937, 2.534363, 2.54248, 2.547577, 
    2.472626, 2.52179, 2.519318, 2.568207, 2.536896, 2.537354, 2.458771, 
    2.388702, 2.345795, 2.493561, 3.227356, 2.210052, 2.196472, 2.315308, 
    2.300201, 2.30249, 2.270996, 2.269257, 2.274109, 2.25531, 2.204529, 
    2.196503, 2.231476, 2.266632, 2.335632, 2.409454, 2.468719, 2.539825, 
    2.555176, 2.595947, 2.60791, 2.593079, 2.553162, 2.529907, 2.475433, 
    2.451477, 2.410126, 2.405243, 2.401642, 2.406677, 2.445343, 2.487335, 
    2.50531, 2.54007, 2.670197, 2.707336, 2.738251, 3.128937, 3.258881, 
    3.593933, 3.448792, 3.162903, 2.904327, 2.968658, 3.085571, 3.677246, 
    3.630096, 3.88974, 3.75708, 2.291962, 2.384155, 2.402649, 2.364868, 
    2.463715, 2.450287, 2.51416, 2.534271, 2.562897,
  2.760315, 2.761505, 2.773651, 2.625092, 4.114441, 3.533966, 2.919952, 
    2.830017, 2.836029, 3.383362, 3.442352, 2.307892, 2.310394, 2.422455, 
    2.532257, 2.535858, 2.556366, 2.527374, 2.443604, 2.461945, 2.456604, 
    2.455414, 2.45578, 2.549255, 2.587402, 2.631409, 2.67868, 2.690063, 
    2.23114, 2.561737, 2.528748, 2.523865, 2.507843, 2.438904, 2.474976, 
    2.393646, 2.330719, 3.10434, 2.927399, 2.77417, 2.324005, 2.316193, 
    2.263763, 2.186493, 2.147247, 2.174683, 2.228699, 2.340576, 2.486084, 
    2.597687, 2.698151, 2.731812, 2.745819, 2.722382, 2.745148, 2.774719, 
    2.781677, 2.77771, 2.762604, 2.734985, 2.704071, 2.695801, 2.693909, 
    2.719818, 2.720978, 2.709717, 2.718079, 2.692108, 2.705109, 2.710602, 
    2.738586, 2.82547, 2.814697, 2.773621, 2.637268, 3.240997, 3.56839, 
    3.313263, 3.597961, 3.09317, 3.365143, 3.785004, 3.994995, 4.034271, 
    3.594391, 3.3591, 3.599518, 2.456146, 2.569122, 2.517151, 2.51767, 
    2.59079, 2.596497, 2.660522, 2.668274, 2.731079,
  2.693604, 2.686707, 2.658752, 2.934387, 3.358246, 3.047546, 2.932648, 
    3.023132, 2.745544, 2.257111, 2.572174, 3.359344, 2.409393, 2.396698, 
    2.471893, 2.459473, 2.428467, 2.376343, 2.39035, 2.401062, 2.417725, 
    2.396332, 2.429718, 2.526733, 2.598022, 2.655945, 2.610046, 2.704132, 
    2.341125, 2.499573, 2.468597, 2.716736, 2.75824, 2.260193, 2.342499, 
    2.94046, 3.055786, 2.817932, 2.643524, 2.362061, 2.349579, 2.271912, 
    2.261108, 2.228363, 2.341492, 2.505035, 2.754944, 3.137085, 3.388428, 
    3.418182, 3.399902, 3.332977, 3.286224, 3.284088, 3.268066, 3.221008, 
    3.170166, 3.116058, 3.071075, 3.009216, 2.976837, 2.96991, 3.013245, 
    3.025269, 3.044647, 3.00824, 2.968079, 2.940613, 2.879456, 2.855957, 
    2.790344, 2.71051, 2.51886, 2.370087, 2.218658, 3.125305, 3.587463, 
    3.351532, 3.48056, 3.699066, 3.944061, 5.122437, 4.052704, 3.615387, 
    3.374268, 2.507385, 2.538452, 2.533051, 2.617218, 2.597229, 2.654968, 
    2.592133, 2.635101, 2.675537, 2.682861, 2.709869,
  2.523346, 2.740997, 2.601074, 2.902191, 3.179382, 3.144562, 2.984985, 
    2.693085, 2.39859, 2.197815, 2.145935, 2.733368, 2.742218, 2.460754, 
    2.473419, 2.498474, 2.524384, 2.449524, 2.381409, 2.310455, 2.310638, 
    2.291046, 2.307068, 2.337402, 2.418243, 2.462982, 2.446381, 2.591675, 
    2.304382, 2.355804, 2.36853, 2.645355, 2.741974, 2.184479, 2.12561, 
    2.069458, 2.003357, 2.135376, 2.315704, 2.346893, 2.27179, 2.275482, 
    2.241241, 2.25824, 2.372192, 2.527435, 2.797699, 3.222382, 3.484863, 
    3.550629, 3.57605, 3.575684, 3.514099, 3.46756, 3.412537, 3.352112, 
    3.296143, 3.211365, 3.147614, 3.052826, 2.998871, 2.94873, 2.965912, 
    2.965332, 2.957123, 2.903229, 2.834015, 2.818329, 2.765778, 2.716766, 
    2.60968, 2.488953, 2.272156, 2.045288, 1.841187, 2.842224, 3.915283, 
    3.712921, 3.573059, 4.145996, 4.577576, 3.969635, 3.597107, 2.407013, 
    2.41748, 2.3591, 2.430389, 2.402313, 2.407135, 2.438782, 2.471069, 
    2.440979, 2.540771, 2.521057, 2.550354, 2.455627,
  3.000061, 2.900879, 3.048462, 3.321594, 3.349365, 3.227417, 3.036621, 
    2.599823, 2.559418, 2.671265, 2.634003, 2.698883, 2.285461, 2.349243, 
    2.396973, 2.462769, 2.55249, 2.593781, 2.548981, 2.50528, 2.428864, 
    2.384735, 2.301666, 2.295288, 2.327484, 2.325226, 2.916504, 2.819824, 
    2.320465, 2.277069, 2.286682, 2.865479, 2.167603, 2.246704, 2.261688, 
    2.152557, 2.144379, 2.251312, 2.303345, 2.289093, 2.276733, 2.274445, 
    2.174774, 2.107452, 2.082581, 2.118317, 2.246246, 2.355499, 2.515869, 
    2.672943, 2.77652, 2.859406, 2.885986, 2.922424, 2.956665, 2.925293, 
    2.867798, 2.77063, 2.680176, 2.621826, 2.567535, 2.52478, 2.510773, 
    2.527893, 2.493011, 2.535889, 2.517548, 2.532257, 2.592804, 2.608429, 
    2.626709, 2.47757, 2.292938, 2.210114, 2.216248, 3.251648, 3.656616, 
    3.696075, 4.179993, 4.865967, 3.557861, 3.046234, 2.620544, 2.493011, 
    2.481567, 2.468842, 2.438507, 2.410187, 2.440979, 2.392792, 2.40799, 
    2.421112, 2.448547, 2.419769, 3.009003, 2.966614,
  3.39325, 3.162262, 3.41626, 3.704803, 3.922638, 3.851532, 3.234741, 
    3.201141, 3.031921, 2.963745, 3.026855, 2.825012, 2.272278, 1.883301, 
    2.398865, 2.453033, 2.573395, 2.546387, 2.489227, 2.40271, 2.423279, 
    2.747162, 2.467865, 2.319305, 2.296051, 2.16864, 2.17868, 2.992737, 
    2.385071, 2.315094, 2.283966, 2.315674, 2.337494, 2.845215, 2.302246, 
    2.268188, 2.306915, 2.263184, 2.26767, 2.266174, 2.26181, 2.251465, 
    2.173187, 2.115204, 2.111755, 2.177368, 2.170807, 2.135254, 2.177643, 
    2.223663, 2.219116, 2.222778, 2.238647, 2.29718, 2.353882, 2.371368, 
    2.329407, 2.278442, 2.239288, 2.276093, 2.289551, 2.353546, 2.420288, 
    2.506104, 2.52829, 2.612732, 2.673798, 2.698792, 2.69104, 2.686035, 
    2.66272, 2.560425, 2.76767, 2.796326, 3.331482, 3.457794, 3.430237, 
    3.997772, 4.341553, 3.781128, 2.314758, 2.362946, 2.348663, 2.382843, 
    2.390472, 2.371765, 2.395203, 2.442657, 2.482361, 2.439697, 2.42868, 
    2.329376, 2.443268, 3.33786, 3.357117, 3.393707,
  3.786316, 3.412415, 3.115936, 2.893005, 3.344574, 3.79599, 3.975616, 
    4.700165, 3.993256, 4.261353, 4.10675, 4.422882, 3.331116, 2.918457, 
    2.471313, 2.46521, 2.537262, 2.478546, 2.435577, 2.367157, 3.106293, 
    3.124329, 2.473724, 2.438507, 2.376831, 2.163574, 1.940155, 2.680878, 
    2.643188, 2.586212, 2.308472, 2.366241, 2.3508, 2.730499, 2.22406, 
    2.221588, 2.245941, 2.231628, 2.234161, 2.244873, 2.276123, 2.266205, 
    2.216919, 2.221832, 2.238068, 2.275055, 2.264618, 2.295929, 2.377777, 
    2.446899, 2.458038, 2.449524, 2.424438, 2.445526, 2.43573, 2.43631, 
    2.389221, 2.374847, 2.353882, 2.354462, 2.365204, 2.424316, 2.472229, 
    2.504456, 2.528168, 2.634583, 2.772705, 2.861359, 2.740997, 2.701721, 
    2.700623, 2.875092, 3.929932, 3.723938, 2.383606, 2.288788, 2.189026, 
    2.17157, 2.197174, 2.293335, 2.305115, 2.334473, 2.290802, 2.279144, 
    2.215271, 2.287933, 2.281067, 2.326935, 2.385498, 2.489014, 2.448212, 
    2.472961, 4.138428, 4.375244, 4.1492, 3.532257,
  3.737854, 3.505249, 3.045197, 2.99118, 3.088501, 3.005493, 3.145355, 
    2.998291, 3.059418, 3.535919, 3.997437, 4.466095, 3.509338, 3.118256, 
    2.610382, 2.448151, 2.479706, 2.473083, 2.443726, 2.462463, 3.681061, 
    3.656799, 2.619232, 2.601471, 2.359863, 2.199585, 2.880615, 2.633545, 
    2.02594, 1.925568, 2.248657, 2.382904, 2.298157, 2.103699, 2.222168, 
    2.215607, 2.188965, 2.239655, 2.267609, 2.256958, 2.257599, 2.239868, 
    2.218445, 2.248016, 2.27652, 2.308502, 2.347839, 2.383698, 2.423859, 
    2.416809, 2.406677, 2.386902, 2.358307, 2.366302, 2.354462, 2.360199, 
    2.363098, 2.377777, 2.359253, 2.331207, 2.285004, 2.228271, 2.188812, 
    2.195801, 2.28299, 2.522949, 2.711945, 2.680176, 2.609222, 3.493927, 
    3.84549, 4.183563, 4.023285, 2.338562, 2.390259, 2.353027, 2.286224, 
    2.303741, 2.276398, 2.323669, 2.2547, 2.237671, 2.208252, 2.185699, 
    2.152832, 2.172424, 2.132904, 2.230957, 2.27771, 2.426788, 2.403961, 
    2.540985, 3.990448, 3.9505, 3.684814, 3.482849,
  3.436737, 3.213623, 3.070343, 2.930359, 2.904114, 3.00882, 3.108887, 
    3.019714, 3.165009, 3.154419, 2.682465, 4.093842, 4.043274, 4.456421, 
    4.244263, 3.235138, 2.331665, 2.418701, 2.533905, 2.487335, 3.748901, 
    3.667419, 3.788055, 3.477173, 2.416565, 2.845734, 3.040009, 2.381531, 
    1.924103, 2.003235, 2.04599, 2.261688, 2.317108, 2.187195, 2.247925, 
    2.290466, 2.244812, 2.207336, 2.185242, 2.201141, 2.227966, 2.203369, 
    2.226593, 2.256805, 2.291626, 2.342346, 2.374146, 2.375305, 2.370667, 
    2.376617, 2.364014, 2.376404, 2.362885, 2.328339, 2.321381, 2.311371, 
    2.326599, 2.322357, 2.314545, 2.300293, 2.256683, 2.126312, 1.959991, 
    1.844055, 1.869629, 2.079895, 2.438904, 2.669708, 3.37561, 3.498993, 
    3.864929, 4.159027, 3.971405, 2.29657, 2.402557, 2.38324, 2.294434, 
    2.345032, 2.315521, 2.284943, 2.243256, 2.273102, 2.239166, 2.186768, 
    2.092224, 2.049652, 2.053345, 2.071259, 2.021576, 2.153564, 2.202942, 
    2.56546, 4.05426, 3.9823, 3.822174, 3.814728,
  3.977753, 3.629395, 3.072235, 2.929138, 2.727692, 2.468872, 2.685852, 
    3.062805, 3.420074, 3.616058, 2.878296, 4.475616, 4.246643, 4.617889, 
    4.806305, 4.107635, 2.516418, 2.659943, 3.514862, 3.097382, 3.080017, 
    3.314484, 3.066345, 3.226135, 2.96228, 3.216034, 3.243866, 2.55072, 
    1.740601, 2.032898, 2.184479, 1.957245, 2.148071, 2.231873, 2.240967, 
    2.301788, 2.291565, 2.207642, 2.156799, 2.151123, 2.169769, 2.18219, 
    2.220337, 2.224396, 2.279541, 2.329254, 2.356415, 2.363708, 2.358063, 
    2.382263, 2.334839, 2.284363, 2.233246, 2.173401, 2.189667, 2.173279, 
    2.159088, 2.133118, 2.142609, 2.138184, 2.143158, 2.070526, 1.953156, 
    1.794373, 1.700562, 1.774719, 2.312744, 4.006195, 4.030304, 3.635895, 
    3.756042, 2.546326, 2.302704, 2.386414, 2.433563, 2.359344, 2.298737, 
    2.371185, 2.421509, 2.435516, 2.393127, 2.357697, 2.318634, 2.290344, 
    2.21344, 2.200073, 2.136902, 2.071716, 2.064087, 2.024902, 1.929718, 
    2.423859, 4.364624, 4.696381, 4.50354, 4.178223,
  3.969238, 3.699066, 3.123199, 3.044373, 3.069092, 2.790924, 3.259613, 
    3.305115, 3.400085, 3.584229, 4.124451, 4.099823, 3.898804, 4.26593, 
    4.536957, 4.135468, 4.163391, 4.312897, 4.292542, 3.593475, 3.008942, 
    3.223907, 3.445984, 2.907593, 2.904663, 2.790344, 3.022247, 2.767944, 
    1.989044, 1.724335, 1.711578, 1.605194, 1.813507, 2.19165, 2.170044, 
    2.205109, 2.29953, 2.355164, 2.296326, 2.203491, 2.160645, 2.165375, 
    2.220459, 2.240387, 2.245422, 2.26593, 2.262573, 2.269104, 2.279388, 
    2.309082, 2.364685, 2.391235, 2.373413, 2.327118, 2.279541, 2.231232, 
    2.170471, 2.120148, 2.085449, 2.111816, 2.088043, 2.025665, 1.943726, 
    1.782257, 1.696899, 1.94812, 3.577637, 4.098206, 3.926819, 3.341064, 
    3.442688, 2.77594, 2.835663, 2.927032, 3.309601, 2.372375, 2.306549, 
    2.337799, 2.402832, 2.386108, 2.349976, 2.328033, 2.32959, 2.324249, 
    2.301544, 2.27829, 2.241913, 2.249634, 2.194763, 2.078918, 1.970734, 
    1.996582, 2.437469, 4.195282, 4.396454, 3.937805,
  3.375092, 3.592407, 3.299194, 3.317596, 3.179199, 2.387665, 3.12262, 
    3.166382, 2.426575, 3.453278, 3.580566, 3.697479, 3.91391, 4.277191, 
    4.247375, 3.804199, 3.885193, 4.250214, 4.282318, 4.270782, 4.093781, 
    3.999451, 3.74353, 3.464233, 3.37854, 2.695862, 2.334015, 2.853363, 
    2.98056, 2.670258, 2.272888, 1.884277, 1.806213, 1.946472, 2.047119, 
    2.236603, 2.383606, 2.439362, 2.41684, 2.302856, 2.218842, 2.135315, 
    2.138824, 2.150513, 2.178009, 2.214539, 2.243256, 2.256409, 2.297485, 
    2.34137, 2.386383, 2.387268, 2.419312, 2.463165, 2.461243, 2.422028, 
    2.324768, 2.236176, 2.11853, 2.086884, 2.002045, 1.926117, 1.904846, 
    1.883301, 1.973999, 3.084076, 3.573456, 3.520996, 3.35379, 3.109802, 
    3.145996, 3.634125, 4.179901, 4.188446, 3.743988, 2.502014, 2.316376, 
    2.212189, 2.215118, 2.234283, 2.296051, 2.276184, 2.22641, 2.202515, 
    2.197296, 2.180237, 2.225555, 2.320526, 2.337463, 2.30191, 2.223999, 
    2.026276, 2.100372, 2.620544, 4.170288, 3.427155,
  3.399841, 3.387512, 3.239624, 2.789917, 2.591156, 2.374847, 2.125397, 
    2.14743, 2.40686, 2.584564, 2.957642, 3.479584, 3.759277, 3.972748, 
    3.890137, 3.731873, 3.61026, 3.779266, 3.710022, 4.028961, 3.60025, 
    4.065796, 3.342621, 3.721832, 3.568695, 3.164734, 2.207977, 2.754944, 
    3.441315, 3.601471, 2.442322, 2.032074, 1.953796, 2.027679, 2.290192, 
    2.201202, 2.849701, 2.93277, 2.525421, 2.463196, 2.361176, 2.274902, 
    2.246887, 2.202393, 2.142334, 2.120819, 2.175232, 2.253204, 2.311401, 
    2.375336, 2.424194, 2.469025, 2.537262, 2.568848, 2.571655, 2.581665, 
    2.473267, 2.329315, 2.231537, 2.15094, 2.043213, 1.931549, 1.918121, 
    1.990845, 2.554932, 2.776672, 2.837982, 2.898468, 3.210358, 3.250946, 
    2.727631, 3.035492, 3.575104, 3.710327, 3.571136, 3.459595, 2.671844, 
    2.398804, 2.204224, 2.134888, 2.063843, 2.021759, 2.122101, 2.156555, 
    2.079803, 2.036163, 1.996796, 2.148621, 2.402313, 2.504852, 2.398651, 
    2.220367, 2.055695, 2.200104, 2.637909, 2.950867,
  2.70401, 2.793549, 2.762787, 2.641479, 2.573425, 2.564209, 3.126526, 
    2.849976, 2.82431, 2.691559, 2.49054, 2.786896, 3.064026, 3.028076, 
    2.376465, 3.129333, 3.285767, 3.512329, 3.434418, 4.228333, 4.794891, 
    3.402588, 2.86377, 2.931427, 3.644379, 2.783173, 2.935822, 1.959137, 
    1.900055, 2.098938, 2.176331, 2.337189, 1.920563, 2.127441, 2.006622, 
    2.437653, 2.566101, 2.895935, 2.495789, 2.50296, 2.478027, 2.466644, 
    2.507782, 2.583893, 2.617615, 2.530579, 2.432343, 2.431915, 2.4758, 
    2.513428, 2.504852, 2.498413, 2.544708, 2.555603, 2.522827, 2.510315, 
    2.444061, 2.397186, 2.326508, 2.199585, 2.022491, 1.84613, 1.889526, 
    2.155548, 2.159424, 1.981049, 2.191254, 2.10968, 2.296204, 2.618591, 
    2.556671, 2.764038, 3.058105, 3.264038, 3.41095, 3.452759, 3.396912, 
    3.099823, 2.797028, 2.522888, 2.212189, 2.035706, 2.199768, 2.272491, 
    2.127563, 1.947418, 1.748596, 1.686218, 1.958099, 2.267426, 2.430695, 
    2.331146, 2.096863, 2.162781, 2.517181, 2.7341,
  2.689423, 2.552643, 2.661102, 2.627991, 2.704498, 2.975677, 3.638, 
    3.264282, 3.101013, 2.907867, 3.086548, 3.004211, 2.871765, 2.368835, 
    2.946564, 3.183319, 3.114105, 2.847626, 2.784943, 3.143982, 3.465332, 
    3.191467, 3.082672, 3.026398, 3.198822, 3.32489, 3.664215, 3.242279, 
    2.910828, 2.441376, 2.220551, 2.125336, 2.023804, 2.082642, 2.334137, 
    2.346527, 2.628998, 2.723541, 2.914886, 3.074524, 2.815735, 2.700165, 
    2.553345, 2.446106, 2.424316, 2.43219, 2.442688, 2.424713, 2.405304, 
    2.41983, 2.454987, 2.514008, 2.565063, 2.573456, 2.515137, 2.408691, 
    2.314758, 2.264343, 2.212677, 2.166718, 2.098816, 1.932922, 1.870087, 
    1.969604, 2.00769, 2.011322, 1.972687, 1.512024, 1.625122, 2.098602, 
    2.272675, 2.187744, 2.471252, 2.936859, 3.205627, 3.071198, 3.084564, 
    3.206421, 3.291962, 3.128082, 2.770996, 2.50119, 2.509735, 2.247925, 
    1.994293, 1.82254, 1.571625, 1.327515, 1.46814, 1.789185, 2.101135, 
    2.198059, 2.057007, 2.097626, 2.507019, 2.680237,
  2.668915, 2.345001, 2.242218, 2.499969, 2.486572, 2.709717, 3.184692, 
    2.973602, 2.983948, 3.009155, 2.854401, 2.733948, 2.577759, 2.598267, 
    2.21051, 2.545868, 2.539703, 2.541199, 2.536896, 2.541199, 2.720612, 
    3.222229, 3.982971, 4.173401, 4.505829, 4.625488, 4.627502, 4.237274, 
    3.422119, 2.940125, 2.88089, 2.833771, 2.861481, 3.050812, 3.11795, 
    3.079071, 3.215332, 2.896759, 2.898865, 2.706268, 2.514923, 2.475616, 
    2.389343, 2.274963, 2.199768, 2.215668, 2.275421, 2.324524, 2.357971, 
    2.408295, 2.457123, 2.450806, 2.449646, 2.473541, 2.491638, 2.48468, 
    2.457184, 2.385895, 2.290527, 2.178741, 2.058167, 1.907318, 1.879456, 
    1.886536, 2.124176, 2.117798, 1.813721, 1.68335, 1.85083, 2.031677, 
    2.004669, 2.106628, 2.333466, 3.062012, 2.930756, 3.106476, 3.197571, 
    3.362274, 3.365936, 3.344177, 3.098267, 2.69397, 2.036499, 1.801453, 
    1.813232, 1.740387, 1.458649, 1.0961, 1.013, 1.264221, 1.565521, 
    1.879974, 1.948669, 1.929596, 2.067749, 2.555634,
  2.125549, 2.339569, 2.454498, 2.463501, 2.243256, 2.269623, 2.426208, 
    2.423737, 2.634857, 2.600372, 2.513641, 2.483459, 2.389099, 2.44751, 
    2.345367, 2.194885, 2.008942, 2.143982, 2.280823, 2.204407, 2.366821, 
    2.755371, 3.341766, 3.392883, 3.58313, 3.523346, 3.430969, 3.244324, 
    3.558563, 4.279388, 3.827118, 4.30426, 4.566895, 4.659393, 4.837921, 
    4.845947, 5.121979, 4.713196, 2.675079, 2.432526, 2.484985, 2.483887, 
    2.446228, 2.268127, 2.157318, 2.181671, 2.22644, 2.278351, 2.343994, 
    2.390198, 2.420166, 2.462341, 2.566498, 2.667542, 2.699982, 2.655365, 
    2.574432, 2.467987, 2.357697, 2.222168, 2.045685, 1.956421, 2.208832, 
    2.539307, 3.009491, 2.541565, 2.048553, 1.875244, 2.014893, 2.301361, 
    2.539307, 2.630249, 2.824463, 2.88797, 3.040009, 3.363525, 3.68689, 
    3.918579, 4.205048, 3.971985, 3.252258, 3.082916, 2.29834, 2.068329, 
    1.855896, 1.568237, 1.080444, 0.4162292, 0.07055664, 0.2893677, 
    0.8170776, 1.330048, 1.558441, 1.573456, 1.685791, 1.945862,
  1.565582, 1.870544, 2.419159, 2.548035, 2.37027, 2.38382, 2.605103, 
    2.569519, 2.432159, 2.368591, 2.330048, 2.370605, 2.462921, 2.36554, 
    2.584351, 2.671783, 2.451843, 2.353333, 2.445984, 2.424591, 2.490387, 
    2.992798, 3.568329, 3.782379, 3.906342, 3.706482, 4.063049, 4.190369, 
    4.351135, 4.59053, 3.930115, 4.196976, 4.914734, 5.986938, 5.510834, 
    5.441315, 5.670364, 4.931152, 2.557526, 2.220734, 2.327515, 2.459412, 
    2.5914, 2.089294, 2.040131, 2.208313, 2.301453, 2.416565, 2.506409, 
    2.536316, 2.561127, 2.657471, 2.798798, 2.890198, 2.838837, 2.752594, 
    2.68219, 2.550354, 2.378418, 2.23819, 2.113464, 2.61676, 3.113708, 
    3.414307, 2.982178, 2.540771, 2.325104, 2.659607, 3.003021, 3.076935, 
    3.210815, 3.572235, 3.566376, 3.507874, 3.497681, 3.6492, 4.666199, 
    5.251801, 5.73349, 5.50412, 4.545471, 2.574036, 2.131805, 1.730225, 
    1.562134, 1.543976, 1.226196, 0.5753174, -0.009033203, -0.0425415, 
    0.4301147, 0.9837036, 1.265411, 1.379059, 1.454651, 1.486145,
  1.280548, 1.624176, 1.638885, 1.927185, 1.899628, 2.054993, 2.055298, 
    2.421722, 2.616302, 2.736084, 2.643524, 2.69928, 2.78299, 2.967926, 
    3.113922, 3.38855, 3.469696, 3.572113, 3.46701, 3.474121, 3.562866, 
    3.836639, 4.300232, 4.348785, 4.324951, 4.265198, 4.533386, 5.04364, 
    5.638596, 5.074646, 4.864182, 5.030533, 5.049194, 5.149078, 5.384811, 
    5.557083, 5.515015, 4.727264, 2.511261, 2.293213, 2.452087, 2.621735, 
    3.534424, 3.344635, 2.401154, 2.649261, 2.722046, 2.695404, 2.869781, 
    3.052246, 3.200104, 3.299957, 3.308167, 3.3172, 3.429413, 2.792694, 
    2.657135, 2.553894, 2.47049, 2.404388, 3.259216, 4.160461, 4.216766, 
    3.87262, 3.135193, 2.686554, 2.617035, 3.403473, 3.902893, 4.259979, 
    4.146515, 4.206085, 3.542816, 3.564056, 3.789429, 4.277527, 5.935455, 
    6.257965, 6.409729, 5.723022, 2.575897, 2.03833, 1.686829, 1.588104, 
    1.700104, 1.613708, 1.565674, 1.242859, 0.777771, 0.6105347, 0.7743835, 
    1.015656, 1.168976, 1.248535, 1.29541, 1.455627,
  1.18161, 1.513977, 1.4245, 2.115631, 2.265594, 1.768768, 1.809082, 
    1.751007, 1.932922, 2.172028, 2.565704, 3.058807, 3.511566, 3.862854, 
    4.139923, 4.210449, 4.507904, 4.578674, 4.649048, 4.864136, 5.202179, 
    5.466675, 5.569183, 5.43988, 5.257523, 5.247559, 5.635391, 6.022934, 
    6.307571, 5.938126, 6.239624, 6.368805, 6.734238, 6.926926, 7.406693, 
    7.224258, 6.380722, 5.184891, 4.898087, 4.871979, 5.394379, 5.14061, 
    5.150116, 5.50708, 5.305969, 4.91507, 4.839996, 3.350159, 3.861938, 
    4.218536, 4.222107, 4.02536, 5.210754, 5.537872, 5.792816, 5.731018, 
    5.60025, 5.104767, 4.636688, 4.467102, 4.70752, 4.765686, 4.587524, 
    3.869873, 3.531555, 3.495239, 4.005371, 4.821533, 5.194, 5.368011, 
    5.383514, 4.029022, 4.391418, 4.888, 5.856018, 6.487488, 7.56665, 
    7.688263, 6.352722, 4.344818, 2.520111, 1.917816, 1.645294, 1.591827, 
    2.717834, 1.279327, 1.507568, 1.399506, 1.36084, 1.319244, 1.253937, 
    1.111938, 0.875946, 0.7355042, 0.918457, 1.055298,
  0.8235168, 0.8989868, 0.8092957, 1.092346, 1.214233, 1.381958, 1.479645, 
    2.087006, 2.440216, 2.834412, 3.213043, 3.549988, 3.914551, 4.327118, 
    4.655945, 5.035461, 5.263794, 5.410187, 5.651215, 6.006226, 6.456482, 
    6.719955, 6.676529, 6.473236, 6.156433, 5.699539, 5.512039, 5.553375, 
    5.819321, 7.510269, 7.380905, 7.093658, 7.416382, 8.195694, 7.622437, 
    6.868469, 5.088989, 5.404221, 5.566071, 5.426086, 5.697968, 5.600769, 
    5.863525, 5.853165, 5.711182, 5.774063, 6.985275, 7.730621, 9.246643, 
    10.36168, 10.22147, 6.739044, 7.101135, 6.063446, 5.482758, 5.12793, 
    4.793671, 4.553833, 4.3078, 4.435913, 4.463409, 4.509277, 4.429291, 
    4.123413, 3.934814, 4.169434, 4.683777, 5.520752, 6.322433, 7.165726, 
    7.59758, 8.056503, 8.852112, 9.979538, 11.91638, 11.86896, 11.55322, 
    9.944244, 8.628998, 7.11377, 3.798645, 2.626007, 3.870087, 3.374908, 
    2.995483, 2.503387, 2.162872, 0.970459, 0.9671631, 0.8794556, 0.9573669, 
    1.285187, 0.9101868, 0.6324158, 0.6018982, 0.6486816,
  0.942749, 0.8336792, 0.7754211, 0.8567505, 0.9456787, 1.396515, 1.905701, 
    2.403198, 2.721771, 2.899994, 2.96286, 1.946625, 2.074066, 2.435852, 
    4.6604, 6.027374, 6.966705, 7.522049, 7.820023, 7.732651, 7.534088, 
    7.394592, 7.356308, 7.359161, 7.307938, 6.477066, 6.499786, 6.995682, 
    7.071915, 6.921799, 6.907272, 6.784042, 6.848221, 6.668213, 5.792496, 
    6.006042, 7.412537, 6.602203, 7.833389, 8.503952, 8.843933, 8.553116, 
    8.637421, 8.443085, 6.760452, 6.485931, 6.634811, 7.86261, 9.799789, 
    15.5941, 16.79744, 14.63214, 13.11435, 9.240921, 7.96489, 7.448471, 
    7.308182, 7.12381, 6.269775, 6.913773, 6.717819, 6.411636, 6.184357, 
    5.900314, 6.191528, 6.284866, 6.709366, 7.626633, 8.469238, 8.707886, 
    9.500702, 9.389572, 9.814224, 11.88016, 11.11833, 11.53563, 11.79295, 
    11.33324, 10.15485, 9.42392, 6.458771, 4.359039, 4.438049, 3.958786, 
    3.619644, 3.827011, 3.560791, 3.348755, 3.360855, 3.471466, 3.721649, 
    3.269928, 2.41684, 2.153381, 1.569763, 1.179657,
  2.170471, 1.707581, 1.369232, 1.187408, 1.051422, 1.156494, 1.656891, 
    2.254578, 2.59491, 2.691376, 2.65509, 2.624329, 2.930267, 4.302704, 
    6.528564, 9.233643, 11.71326, 12.55739, 12.41704, 9.748611, 8.936264, 
    8.382217, 8.319458, 7.892105, 7.412872, 6.88768, 6.617569, 6.492569, 
    6.492035, 6.853897, 6.437943, 6.792313, 7.30838, 8.080261, 8.983444, 
    10.19205, 11.01099, 11.44667, 8.799271, 8.291916, 9.773819, 9.791641, 
    9.655457, 9.555771, 9.236374, 8.633377, 8.093475, 8.04158, 8.602722, 
    9.532608, 10.29431, 10.43214, 10.30325, 10.03799, 9.788071, 9.754593, 
    9.868271, 9.972763, 9.902771, 9.583725, 9.107742, 8.392303, 7.346924, 
    6.672958, 6.405777, 6.448883, 6.972656, 7.814896, 8.729034, 11.24026, 
    9.895432, 10.01015, 11.98418, 9.514297, 9.87941, 10.27071, 11.19518, 
    13.258, 13.3488, 11.63602, 8.703613, 6.668137, 5.30513, 4.038651, 
    3.201096, 2.789566, 2.417236, 2.780518, 3.678757, 4.844193, 6.13826, 
    9.13356, 9.039673, 6.936157, 3.829254, 2.685486,
  4.187805, 2.371674, 2.179535, 2.163513, 1.987427, 2.50116, 3.943604, 
    5.945404, 7.540588, 8.484283, 9.314423, 9.973297, 10.67368, 11.24445, 
    11.416, 11.6833, 12.00807, 12.07166, 11.79756, 11.34256, 10.65195, 
    9.882736, 9.296143, 8.643982, 7.847427, 8.047379, 7.901413, 7.694122, 
    7.622894, 7.868271, 7.753632, 7.95813, 8.376999, 8.82283, 9.020355, 
    8.988663, 8.897125, 8.555649, 7.968811, 7.649582, 7.575439, 7.629944, 
    7.765228, 7.935471, 8.068542, 8.081955, 7.933578, 7.809875, 7.73996, 
    7.734558, 7.837753, 8.071533, 8.332794, 8.519714, 8.650314, 8.682922, 
    8.671005, 8.667572, 8.627716, 8.613922, 8.585342, 8.47699, 8.243149, 
    7.996414, 7.49086, 7.520294, 7.578308, 7.591324, 7.679276, 7.944138, 
    8.188004, 8.896133, 8.707077, 8.705841, 8.619507, 9.022293, 9.554276, 
    9.329163, 7.82283, 6.947189, 5.966583, 5.221008, 4.64537, 4.309875, 
    4.119385, 3.681427, 3.308838, 3.380127, 3.929596, 4.760651, 5.691589, 
    6.388916, 7.189774, 7.622833, 7.490265, 6.836639,
  6.376297, 6.108109, 5.739105, 5.272614, 5.708694, 5.886185, 6.162735, 
    6.780762, 7.294388, 7.654068, 7.941116, 8.168137, 8.354858, 8.449448, 
    8.443283, 8.3806, 8.328384, 8.242905, 8.18071, 8.173431, 8.114487, 
    8.067566, 7.996597, 7.864883, 7.611313, 7.784683, 7.784683, 7.570282, 
    7.658768, 7.678436, 7.651352, 7.600311, 7.637939, 7.667557, 7.613266, 
    7.545486, 7.470367, 7.374191, 7.249069, 7.14035, 7.086899, 7.07811, 
    7.025894, 7.021011, 7.054214, 7.15506, 7.254272, 7.38266, 7.541321, 
    7.658829, 7.773285, 7.862625, 7.90831, 7.925644, 7.882339, 7.811951, 
    7.717163, 7.62915, 7.581436, 7.629471, 7.726547, 7.879074, 7.990738, 
    8.10318, 8.191132, 8.20578, 8.226929, 8.127655, 7.862549, 7.774002, 
    7.601486, 6.908188, 6.956497, 7.122894, 7.034225, 6.889435, 6.689117, 
    6.414246, 6.150177, 5.871597, 5.578629, 5.268799, 5.001495, 4.801422, 
    4.650513, 4.534622, 4.469589, 4.707794, 5.049393, 5.493469, 5.793991, 
    6.098419, 6.772049, 6.85701, 6.879791, 6.733261,
  6.43103, 6.326752, 6.327988, 6.328308, 6.303177, 6.347961, 6.352844, 
    6.450241, 6.543594, 6.628891, 6.728439, 6.801422, 6.861237, 6.913132, 
    6.95488, 6.95961, 6.95903, 6.98703, 7.015869, 7.056824, 7.077652, 
    7.082336, 7.06163, 7.05629, 7.083771, 7.060532, 7.127655, 7.085068, 
    7.138077, 7.210922, 7.291916, 7.350372, 7.403488, 7.453949, 7.539886, 
    7.579147, 7.543076, 7.503174, 7.480194, 7.474991, 7.449921, 7.43103, 
    7.406174, 7.326935, 7.249924, 7.185913, 7.128693, 7.093155, 7.046402, 
    7.011963, 6.938522, 6.881638, 6.883957, 6.8992, 6.964767, 7.016769, 
    7.011307, 7.091324, 7.223679, 7.358826, 7.520554, 7.697433, 7.795822, 
    7.871658, 7.91925, 7.904541, 7.889175, 7.845047, 7.839691, 7.840347, 
    7.831619, 7.820099, 7.848434, 7.960663, 7.956039, 7.948349, 7.954086, 
    8.147308, 8.336319, 8.327515, 8.292435, 8.179672, 8.053955, 7.884094, 
    7.990479, 8.10759, 8.173431, 8.090347, 8.101349, 7.832077, 7.715546, 
    7.594055, 7.223816, 6.929611, 6.70285, 6.575363,
  6.631561, 6.507019, 6.496216, 6.503036, 6.495483, 6.55571, 6.566452, 
    6.554932, 6.545166, 6.564499, 6.552002, 6.545547, 6.560272, 6.575897, 
    6.572189, 6.556488, 6.505127, 6.452271, 6.425308, 6.432999, 6.455261, 
    6.491852, 6.520035, 6.539963, 6.557938, 6.557343, 6.567307, 6.581879, 
    6.579468, 6.57283, 6.593079, 6.638657, 6.668335, 6.719788, 6.753311, 
    6.793213, 6.815353, 6.852066, 6.882019, 6.91835, 6.92485, 6.943405, 
    6.954025, 6.962494, 6.970947, 6.95285, 6.937347, 6.951294, 6.97316, 
    6.974274, 7.003174, 6.982407, 6.988083, 7.000702, 7.020172, 7.047714, 
    7.140945, 7.183701, 7.24205, 7.273743, 7.299194, 7.37999, 7.426147, 
    7.502197, 7.551865, 7.579605, 7.61673, 7.594513, 7.569199, 7.574188, 
    7.576096, 7.5867, 7.577393, 7.575378, 7.627975, 7.646011, 7.676086, 
    7.696533, 7.715088, 7.727203, 7.728104, 7.708374, 7.661896, 7.604874, 
    7.538147, 7.48494, 7.431808, 7.395233, 7.365021, 7.306824, 7.207596, 
    7.085785, 6.98085, 6.852066, 6.733582, 6.668289,
  1.718872, 1.701111, 1.689835, 1.67662, 1.666412, 1.651489, 1.641479, 
    1.634705, 1.630539, 1.62175, 1.609634, 1.598373, 1.595963, 1.601044, 
    1.607285, 1.611465, 1.621689, 1.630341, 1.636124, 1.644272, 1.652206, 
    1.661911, 1.66745, 1.675262, 1.681503, 1.682617, 1.682419, 1.67955, 
    1.669861, 1.662766, 1.647903, 1.633652, 1.620636, 1.611389, 1.598694, 
    1.584839, 1.574478, 1.563278, 1.543488, 1.523895, 1.508469, 1.492065, 
    1.474869, 1.464005, 1.458282, 1.458725, 1.455917, 1.462097, 1.4608, 
    1.474609, 1.490356, 1.509064, 1.531784, 1.525528, 1.5457, 1.569016, 
    1.59375, 1.609497, 1.615692, 1.627213, 1.633469, 1.650391, 1.677155, 
    1.691269, 1.710602, 1.728912, 1.746948, 1.773895, 1.804291, 1.8293, 
    1.850067, 1.866791, 1.882416, 1.910278, 1.916214, 1.929489, 1.944412, 
    1.965286, 1.962891, 1.97226, 1.981842, 1.979553, 1.9776, 1.979294, 
    1.971817, 1.967651, 1.955017, 1.941864, 1.919724, 1.894852, 1.865372, 
    1.833008, 1.802872, 1.78067, 1.75592, 1.737366,
  1.891739, 1.885681, 1.87233, 1.837692, 1.794464, 1.760925, 1.739334, 
    1.733994, 1.734634, 1.730347, 1.713745, 1.692123, 1.665237, 1.654434, 
    1.650711, 1.652863, 1.681183, 1.725327, 1.77655, 1.828903, 1.874619, 
    1.905273, 1.922913, 1.933533, 1.937561, 1.933456, 1.905075, 1.860168, 
    1.812042, 1.760666, 1.724533, 1.708206, 1.704102, 1.710678, 1.710342, 
    1.709106, 1.705276, 1.70163, 1.694016, 1.680603, 1.670547, 1.671478, 
    1.69046, 1.692719, 1.682037, 1.719513, 1.727966, 1.754028, 1.770447, 
    1.800812, 1.80838, 1.775818, 1.806702, 1.762268, 1.837372, 1.593933, 
    1.557678, 1.582214, 1.632721, 1.685394, 1.7565, 1.800964, 1.821472, 
    1.84375, 1.853516, 1.857147, 1.890594, 1.943802, 1.966019, 1.950897, 
    1.94751, 1.999405, 2.071716, 2.131989, 2.165466, 2.153107, 2.11908, 
    2.082367, 2.087433, 2.090912, 2.055756, 2.036682, 2.016022, 2.01889, 
    2.032867, 2.054413, 2.043579, 2.01828, 2.00174, 1.976608, 1.946472, 
    1.915375, 1.901108, 1.905655, 1.914001, 1.901291,
  1.879089, 1.867188, 1.82193, 1.759888, 1.70665, 1.648438, 1.588867, 
    1.545105, 1.572983, 1.663742, 1.781448, 1.879745, 1.906052, 1.902145, 
    1.870255, 1.821945, 1.809174, 1.825134, 1.845642, 1.871231, 1.901169, 
    1.913681, 1.888031, 1.848236, 1.810745, 1.79863, 1.797134, 1.798309, 
    1.815308, 1.801239, 1.796234, 1.802414, 1.8125, 1.847198, 1.871552, 
    1.896225, 1.927795, 1.977615, 2.030014, 2.064697, 2.098633, 2.117493, 
    2.096527, 2.027832, 1.95639, 1.858185, 1.817627, 1.843994, 1.869324, 
    1.843201, 1.776611, 1.672455, 1.619843, 1.559937, 1.570709, 1.687988, 
    1.682098, 1.635315, 1.672241, 1.776672, 1.820251, 1.813904, 1.819763, 
    1.843658, 1.867096, 1.869919, 1.860779, 1.816589, 1.882202, 1.997955, 
    2.063339, 2.137817, 2.163544, 2.146484, 2.134827, 2.101013, 2.120941, 
    2.013275, 1.957153, 1.9198, 1.899353, 1.876282, 1.826538, 1.796143, 
    1.748505, 1.755798, 1.779297, 1.820862, 1.90213, 1.944122, 1.91626, 
    1.893799, 1.873428, 1.872009, 1.840103, 1.851563,
  2.022919, 2.072723, 2.105804, 2.066605, 2.003326, 1.907227, 1.819336, 
    1.765945, 1.714706, 1.731705, 1.757034, 1.775726, 1.77948, 1.817444, 
    1.882217, 1.893829, 1.881836, 1.877075, 1.919922, 1.943817, 1.958725, 
    1.926498, 1.865952, 1.808395, 1.714844, 1.657745, 1.707809, 1.818497, 
    1.941864, 1.998825, 2.017319, 2.012436, 1.978775, 1.976044, 1.981964, 
    2.004807, 1.996353, 1.987503, 2.022919, 2.063477, 2.086975, 2.074402, 
    2.054932, 1.979736, 1.921509, 1.919189, 1.186249, 1.327728, 1.309357, 
    1.236572, 1.170593, 1.097656, 0.9614258, 0.9257202, 0.9371338, 0.9135742, 
    0.8670959, 1.217438, 1.294403, 1.420959, 1.58252, 1.654297, 1.805695, 
    1.862213, 1.893677, 1.896393, 1.853821, 1.819794, 1.843353, 1.857147, 
    1.872894, 1.94101, 1.99353, 2.010468, 1.973511, 1.862091, 1.792175, 
    1.792572, 1.756683, 1.833984, 1.537689, 1.503784, 1.493652, 1.529083, 
    1.576416, 1.557281, 1.468353, 1.346008, 1.328796, 1.507996, 1.590759, 
    1.674988, 1.772888, 1.774948, 1.807693, 1.912308,
  1.887787, 1.945694, 2.066772, 2.10463, 2.12207, 2.041153, 2.002609, 
    1.924225, 1.856003, 1.85083, 1.822784, 1.835541, 1.837311, 1.855865, 
    1.833466, 1.858139, 1.874023, 1.866531, 1.85051, 1.849213, 1.893997, 
    1.913727, 1.861465, 1.855804, 1.861526, 1.868164, 1.913742, 2.0392, 
    2.069336, 2.061783, 2.044922, 2.064194, 2.095383, 2.129623, 2.129501, 
    2.086914, 2.077286, 2.045578, 2.022339, 2.021942, 1.992447, 1.972885, 
    1.972321, 1.991089, 1.952637, 1.930573, 1.220642, 1.223419, 1.132385, 
    1.044128, 0.9141846, 0.8389893, 0.811615, 0.8339844, 0.8468628, 
    0.8405457, 0.8505554, 0.8747864, 0.8536987, 0.8529968, 0.8690186, 
    0.8504333, 0.8981628, 0.9721069, 0.984314, 1.037994, 1.027252, 0.9372864, 
    0.7437439, 0.5198364, 1.071075, 0.8531799, 0.9985657, 1.061829, 1.083252, 
    0.9375, 1.525391, 1.523102, 1.598358, 1.664948, 1.354736, 1.353088, 
    1.391785, 1.473877, 1.551941, 1.557556, 1.620483, 1.573334, 1.491058, 
    1.381561, 1.402771, 1.737671, 1.686615, 1.756775, 1.788269, 1.824463,
  1.19574, 0.9529724, 1.866516, 1.933838, 1.942932, 1.922913, 1.891083, 
    1.87558, 1.870483, 1.837341, 1.962769, 2.00174, 1.917694, 1.917175, 
    1.911102, 1.882782, 1.813263, 1.670319, 1.549469, 1.579773, 1.597351, 
    1.641632, 1.684479, 1.710083, 1.755737, 1.776672, 1.767761, 1.798035, 
    1.840088, 1.743805, 1.613708, 1.476257, 1.537292, 1.638702, 1.581757, 
    1.518341, 1.516785, 1.485657, 1.496338, 1.533173, 1.601624, 1.753113, 
    1.70636, 1.455139, 0.8734131, 0.8919983, 0.936554, 0.8503723, 0.652771, 
    0.5447083, 0.4343567, 0.4076538, 0.4021301, 0.3693237, 0.3832092, 
    0.4152832, 0.4664307, 0.5297546, 0.5603943, 0.5895081, 0.6255798, 
    0.6704712, 0.6385193, 0.6383362, 0.6251831, 0.6166992, 0.5924377, 
    0.5461426, 0.5267334, 0.5506287, 0.6591492, 0.7986145, 0.8746643, 
    0.9473572, 0.9624023, 0.87677, 0.7316284, 0.5986938, 1.324799, 1.408173, 
    1.235779, 1.28833, 1.261383, 1.218201, 1.282288, 1.343811, 1.390991, 
    1.406311, 1.433502, 1.429993, 1.415802, 1.378876, 1.345551, 1.271912, 
    1.242249, 1.2677,
  0.9569702, 1.03418, 1.203308, 1.351227, 1.453705, 1.413086, 1.376221, 
    1.405914, 1.436188, 1.453613, 1.449799, 1.420441, 1.47641, 1.529449, 
    1.574677, 1.495972, 1.326355, 1.142242, 0.9647217, 0.8876953, 0.879364, 
    0.9115601, 1.032867, 1.172058, 1.149078, 1.061584, 0.924469, 0.7615662, 
    0.6633911, 0.5419006, 0.4844055, 0.4067688, 0.3822021, 1.35025, 1.485596, 
    1.552338, 0.9785461, 0.8111877, 0.6152039, 0.4996033, 0.4593506, 
    0.4042053, 0.3257141, 0.3225098, 0.351532, 0.3060913, 0.2131958, 
    0.1372681, 0.09014893, 0.1052551, 0.1490479, 0.1363831, 0.08233643, 
    0.03292847, -0.009155273, 0.02856445, 0.2018127, 0.3303223, 0.3803711, 
    0.4301147, 0.5059814, 0.5685425, 0.5773926, 0.6596069, 0.7564087, 
    0.8786926, 0.8922424, 0.9347534, 0.9830017, 1.036285, 1.104858, 1.156555, 
    1.22226, 1.198242, 1.149353, 1.075378, 0.9884338, 0.9649048, 1.099915, 
    1.257446, 0.9371033, 0.7403564, 0.6646423, 0.6730042, 0.7902832, 
    0.8812256, 0.8959656, 0.8874817, 0.9867249, 1.107513, 1.19223, 1.204346, 
    1.170105, 1.14093, 1.058502, 1.03183,
  0.7252502, 0.6498413, 0.6366577, 0.6838379, 0.708374, 0.685791, 0.7396851, 
    0.8741455, 1.006561, 1.084595, 1.08902, 1.127045, 1.217621, 1.237885, 
    1.212555, 1.144318, 1.132751, 1.143219, 1.027924, 0.8695679, 0.7600708, 
    0.7063599, 0.6976013, 0.727417, 0.7547302, 0.7680054, 0.6878052, 
    0.6063843, 0.556488, 0.5107727, 0.4273376, 0.4384766, 0.4814453, 
    0.5705566, 0.6653137, 0.846405, 0.9303589, 0.8892822, 0.842865, 0.821106, 
    0.8128357, 0.8466187, 0.9447937, 1.004364, 0.9651794, 0.7903137, 
    0.5024719, 0.2922363, 0.1158142, -0.1164551, -0.3583984, -0.5137329, 
    -0.6070557, -0.6642456, -0.5093079, -0.2617188, 0.004821777, 0.1333313, 
    0.2254944, 0.367981, 0.5584717, 0.6677551, 0.7496948, 0.8964844, 
    1.090363, 1.273102, 1.419006, 1.536774, 1.644196, 1.849609, 2.084839, 
    2.2565, 2.331329, 2.327728, 2.311829, 2.2612, 2.173706, 2.046234, 
    1.920898, 1.735474, 1.555786, 1.345184, 1.102203, 1.050476, 1.102875, 
    1.054535, 0.9751587, 0.9012756, 0.8244019, 0.7663879, 0.7705688, 
    0.8085022, 0.8678894, 0.9151001, 0.8785706, 0.8033752,
  1.095856, 0.9676514, 0.91745, 0.9365845, 1.00293, 1.050262, 1.100006, 
    1.142822, 1.151367, 1.167114, 1.233917, 1.366455, 1.443359, 1.47641, 
    1.513214, 1.572205, 1.637085, 1.640289, 1.576324, 1.53125, 1.521484, 
    1.431641, 1.359314, 1.345642, 1.367462, 1.366608, 1.307739, 1.264343, 
    1.20401, 1.12323, 0.9724426, 0.8125, 0.7424622, 0.6667175, 0.5335083, 
    0.4553833, 0.625, 0.9338074, 1.151062, 1.234711, 1.218567, 1.333984, 
    1.572601, 1.661469, 1.60144, 1.533508, 1.303833, 0.8744202, 0.3769531, 
    -0.09967041, -0.3970642, -0.4658813, -0.4697876, -0.5359802, -0.5901794, 
    -0.5175781, -0.4101563, -0.3997498, -0.3699646, 0.01031494, 0.4760437, 
    0.7495422, 0.966156, 1.261047, 1.554108, 1.696533, 1.818298, 1.995331, 
    2.100067, 2.176056, 2.282898, 2.375183, 2.407166, 2.365692, 2.240295, 
    1.999481, 1.613281, 1.503448, 1.556702, 1.694458, 1.812561, 1.811005, 
    1.618164, 1.288544, 1.13797, 1.153259, 1.224335, 1.267059, 1.231049, 
    1.194275, 1.27713, 1.379211, 1.395172, 1.303986, 1.230988, 1.192963,
  1.458618, 1.553314, 1.674866, 1.801758, 1.864471, 1.888824, 1.90332, 
    1.896179, 1.912781, 1.929169, 1.923553, 1.946106, 1.927795, 1.982086, 
    2.135803, 2.275848, 2.419922, 2.550964, 2.439209, 1.954315, 1.672729, 
    1.623047, 1.566925, 1.538361, 1.630676, 1.76178, 1.856659, 1.918182, 
    1.940765, 1.975647, 1.905273, 1.693024, 1.476166, 1.303986, 1.162933, 
    1.139862, 1.29129, 1.495728, 1.638214, 1.647858, 1.631714, 1.699615, 
    1.779755, 1.696716, 1.638397, 1.643768, 1.59317, 1.341278, 1.01535, 
    0.755127, 0.5991821, 0.5859985, 0.5033875, 0.3504028, 0.2325439, 
    0.1665955, 0.136261, 0.1413879, 0.1947327, 0.4028625, 0.6965332, 
    0.8743591, 1.027283, 1.259003, 1.466675, 1.489563, 1.538208, 1.692719, 
    1.785553, 1.824799, 1.881226, 1.931396, 1.938354, 1.885864, 1.688751, 
    1.275513, 1.227203, 1.472809, 1.646301, 1.736603, 1.708649, 1.644318, 
    1.598175, 1.42807, 1.328644, 1.425049, 1.633972, 1.754364, 1.70755, 
    1.656982, 1.65509, 1.679749, 1.671265, 1.607727, 1.529114, 1.460815,
  1.865509, 2.023956, 2.188416, 2.326965, 2.447083, 2.529541, 2.571594, 
    2.613892, 2.633606, 2.72995, 2.882813, 2.921997, 2.897186, 2.896698, 
    2.92337, 2.950439, 3.015472, 3.21756, 3.234375, 2.92981, 2.660095, 
    2.610291, 2.48822, 2.30423, 2.272858, 2.464783, 2.611725, 2.562225, 
    2.463013, 2.478577, 2.49173, 2.347534, 2.100525, 1.859589, 1.695038, 
    1.620636, 1.619537, 1.615356, 1.572083, 1.602936, 1.752136, 1.892365, 
    1.869965, 1.780548, 1.789612, 1.848267, 1.818451, 1.694824, 1.565216, 
    1.491699, 1.500488, 1.450684, 1.284607, 1.122101, 1.057709, 0.993988, 
    0.9331055, 0.9238586, 0.9451599, 1.029144, 1.175812, 1.285645, 1.354553, 
    1.44043, 1.533875, 1.53418, 1.540558, 1.577606, 1.598053, 1.643188, 
    1.670776, 1.636078, 1.56076, 1.467865, 1.298096, 1.217407, 1.395508, 
    1.69812, 1.949097, 1.999054, 1.804047, 1.667175, 1.601868, 1.533386, 
    1.494263, 1.672516, 1.928558, 2.135284, 2.221619, 2.227661, 2.165894, 
    2.028229, 1.921143, 1.912109, 1.889191, 1.827667,
  1.943878, 2.124329, 2.283997, 2.380005, 2.473511, 2.627289, 2.870789, 
    3.09024, 3.154755, 3.248657, 3.450836, 3.567383, 3.556, 3.468353, 
    3.317047, 3.144745, 3.08606, 3.146271, 3.166931, 3.172852, 3.303802, 
    3.371185, 3.229065, 2.933624, 2.799652, 2.737396, 2.596832, 2.416901, 
    2.299316, 2.253204, 2.240601, 2.151093, 1.967285, 1.841064, 1.769257, 
    1.734344, 1.73996, 1.612457, 1.437775, 1.535126, 1.919952, 2.091309, 
    2.099701, 2.054321, 2.163391, 2.189545, 2.331238, 2.258179, 2.119232, 
    2.111572, 2.236298, 2.240723, 2.056213, 1.857391, 1.744354, 1.652039, 
    1.588379, 1.590057, 1.598145, 1.575378, 1.576294, 1.582184, 1.550598, 
    1.519165, 1.524384, 1.546722, 1.579407, 1.585968, 1.530182, 1.455902, 
    1.414398, 1.417816, 1.417267, 1.340698, 1.279846, 1.283508, 1.599884, 
    2.013336, 2.545013, 1.967743, 1.717804, 1.529388, 1.602234, 1.687866, 
    1.748169, 1.860016, 1.93399, 1.965424, 2.0448, 2.075592, 2.001129, 
    1.913147, 1.832947, 1.767456, 1.785431, 1.844116,
  2.024963, 2.185577, 2.372955, 2.485077, 2.641846, 2.997681, 3.491577, 
    3.860107, 4.087402, 4.341949, 4.576538, 4.48584, 4.075623, 3.719757, 
    3.389801, 3.130615, 3.008057, 2.947357, 2.928101, 2.93869, 2.862854, 
    2.698395, 2.462494, 2.190063, 2.039612, 1.996582, 1.961487, 1.947021, 
    1.959686, 1.94754, 1.934845, 1.930084, 1.915405, 1.896912, 1.809998, 
    1.752106, 1.741119, 1.572571, 1.554657, 1.902588, 2.311554, 2.376068, 
    2.390076, 2.41568, 2.503326, 2.660919, 3.202972, 2.693787, 2.695099, 
    2.701324, 2.860962, 2.812531, 2.566101, 2.297607, 2.119629, 2.004211, 
    1.905914, 1.831543, 1.759613, 1.697418, 1.671112, 1.66333, 1.645233, 
    1.652771, 1.670013, 1.634796, 1.629578, 1.600159, 1.54184, 1.542542, 
    1.514465, 1.547485, 1.585968, 1.484863, 1.389679, 1.325043, 1.516235, 
    2.159332, 2.888184, 2.034668, 1.784576, 1.594299, 1.712463, 2.051208, 
    2.176208, 2.105255, 1.977295, 1.898163, 1.995667, 2.046082, 1.961609, 
    1.934143, 1.929657, 1.870026, 1.88974, 1.951263,
  2.044891, 2.168396, 2.215271, 2.300293, 2.550873, 2.969574, 3.270935, 
    3.821381, 4.050079, 3.788422, 3.400085, 3.047058, 2.662598, 2.40329, 
    2.249969, 2.182281, 2.144623, 2.051422, 1.966064, 1.83493, 1.705292, 
    1.657501, 1.617584, 1.509338, 1.388306, 1.420074, 1.516632, 1.538818, 
    1.641815, 1.818848, 2.017029, 2.027893, 1.892914, 1.736237, 1.659729, 
    1.706757, 1.838837, 1.908844, 2.198792, 3.808502, 2.601929, 2.672607, 
    2.954865, 2.874969, 2.714935, 2.763428, 2.838257, 2.998413, 2.690399, 
    2.533478, 2.399902, 2.3255, 2.257629, 2.181885, 2.035645, 1.973541, 
    1.916504, 1.833221, 1.780396, 1.764221, 1.78009, 1.785767, 1.765411, 
    1.771667, 1.788177, 1.771515, 1.806427, 1.79248, 1.746216, 1.804138, 
    1.753937, 1.715271, 1.689758, 1.587341, 1.497284, 1.299896, 1.458557, 
    3.157837, 3.386566, 2.622192, 1.697083, 1.695282, 2.061554, 2.394287, 
    2.339203, 2.122681, 2.054749, 2.004852, 2.010345, 1.988373, 1.934204, 
    1.948669, 1.904083, 1.861938, 1.867493, 1.90387,
  1.890594, 1.829681, 1.863068, 2.065979, 2.327972, 2.436249, 2.558105, 
    2.786621, 2.949341, 2.602936, 1.97226, 1.787201, 1.757446, 1.836365, 
    1.803741, 1.739746, 1.671448, 1.538116, 1.480072, 1.39563, 1.367737, 
    1.359863, 1.283295, 1.319122, 1.349579, 1.477203, 1.662384, 1.78598, 
    2.06488, 2.221832, 1.989838, 2.04599, 1.945953, 1.819244, 1.82196, 
    1.868866, 1.984283, 3.132599, 3.773376, 3.961792, 2.911194, 2.800507, 
    3.354919, 3.149048, 2.926483, 2.947388, 2.793182, 2.529053, 2.246338, 
    1.921204, 1.788391, 1.774323, 1.799622, 1.813904, 1.814026, 1.84259, 
    1.832062, 1.804016, 1.809662, 1.842865, 1.908508, 1.939789, 1.948975, 
    1.960785, 1.98761, 1.925232, 1.862793, 1.831299, 1.805237, 1.741791, 
    1.695221, 1.675568, 1.546326, 1.345215, 1.27713, 1.099243, 1.374817, 
    4.23468, 3.647034, 1.153046, 0.8424988, 1.725647, 2.008698, 2.375671, 
    2.258484, 2.014435, 2.013489, 2.043182, 1.996521, 1.825104, 1.760254, 
    1.801514, 1.741577, 1.777588, 1.825287, 1.840576,
  1.70636, 1.641571, 1.694672, 1.808289, 2.047791, 3.885681, 4.429413, 
    3.557373, 2.728119, 2.248199, 2.17157, 2.261139, 2.247314, 2.19754, 
    2.091614, 2.04538, 2.067749, 1.988464, 1.939514, 1.911285, 1.916443, 
    1.962006, 2.022034, 2.087646, 2.129852, 2.19632, 2.336548, 2.36142, 
    2.259064, 1.865814, 2.164642, 4.293091, 3.868164, 3.393738, 3.536652, 
    3.48587, 3.456116, 3.589722, 3.787903, 3.56665, 2.800964, 2.08255, 
    1.816345, 1.903442, 2.201294, 2.376556, 2.143036, 1.710175, 1.655792, 
    1.712616, 1.752594, 1.847382, 1.891815, 1.908356, 1.878357, 1.872803, 
    1.870422, 1.868378, 1.862671, 1.907532, 1.929993, 1.918274, 1.927307, 
    1.845673, 1.830597, 1.748566, 1.632416, 1.524353, 1.456757, 1.386627, 
    1.286804, 1.268341, 1.174316, 1.093384, 1.005432, 0.9007874, 1.199188, 
    3.069641, 3.364838, 1.642334, 1.791718, 2.5112, 2.343018, 2.221161, 
    2.135223, 1.997253, 2.005737, 1.920105, 1.922455, 1.893219, 1.856964, 
    1.841583, 1.754364, 1.73468, 1.727509, 1.740326,
  1.501038, 1.479614, 1.654907, 1.739044, 2.442871, 4.052521, 3.942535, 
    3.256958, 2.75589, 2.227478, 2.215179, 2.370728, 2.301086, 2.282623, 
    2.4487, 2.545624, 2.596558, 2.52774, 2.451233, 2.4599, 2.406586, 
    2.368164, 2.307434, 2.261261, 2.208923, 2.124542, 2.062286, 1.949921, 
    1.940308, 1.900391, 2.60611, 5.054413, 4.597321, 4.050201, 3.988861, 
    3.824402, 4.035156, 3.826477, 3.602203, 3.392273, 2.435822, 1.593994, 
    1.277283, 1.439911, 1.768494, 1.963623, 2.006897, 2.009888, 2.07962, 
    2.168671, 2.172791, 2.084503, 2.023163, 1.942535, 1.854767, 1.752136, 
    1.696625, 1.695984, 1.6763, 1.703125, 1.698181, 1.659637, 1.59201, 
    1.427216, 1.357361, 1.317719, 1.2995, 1.194794, 1.138977, 1.113403, 
    1.026306, 1.049072, 1.000397, 0.9554443, 0.7951965, 1.019379, 1.524689, 
    2.840637, 3.977234, 2.633545, 2.185425, 2.867126, 3.025848, 2.913147, 
    2.311188, 2.098694, 2.124786, 2.035309, 1.974152, 1.916748, 1.906189, 
    1.837616, 1.775909, 1.742523, 1.616669, 1.591614,
  1.614471, 1.728912, 1.938416, 2.265381, 3.509491, 3.459442, 2.809204, 
    3.247406, 3.080841, 2.61615, 2.3367, 2.477081, 2.920563, 2.326416, 
    2.312561, 2.47702, 2.328583, 2.265015, 2.166534, 2.093811, 2.040955, 
    2.001556, 1.978455, 1.95697, 1.960938, 1.926117, 1.882996, 1.90155, 
    2.045776, 2.097504, 2.471436, 4.386841, 4.585114, 4.430054, 4.067566, 
    3.548248, 3.934967, 3.735962, 3.431854, 3.184631, 2.296173, 1.661133, 
    1.794342, 2.05011, 2.111206, 2.147522, 2.172058, 2.223175, 2.186859, 
    2.150787, 2.09848, 1.989319, 1.917206, 1.816345, 1.725189, 1.659821, 
    1.614075, 1.648499, 1.630127, 1.569855, 1.510986, 1.392365, 1.325531, 
    1.260437, 1.262115, 1.234375, 1.21756, 1.117706, 1.093231, 1.013519, 
    1.046173, 1.057617, 0.8429565, 0.9199524, 0.9476929, 1.515137, 2.328278, 
    3.733978, 5.32132, 3.254211, 2.349792, 3.041534, 3.187897, 3.197876, 
    3.1362, 2.344727, 2.082825, 2.098419, 2.045197, 1.895721, 1.796356, 
    1.683716, 1.605408, 1.572662, 1.555267, 1.575043,
  1.940247, 2.085083, 2.19928, 2.325989, 3.53064, 3.365021, 3.172272, 
    3.624817, 3.444153, 3.02359, 2.458984, 2.408478, 2.839508, 2.843689, 
    2.186707, 2.196411, 2.088135, 2.111572, 2.105316, 2.057678, 2.057434, 
    2.0401, 2.041016, 1.99884, 1.987122, 1.989197, 2.064117, 2.145172, 
    2.280914, 2.315948, 2.303497, 2.775055, 4.170441, 4.753906, 4.269531, 
    3.605011, 3.429749, 3.060944, 3.018036, 2.781647, 1.891083, 1.938141, 
    2.077789, 2.163666, 2.209503, 2.266327, 2.292053, 2.31192, 2.274567, 
    2.274292, 2.217896, 2.133392, 2.039246, 1.980255, 1.9487, 1.889648, 
    1.842255, 1.819794, 1.806305, 1.745575, 1.704224, 1.647278, 1.675781, 
    1.61908, 1.53833, 1.471283, 1.415619, 1.356445, 1.34494, 1.301575, 
    1.260101, 1.30835, 1.281128, 1.542389, 1.486908, 1.693451, 2.504242, 
    4.379944, 5.641693, 3.634613, 2.712036, 3.064117, 2.945831, 3.242981, 
    4.045715, 4.471497, 2.08432, 2.049744, 1.968445, 1.859283, 1.776764, 
    1.714203, 1.705139, 1.70755, 1.769226, 1.872406,
  2.307404, 2.416718, 2.588684, 2.583649, 3.05072, 2.907471, 2.823029, 
    3.201508, 3.699097, 3.943604, 3.838013, 2.393097, 2.685211, 3.152863, 
    2.261963, 2.210815, 2.191528, 2.212158, 2.226685, 2.224548, 2.246033, 
    2.222992, 2.232758, 2.240997, 2.24585, 2.275726, 2.343811, 2.428894, 
    2.4664, 2.445831, 2.327545, 2.35321, 2.573761, 3.725769, 3.819611, 
    3.654297, 3.486847, 2.349365, 2.74942, 2.00351, 1.962433, 2.174927, 
    2.219147, 2.26886, 2.288849, 2.341553, 2.399353, 2.41037, 2.355865, 
    2.309357, 2.227997, 2.184509, 2.193268, 2.210663, 2.205139, 2.197205, 
    2.153595, 2.104492, 2.120514, 2.132416, 2.112305, 2.106262, 2.097321, 
    2.011017, 1.93515, 1.911652, 1.834564, 1.831909, 1.813812, 1.850922, 
    1.84967, 1.883728, 1.875183, 1.904755, 1.82724, 2.349609, 4.351501, 
    5.680756, 4.491028, 3.313416, 2.961243, 3.269714, 3.254547, 3.17688, 
    4.557343, 4.820374, 1.985504, 2.069794, 1.999023, 1.949738, 2.018982, 
    2.005646, 2.113556, 2.165375, 2.243561, 2.301392,
  2.555267, 2.612305, 2.777344, 2.619141, 2.919586, 2.911713, 2.708527, 
    2.885742, 3.518433, 4.028198, 4.291656, 2.391541, 2.285156, 2.345825, 
    2.334381, 2.415314, 2.331757, 2.31192, 2.303436, 2.335693, 2.347961, 
    2.352142, 2.365753, 2.3573, 2.34317, 2.38678, 2.443237, 2.517517, 
    2.53241, 2.532104, 2.521088, 2.524292, 2.461914, 2.433899, 2.359161, 
    3.019135, 3.208801, 2.36731, 2.133331, 2.085327, 2.08255, 2.320251, 
    2.286713, 2.303619, 2.342346, 2.387054, 2.423676, 2.343353, 2.243622, 
    2.199982, 2.224091, 2.238342, 2.253754, 2.305267, 2.334503, 2.325867, 
    2.353271, 2.378723, 2.420837, 2.431122, 2.41452, 2.393036, 2.313538, 
    2.276947, 2.217651, 2.205658, 2.156128, 2.210602, 2.209778, 2.22937, 
    2.25177, 2.270691, 2.387817, 2.404449, 2.597656, 3.984711, 3.899841, 
    4.061493, 3.496063, 3.11795, 3.204498, 3.44043, 3.577148, 3.286072, 
    4.009766, 4.224152, 2.026642, 2.159912, 2.222015, 2.185272, 2.254761, 
    2.303711, 2.360016, 2.436981, 2.473694, 2.528961,
  2.703461, 2.702789, 2.692108, 2.494476, 3.093567, 3.0867, 2.796417, 
    2.606598, 2.921021, 3.636108, 3.544708, 2.322357, 2.4487, 2.48938, 
    2.464203, 2.56192, 2.461304, 2.388336, 2.319916, 2.354279, 2.374207, 
    2.399536, 2.399811, 2.456238, 2.480225, 2.472656, 2.472778, 2.451447, 
    2.436646, 2.498718, 2.451874, 2.497467, 2.540802, 2.474884, 2.470703, 
    2.360657, 2.338348, 2.371277, 2.253113, 2.125824, 2.164886, 2.33429, 
    2.226044, 2.176117, 2.155609, 2.151611, 2.193115, 2.181854, 2.137939, 
    2.144012, 2.239014, 2.276154, 2.29837, 2.363403, 2.395081, 2.404297, 
    2.42865, 2.489594, 2.493347, 2.52182, 2.518311, 2.5289, 2.503052, 
    2.488647, 2.458679, 2.477997, 2.491669, 2.473328, 2.522766, 2.559174, 
    2.626434, 2.652466, 2.757355, 2.705017, 2.652924, 3.11438, 3.380493, 
    3.610138, 3.744446, 3.454437, 3.25827, 3.333069, 3.527039, 3.549622, 
    3.200439, 3.656647, 3.420563, 2.340881, 2.384247, 2.385925, 2.370239, 
    2.450317, 2.467133, 2.579041, 2.627197, 2.66333,
  2.785095, 2.770386, 2.688019, 2.534241, 3.111328, 3.100708, 3.030914, 
    2.972351, 2.905243, 3.339172, 3.242249, 2.3638, 2.414337, 2.475769, 
    2.458588, 2.520691, 2.494019, 2.430359, 2.412231, 2.387177, 2.360992, 
    2.40567, 2.436371, 2.526764, 2.533997, 2.487244, 2.524078, 2.470184, 
    2.135223, 2.492706, 2.463165, 2.409912, 2.410492, 2.361206, 2.421265, 
    2.392761, 2.324036, 3.058136, 2.72171, 2.353455, 2.140747, 2.268768, 
    2.202423, 2.138, 2.035309, 2.101105, 2.245575, 2.355286, 2.496765, 
    2.582031, 2.630554, 2.684906, 2.717377, 2.725342, 2.730621, 2.746613, 
    2.755737, 2.775208, 2.73111, 2.743927, 2.743225, 2.767853, 2.782623, 
    2.784821, 2.788544, 2.754181, 2.766205, 2.74823, 2.797668, 2.779114, 
    2.821411, 2.856049, 2.799225, 2.699554, 2.625305, 3.504364, 4.026245, 
    3.658722, 3.649109, 3.254974, 3.570953, 3.611633, 3.722778, 4.212433, 
    3.303558, 2.930847, 3.243042, 2.430969, 2.493225, 2.455139, 2.459717, 
    2.554474, 2.580353, 2.67746, 2.699493, 2.740875,
  2.600128, 2.577362, 2.537872, 2.798187, 2.933197, 2.973633, 3.010071, 
    2.850037, 2.734558, 2.709808, 2.917084, 3.499603, 2.545135, 2.443878, 
    2.470184, 2.49408, 2.493378, 2.412201, 2.44812, 2.481628, 2.455353, 
    2.47879, 2.523224, 2.557617, 2.558594, 2.493744, 2.422333, 2.696106, 
    2.471436, 2.397308, 2.436371, 2.189117, 2.075195, 2.199219, 2.229309, 
    2.683258, 2.612885, 2.822723, 2.687408, 2.18457, 2.253632, 2.26947, 
    2.299408, 2.335297, 2.327423, 2.498108, 2.768829, 3.053925, 3.206116, 
    3.222137, 3.251099, 3.249481, 3.241272, 3.282104, 3.302155, 3.306976, 
    3.303192, 3.294983, 3.296967, 3.28775, 3.278259, 3.214264, 3.155212, 
    3.059784, 3.022614, 2.938538, 2.90802, 2.84668, 2.808258, 2.799408, 
    2.787781, 2.698517, 2.538727, 2.383514, 2.386078, 3.290039, 3.436188, 
    3.382965, 3.358215, 3.639069, 3.975739, 5.112762, 4.446442, 4.201843, 
    3.529816, 2.496155, 2.501373, 2.535095, 2.600586, 2.593231, 2.645569, 
    2.600922, 2.637482, 2.684448, 2.679352, 2.631836,
  2.471954, 2.699371, 2.5979, 3.026581, 2.997772, 2.930786, 2.698883, 
    2.517456, 2.537231, 2.910278, 2.49765, 3.425323, 3.464386, 2.575775, 
    2.561249, 2.475067, 2.489349, 2.479309, 2.446564, 2.447327, 2.436768, 
    2.335236, 2.384247, 2.41687, 2.465118, 2.367004, 2.245544, 2.806488, 
    2.204376, 2.315552, 2.319, 2.310242, 2.369415, 2.156952, 2.130249, 
    2.117249, 2.040161, 2.109375, 2.208405, 2.232819, 2.176086, 2.182037, 
    2.220398, 2.249268, 2.294128, 2.439392, 2.723175, 3.016663, 3.140167, 
    3.153656, 3.18103, 3.219727, 3.197266, 3.171509, 3.141266, 3.14325, 
    3.214691, 3.218323, 3.252014, 3.19342, 3.186005, 3.080597, 3.023621, 
    2.941071, 2.884308, 2.816559, 2.734497, 2.723724, 2.734436, 2.723694, 
    2.67572, 2.577148, 2.390503, 2.129028, 2.0065, 2.879425, 3.636932, 
    4.009705, 3.294678, 3.864899, 4.736145, 4.457092, 3.790833, 2.416809, 
    2.358521, 2.337952, 2.358734, 2.426575, 2.454773, 2.516327, 2.548431, 
    2.542511, 2.613953, 2.532288, 2.532043, 2.429901,
  3.388275, 2.879639, 3.267761, 3.535858, 3.107544, 3.030609, 2.897461, 
    2.689575, 2.921082, 3.167389, 3.057648, 2.708862, 2.856842, 2.527405, 
    2.496033, 2.464844, 2.492126, 2.496857, 2.447266, 2.397797, 2.384552, 
    2.343933, 2.321411, 2.272736, 2.305786, 2.325195, 2.742981, 3.161011, 
    2.240234, 2.229431, 2.19342, 2.888489, 2.27533, 2.296234, 2.215027, 
    2.143188, 2.165375, 2.208405, 2.212708, 2.164063, 2.144775, 2.162567, 
    2.153717, 2.131775, 2.120453, 2.202606, 2.340942, 2.412903, 2.526154, 
    2.63208, 2.683899, 2.759186, 2.782043, 2.800262, 2.816711, 2.756378, 
    2.722473, 2.66745, 2.596069, 2.522278, 2.472321, 2.425201, 2.4375, 
    2.453979, 2.487762, 2.523712, 2.54303, 2.610748, 2.728333, 2.824951, 
    2.913483, 2.759888, 2.462616, 2.286652, 2.357758, 3.131134, 4.300293, 
    4.863983, 4.330994, 5.373505, 4.341675, 3.940765, 2.580292, 2.481232, 
    2.443604, 2.419098, 2.427338, 2.443268, 2.459961, 2.41217, 2.447266, 
    2.419678, 2.425476, 2.476196, 3.179749, 3.285492,
  3.309875, 3.242584, 3.359894, 3.462433, 3.47168, 3.592499, 3.368744, 
    3.573364, 3.50885, 3.02121, 3.460358, 3.209198, 3.326752, 3.020264, 
    2.570526, 2.556702, 2.631439, 2.57428, 2.583252, 2.546997, 2.608276, 
    2.748169, 2.452087, 2.313721, 2.269989, 2.227081, 2.309357, 3.736725, 
    2.516663, 2.374725, 2.314758, 2.223694, 2.258545, 2.827789, 2.305939, 
    2.24585, 2.275726, 2.218597, 2.258087, 2.218689, 2.208923, 2.198975, 
    2.141541, 2.118927, 2.123901, 2.174133, 2.227325, 2.235992, 2.286652, 
    2.307892, 2.339325, 2.378265, 2.429535, 2.48111, 2.515259, 2.529816, 
    2.516998, 2.502716, 2.458527, 2.445892, 2.39798, 2.414795, 2.462616, 
    2.532928, 2.61731, 2.675507, 2.684753, 2.679504, 2.771667, 2.857117, 
    2.847992, 2.787048, 2.868378, 2.752533, 3.257874, 3.383942, 3.862183, 
    4.830811, 4.414764, 4.237457, 2.274414, 2.242706, 2.237823, 2.384247, 
    2.358276, 2.341919, 2.354309, 2.390533, 2.447632, 2.418732, 2.451324, 
    2.353394, 2.507751, 3.289673, 3.368469, 3.180298,
  3.748718, 3.185486, 2.697906, 2.656555, 2.990295, 3.270172, 3.351135, 
    3.663055, 3.827362, 3.977539, 4.113403, 4.491974, 4.071777, 3.531525, 
    2.682617, 2.658081, 2.71048, 2.670685, 2.667572, 2.647003, 3.190002, 
    3.318542, 2.562073, 2.437836, 2.334167, 2.234192, 2.2435, 3.850281, 
    3.572754, 2.861023, 2.324036, 2.322205, 2.260925, 2.733582, 2.246765, 
    2.203827, 2.186737, 2.193298, 2.247528, 2.259644, 2.239532, 2.220459, 
    2.205475, 2.221954, 2.270691, 2.281006, 2.291718, 2.300049, 2.377075, 
    2.422852, 2.469788, 2.483734, 2.543427, 2.621216, 2.631897, 2.672852, 
    2.633667, 2.618164, 2.556702, 2.526611, 2.522858, 2.528717, 2.539398, 
    2.594788, 2.659973, 2.697205, 2.723267, 2.74231, 2.679047, 2.66452, 
    2.721375, 2.884766, 3.94342, 3.769104, 2.49585, 2.428253, 2.305267, 
    2.274017, 2.260162, 2.282288, 2.310547, 2.372253, 2.295441, 2.281494, 
    2.26004, 2.309875, 2.323639, 2.412872, 2.469788, 2.507141, 2.533356, 
    2.700012, 3.4664, 3.893494, 3.782379, 3.345612,
  3.25647, 3.003082, 2.645325, 2.598938, 2.676331, 2.491486, 2.563812, 
    2.569885, 2.492401, 2.938293, 4.233093, 4.635651, 3.673065, 3.609222, 
    3.27179, 2.677521, 2.724823, 2.759308, 2.718079, 2.691406, 3.46286, 
    3.552246, 2.757568, 2.664703, 2.418945, 2.335541, 3.736603, 3.790649, 
    3.313324, 2.194, 2.22937, 2.268768, 2.136658, 2.074158, 2.219452, 
    2.191071, 2.119202, 2.207245, 2.24585, 2.274689, 2.286133, 2.247253, 
    2.264252, 2.277344, 2.303955, 2.27832, 2.286652, 2.32428, 2.363739, 
    2.384888, 2.40097, 2.43985, 2.459442, 2.483459, 2.470123, 2.436401, 
    2.403717, 2.398254, 2.366028, 2.311646, 2.264984, 2.242523, 2.273773, 
    2.315582, 2.381775, 2.513733, 2.567963, 2.486328, 2.335022, 2.702942, 
    3.212006, 3.117096, 2.733856, 2.309906, 2.388672, 2.345306, 2.350037, 
    2.370819, 2.359375, 2.363953, 2.306427, 2.259888, 2.212769, 2.181305, 
    2.156769, 2.164856, 2.174927, 2.301117, 2.366455, 2.460541, 2.45462, 
    2.731964, 3.645752, 3.545563, 3.633118, 3.317352,
  3.088989, 2.986755, 3.019714, 2.858887, 2.680939, 2.689362, 2.752563, 
    2.82132, 2.621582, 2.439972, 2.503204, 3.875641, 3.772949, 3.865082, 
    3.970917, 3.723297, 2.697662, 2.742065, 2.733124, 2.491028, 3.254547, 
    3.465393, 3.459015, 3.485626, 2.480072, 3.019836, 3.564148, 3.244812, 
    3.264282, 2.853729, 2.239655, 2.246094, 2.135345, 2.118286, 2.173553, 
    2.183594, 2.114258, 2.118286, 2.161652, 2.188538, 2.206818, 2.192383, 
    2.221985, 2.233704, 2.233917, 2.230072, 2.241516, 2.229034, 2.249207, 
    2.279572, 2.323639, 2.388092, 2.408722, 2.446014, 2.446289, 2.439972, 
    2.446014, 2.393768, 2.338593, 2.31308, 2.227234, 2.104309, 2.017334, 
    2.002411, 2.062836, 2.204865, 2.351837, 2.42746, 2.381287, 2.286011, 
    2.037781, 1.603699, 1.624146, 2.137512, 2.432404, 2.477875, 2.502686, 
    2.532013, 2.494476, 2.414703, 2.350372, 2.308136, 2.246399, 2.091919, 
    1.974762, 1.962006, 1.964508, 2.0625, 2.139008, 2.255219, 2.26712, 
    2.645233, 3.87738, 3.878296, 3.713959, 3.574829,
  4.066956, 3.703033, 3.201691, 3.113739, 2.932861, 2.517548, 2.466888, 
    2.825684, 2.975555, 2.867157, 2.448242, 3.630096, 3.369965, 3.40271, 
    3.836426, 3.907379, 2.786835, 2.942169, 4.06424, 3.403931, 2.877838, 
    2.833954, 2.600098, 3.009399, 3.00882, 2.561859, 2.746704, 2.782318, 
    2.882507, 2.969879, 2.748169, 2.672943, 2.162109, 2.139313, 2.127197, 
    2.167786, 2.187897, 2.133453, 2.158783, 2.100403, 2.083191, 2.076752, 
    2.084259, 2.103912, 2.101044, 2.103119, 2.087494, 2.093536, 2.123749, 
    2.164856, 2.186707, 2.183319, 2.178467, 2.18457, 2.226318, 2.247955, 
    2.251434, 2.239563, 2.261536, 2.275787, 2.240448, 2.130005, 2.017395, 
    1.921631, 1.916595, 2.002075, 2.358521, 2.80069, 2.592041, 2.322205, 
    2.270416, 2.048492, 1.951508, 2.063934, 2.227661, 2.31955, 2.37207, 
    2.483734, 2.621735, 2.57663, 2.528381, 2.439331, 2.365112, 2.292603, 
    2.201569, 2.123627, 2.066925, 2.067932, 2.04837, 2.038605, 2.032501, 
    2.312164, 3.636169, 4.127228, 4.032837, 4.145721,
  3.995209, 4.02829, 3.693237, 3.445374, 3.202087, 2.699646, 2.93811, 
    3.033142, 3.049072, 2.879669, 3.054047, 3.011292, 2.945099, 3.162781, 
    3.826874, 3.989655, 3.584747, 3.806396, 4.2948, 3.517822, 2.999908, 
    3.318726, 3.152618, 2.912994, 2.477386, 3.12619, 2.766846, 2.480103, 
    2.950012, 2.632477, 2.315826, 2.215637, 2.403778, 2.262177, 2.180359, 
    2.189758, 2.291351, 2.313599, 2.321747, 2.202087, 2.144958, 2.155151, 
    2.1698, 2.156769, 2.112579, 2.091003, 2.027405, 1.986237, 1.962891, 
    1.928101, 2.001831, 2.095398, 2.151428, 2.156586, 2.177795, 2.237366, 
    2.257355, 2.234375, 2.2117, 2.223877, 2.21701, 2.159363, 2.07486, 
    1.934906, 1.925812, 2.069702, 3.090973, 3.022003, 2.776825, 2.842194, 
    2.512268, 2.306244, 2.273712, 2.324432, 2.069885, 2.140869, 2.272278, 
    2.390411, 2.579224, 2.600861, 2.556976, 2.466614, 2.382996, 2.302216, 
    2.18985, 2.112244, 2.103973, 2.124664, 2.135681, 2.059387, 1.989471, 
    2.032501, 2.42099, 3.819183, 4.113922, 3.810272,
  3.364044, 3.50293, 3.389404, 3.444214, 3.30304, 2.43042, 2.615723, 
    2.650085, 2.269623, 2.543549, 2.381378, 2.712036, 2.752869, 2.944519, 
    2.828918, 3.005127, 3.008911, 3.295654, 4.218811, 3.949615, 3.915192, 
    6.419891, 4.844772, 3.893661, 3.541626, 3.850189, 2.849792, 1.738342, 
    3.019653, 3.618561, 2.475281, 2.253326, 2.437103, 2.05368, 2.057129, 
    2.354187, 2.520081, 2.560181, 2.515778, 2.39978, 2.308868, 2.256561, 
    2.244354, 2.230591, 2.193787, 2.163177, 2.112152, 2.070435, 2.055634, 
    2.041321, 2.0495, 2.012909, 2.056091, 2.163727, 2.223663, 2.279175, 
    2.263123, 2.231812, 2.205231, 2.255493, 2.164612, 2.039307, 1.957977, 
    1.897369, 2.035919, 2.869415, 2.844147, 2.351898, 2.345764, 2.764465, 
    2.464844, 1.962494, 1.594513, 1.698181, 1.95401, 2.066284, 2.149628, 
    2.182281, 2.242706, 2.255066, 2.303131, 2.366669, 2.350769, 2.243225, 
    2.131317, 2.063538, 2.005005, 2.046204, 2.134125, 2.132111, 2.142365, 
    2.079254, 2.115662, 2.476868, 3.806244, 3.254608,
  3.159698, 2.602875, 2.769867, 2.753479, 2.598083, 2.365784, 2.038391, 
    1.945801, 2.153076, 2.342438, 2.128326, 2.432739, 2.303772, 2.514313, 
    2.715668, 2.910858, 2.894928, 3.020844, 4.794891, 4.894318, 5.104141, 
    5.169235, 4.535599, 4.150879, 3.775299, 4.253906, 4.5065, 2.073242, 
    3.868683, 3.907532, 2.312561, 2.314362, 2.256714, 2.391022, 3.081909, 
    2.563965, 3.384979, 3.561005, 2.683228, 2.574768, 2.449951, 2.357452, 
    2.30954, 2.288177, 2.243805, 2.184662, 2.16156, 2.179504, 2.157166, 
    2.12381, 2.138428, 2.141693, 2.204132, 2.286682, 2.34201, 2.424011, 
    2.425659, 2.361938, 2.32251, 2.266174, 2.153564, 2.058441, 1.994263, 
    1.934265, 2.359497, 2.249207, 1.958069, 1.747253, 2.08316, 2.429749, 
    2.284454, 2.119598, 2.137634, 2.115479, 2.210205, 2.393158, 2.424103, 
    2.368713, 2.277588, 2.242249, 2.125275, 1.898315, 1.905151, 2.026184, 
    1.930389, 1.796448, 1.722626, 1.823975, 2.133636, 2.357788, 2.363373, 
    2.262665, 2.193665, 2.402893, 2.64859, 3.164825,
  2.975586, 2.74234, 2.677032, 2.600281, 2.525574, 2.413849, 2.445526, 
    1.831177, 1.763672, 1.656097, 1.917053, 3.030365, 2.772369, 2.370636, 
    2.163391, 2.578125, 2.433594, 2.385101, 2.983643, 5.080383, 5.208054, 
    5.559418, 5.342743, 5.258575, 4.458588, 4.92099, 5.217087, 4.995941, 
    4.026031, 3.524048, 3.183319, 2.740021, 2.498749, 3.349274, 3.589752, 
    2.86676, 2.750549, 3.079956, 2.656464, 2.662842, 2.623138, 2.591187, 
    2.536682, 2.499512, 2.510101, 2.486115, 2.389465, 2.341125, 2.318024, 
    2.276001, 2.23291, 2.20047, 2.246887, 2.309326, 2.352966, 2.401733, 
    2.425476, 2.435059, 2.427185, 2.36731, 2.252777, 2.047028, 1.891632, 
    2.067841, 2.468933, 2.581665, 2.753235, 2.746613, 2.32132, 1.422424, 
    1.710327, 1.906311, 2.159119, 2.134247, 2.166595, 2.538361, 3.097748, 
    3.168213, 2.991577, 2.775757, 2.506073, 2.023804, 1.793396, 1.935242, 
    1.889801, 1.56781, 1.187286, 1.087585, 1.49704, 2.003937, 2.287384, 
    2.292267, 2.208435, 2.319305, 2.699341, 2.950653,
  2.700653, 2.543243, 2.604919, 2.868347, 2.581604, 2.942322, 3.042603, 
    2.464783, 1.820435, 1.676361, 2.131836, 2.898926, 2.541779, 2.048553, 
    2.157562, 2.796478, 3.209625, 2.753326, 2.808075, 4.158386, 4.653687, 
    5.269379, 5.562866, 5.605835, 5.295349, 5.147461, 4.8311, 5.024918, 
    5.671616, 5.489838, 4.839691, 4.542572, 4.301086, 3.751678, 4.405777, 
    4.685455, 3.266449, 2.954224, 3.220367, 3.49585, 3.291138, 2.92572, 
    2.688232, 2.504822, 2.431702, 2.41217, 2.31366, 2.222534, 2.159973, 
    2.125702, 2.124023, 2.153229, 2.254089, 2.398041, 2.440857, 2.395935, 
    2.355896, 2.390198, 2.384399, 2.304016, 2.228821, 2.128357, 2.006805, 
    2.258148, 2.808075, 3.229279, 2.917755, 2.31131, 1.978363, 1.553436, 
    1.499329, 1.557129, 2.069885, 2.221893, 2.828278, 3, 3.18689, 3.171875, 
    3.317841, 3.232361, 2.799255, 2.384857, 2.30484, 1.902313, 1.600342, 
    1.439484, 1.14743, 0.7233276, 0.8927917, 1.415466, 1.873718, 2.147858, 
    2.113129, 2.046753, 2.193817, 2.397919,
  2.263763, 2.419525, 3.114838, 3.342712, 2.81662, 2.501678, 2.556091, 
    1.897522, 1.746948, 1.578918, 1.454803, 1.488861, 1.45578, 1.405853, 
    1.942261, 2.925049, 3.923279, 4.32843, 4.360809, 4.382599, 4.541901, 
    4.761627, 5.090225, 4.795105, 4.448364, 3.856842, 3.471878, 3.356903, 
    3.884247, 4.012405, 3.934799, 4.832397, 5.177719, 5.191238, 4.961624, 
    5.580856, 5.595291, 3.24939, 3.20343, 2.81134, 2.518372, 2.423584, 
    2.386993, 2.318878, 2.217834, 2.163849, 2.153381, 2.176422, 2.210999, 
    2.224365, 2.242645, 2.255463, 2.291382, 2.335083, 2.398163, 2.46582, 
    2.489258, 2.464783, 2.431458, 2.369354, 2.27829, 2.146912, 2.049652, 
    2.408844, 3.410919, 3.485901, 3.164825, 2.533783, 2.20517, 2.017761, 
    2.103119, 2.130188, 2.606445, 2.905731, 3.011963, 3.485474, 3.751221, 
    3.996216, 3.915222, 3.52771, 3.026581, 2.535614, 1.92337, 1.602997, 
    1.460083, 1.349365, 1.028046, 0.4842224, 0.3317261, 0.7064819, 1.154907, 
    1.594238, 1.83194, 1.933441, 2.027924, 2.150146,
  2.02124, 2.158844, 2.732422, 2.952484, 2.754211, 2.684357, 2.353241, 
    1.865875, 1.968323, 2.37204, 2.419403, 2.436493, 2.292816, 2.032196, 
    2.450073, 2.933319, 3.147064, 3.393341, 3.685272, 3.83017, 4.221222, 
    4.738922, 4.521667, 3.526337, 3.954498, 3.208923, 3.008469, 2.729691, 
    3.244461, 3.392899, 3.909302, 4.486588, 4.751038, 4.887512, 4.932159, 
    5.159637, 5.176697, 4.705978, 2.816498, 2.432678, 2.415558, 2.422607, 
    2.446625, 2.244598, 2.158783, 2.176575, 2.20813, 2.239594, 2.300018, 
    2.330475, 2.327087, 2.371277, 2.499084, 2.631378, 2.721893, 2.766449, 
    2.739441, 2.626373, 2.539063, 2.455994, 2.279755, 2.131653, 2.5867, 
    3.431671, 3.503235, 3.320251, 3.220612, 3.091919, 3.356873, 3.540405, 
    3.61853, 3.868286, 4.0914, 4.138458, 4.186493, 4.543274, 4.786652, 
    4.76236, 4.739258, 4.484558, 3.209167, 2.859833, 2.078125, 1.791779, 
    1.536316, 1.210693, 0.6311951, -0.1725464, -0.6008911, -0.2477722, 
    0.505127, 1.200012, 1.527496, 1.68396, 1.799377, 1.864014,
  2.178253, 1.903442, 2.362946, 2.286438, 2.247589, 2.272949, 2.388855, 
    2.197113, 2.048096, 2.155762, 2.210999, 2.41861, 2.687286, 2.946838, 
    3.202332, 3.125183, 3.149445, 3.66803, 3.842621, 3.704468, 4.026154, 
    4.471069, 4.326538, 3.900314, 3.660202, 3.817307, 4.057419, 4.078842, 
    3.93457, 3.6595, 3.702927, 3.674744, 4.220566, 4.814072, 4.81543, 
    4.599533, 4.653778, 4.757492, 3.953064, 2.475281, 2.448761, 2.622009, 
    3.907227, 2.319855, 2.206512, 2.293427, 2.378448, 2.470428, 2.555237, 
    2.611786, 2.622589, 2.692719, 2.849426, 2.980469, 2.972595, 2.976044, 
    2.930725, 2.829895, 2.660828, 2.434235, 2.241272, 3.101959, 3.718658, 
    3.332916, 2.976105, 2.80011, 2.964203, 3.65976, 3.997864, 3.998962, 
    4.173889, 4.291931, 4.906036, 5.559357, 6.073486, 6.725067, 5.837311, 
    5.423859, 5.247574, 5.122192, 4.64563, 2.535339, 1.992371, 1.560425, 
    1.288666, 1.207825, 0.8551941, 0.05404663, -0.6678467, -0.7058716, 
    -0.007720947, 0.9009399, 1.419037, 1.593658, 2.103638, 2.257996,
  1.447723, 1.725067, 1.926758, 3.113922, 2.898499, 2.16333, 2.067566, 
    2.592743, 2.904541, 2.828033, 2.90448, 2.610413, 2.693604, 2.944641, 
    3.387146, 3.578369, 3.529297, 3.750061, 3.99115, 4.290222, 4.536957, 
    4.5755, 4.676086, 4.389618, 4.24263, 4.058578, 4.22493, 3.64238, 
    3.885345, 3.938477, 3.924103, 4.054749, 4.225708, 4.563293, 4.8069, 
    4.698883, 4.876358, 4.961716, 4.868683, 2.705566, 3.004852, 3.957031, 
    5.237808, 4.767548, 2.965607, 3.028961, 3.018799, 3.085938, 3.261444, 
    3.367432, 3.442383, 3.551056, 3.69516, 3.873779, 5.259888, 3.424194, 
    3.060089, 2.741913, 2.613739, 2.624481, 4.133514, 4.495117, 4.191559, 
    3.906433, 3.621582, 3.8862, 4.043854, 4.309509, 4.038986, 4.421082, 
    5.458313, 6.818726, 9.857941, 9.902069, 9.895477, 10.13318, 7.920624, 
    7.302261, 7.400192, 7.004486, 4.689423, 2.3974, 1.968018, 1.818939, 
    1.744415, 1.479706, 1.223053, 0.8671265, 0.4898376, 0.4300232, 0.7432861, 
    1.175568, 1.472382, 1.57077, 1.543488, 1.980652,
  1.327026, 1.685028, 3.205536, 3.800293, 3.779877, 2.217834, 3.067291, 
    3.019897, 3.082489, 3.203247, 3.292358, 3.364594, 3.391968, 3.708527, 
    4.109436, 4.477722, 4.380646, 4.057587, 4.061829, 4.275558, 4.533966, 
    4.825928, 4.785156, 4.846024, 4.946167, 4.416016, 4.47728, 4.713226, 
    5.199997, 5.244278, 5.105728, 5.107819, 5.475449, 5.839584, 6.384125, 
    6.589844, 6.084824, 5.339188, 5.615555, 5.720764, 6.089325, 6.134506, 
    6.517838, 6.958267, 6.983795, 6.691483, 6.79483, 4.755493, 5.950775, 
    6.346954, 6.663422, 7.184448, 8.652344, 8.667053, 8.187943, 7.352356, 
    6.68631, 5.559296, 4.909821, 4.525574, 4.327728, 4.26326, 4.207535, 
    3.999802, 4.254089, 4.514832, 4.741531, 4.976349, 4.943161, 5.774414, 
    7.340683, 11.11185, 12.02692, 13.26703, 14.5527, 14.23299, 10.06425, 
    10.12259, 13.6395, 12.16281, 7.80722, 4.241089, 3.466644, 4.174286, 
    3.229279, 1.748383, 1.583008, 1.381989, 1.249359, 1.293884, 1.317047, 
    1.174347, 0.8695984, 0.6895142, 0.9963074, 1.204681,
  1.025146, 1.246796, 1.118622, 2.913391, 3.219391, 3.421204, 3.319122, 
    4.303497, 4.742737, 4.98233, 4.775635, 4.296448, 4.220306, 4.382599, 
    4.677322, 4.876862, 4.932007, 4.895309, 5.140427, 5.684128, 6.158325, 
    6.15097, 5.719009, 5.566071, 5.502472, 4.625, 4.417389, 4.521805, 
    4.945831, 5.887573, 6.028259, 5.997589, 6.451233, 7.336075, 6.952606, 
    6.593552, 5.972717, 5.869598, 6.905731, 6.792648, 6.469986, 6.248184, 
    6.463547, 6.712372, 6.93782, 7.002411, 7.3862, 7.807098, 9.242065, 
    11.74197, 13.4055, 17.02238, 11.75259, 8.998627, 6.797562, 5.691772, 
    5.302719, 5.252487, 4.936646, 4.632553, 4.294998, 4.220688, 4.454666, 
    4.662674, 4.648499, 4.500397, 4.915756, 5.885742, 6.780914, 7.091339, 
    6.816208, 6.854568, 7.511063, 8.682816, 10.87439, 10.63585, 9.871796, 
    7.894333, 8.968948, 9.950714, 11.90356, 9.402771, 6.676956, 4.427841, 
    3.160416, 2.949402, 2.950775, 1.652649, 1.929962, 2.124298, 2.308472, 
    4.134308, 1.898163, 1.221985, 0.8719788, 0.7738953,
  1.262848, 1.002075, 0.9157715, 0.8839417, 1.131012, 3.586426, 3.969604, 
    4.16098, 4.236572, 4.106995, 4.102997, 2.580322, 3.154663, 4.829346, 
    5.786652, 6.554352, 6.595428, 6.436829, 6.623703, 6.781769, 6.833984, 
    6.917114, 6.881378, 6.641205, 6.378448, 5.539841, 5.350327, 5.533524, 
    5.409103, 5.643036, 6.049469, 6.388474, 6.639206, 6.812897, 6.675781, 
    6.567001, 7.070709, 6.570374, 7.506897, 7.65892, 7.491806, 7.212036, 
    7.239456, 7.748047, 7.520187, 7.047134, 6.739975, 6.948761, 8.233139, 
    11.12233, 14.76099, 16.37321, 14.79105, 9.262634, 7.22435, 6.339645, 
    6.306381, 6.627014, 5.700653, 6.554626, 6.721298, 6.112747, 6.124542, 
    5.764328, 5.690048, 5.643097, 6.510025, 7.696289, 8.786331, 12.58116, 
    9.002808, 8.300781, 7.85379, 10.06334, 7.419983, 7.806503, 7.21991, 
    8.260605, 9.83197, 12.31483, 13.40831, 11.27992, 6.654953, 4.609756, 
    3.778122, 4.120056, 4.285614, 4.766602, 6.221207, 7.366455, 11.76717, 
    10.92941, 7.409363, 4.48587, 2.911774, 1.936127,
  3.249023, 2.404114, 1.768555, 1.439575, 1.163361, 1.365509, 2.087494, 
    2.85379, 3.349426, 3.579681, 3.698242, 4.198883, 6.080536, 8.970215, 
    10.33182, 9.578247, 10.52077, 10.44717, 9.719955, 8.242249, 7.667191, 
    7.302994, 7.275131, 6.968414, 6.645447, 6.253448, 6.139465, 5.896545, 
    5.965942, 6.725723, 6.600464, 6.924744, 7.07663, 7.356583, 7.517319, 
    7.623566, 7.76413, 7.690964, 7.556183, 7.411591, 7.931183, 8.118225, 
    8.270447, 8.334045, 8.239182, 7.974487, 7.437241, 6.966797, 6.950333, 
    7.346939, 7.879944, 8.261719, 8.391144, 8.190765, 8.004227, 7.778183, 
    7.576889, 7.37233, 7.125336, 6.883865, 6.705078, 6.396362, 5.779556, 
    6.306244, 6.290237, 6.321609, 6.612823, 7.122208, 7.834579, 9.693069, 
    8.310608, 8.101822, 8.4384, 6.79863, 6.644531, 6.671478, 7.637039, 
    8.398499, 9.881317, 10.81386, 9.335281, 6.801361, 5.475266, 4.1315, 
    3.48053, 3.083344, 2.604233, 2.79863, 3.777466, 5.312302, 6.849792, 
    8.961319, 9.735596, 10.31931, 8.77832, 4.682037,
  7.974915, 5.616516, 3.655182, 3.134888, 3.015076, 5.035492, 8.706085, 
    11.56448, 12.45552, 12.74529, 12.58403, 12.20433, 11.81229, 11.33891, 
    10.81627, 10.39796, 10.20526, 9.872177, 9.258835, 8.688675, 8.285095, 
    7.844864, 7.502747, 7.072983, 6.484238, 7.420258, 7.467255, 7.227921, 
    7.419724, 7.734772, 7.731262, 7.665634, 7.790436, 7.910599, 7.902145, 
    7.974472, 8.10051, 8.116135, 8.061722, 8.067184, 8.005661, 7.961533, 
    7.969864, 7.998169, 8.077744, 8.064117, 8.033203, 8.000854, 7.994339, 
    7.988098, 8.075714, 8.290558, 8.442245, 8.510544, 8.510483, 8.38327, 
    8.185867, 8.011917, 7.827011, 7.703186, 7.70546, 7.765167, 7.770767, 
    7.547394, 6.995956, 7.623566, 7.527222, 7.439072, 7.355408, 7.2845, 
    7.08197, 7.190887, 6.882813, 6.491928, 5.869202, 5.987564, 5.728592, 
    6.159439, 4.698044, 4.483795, 4.216736, 4.027802, 4.161453, 4.721558, 
    5.04303, 4.649536, 4.319199, 4.316864, 4.620834, 5.24617, 6.350647, 
    7.480667, 8.564301, 9.182999, 9.231888, 8.681473,
  8.091461, 7.653305, 7.134109, 6.378189, 8.338593, 8.713593, 9.08989, 
    9.763916, 9.993927, 10.20584, 10.24348, 10.10043, 9.849396, 9.565735, 
    9.272324, 9.002533, 8.779221, 8.594971, 8.480988, 8.403839, 8.294205, 
    8.126755, 7.941727, 7.667191, 7.228638, 7.587311, 7.488159, 7.359573, 
    7.436005, 7.516479, 7.467575, 7.464523, 7.525909, 7.631119, 7.730789, 
    7.766998, 7.820709, 7.817719, 7.780334, 7.748383, 7.686203, 7.61055, 
    7.61113, 7.692581, 7.856644, 8.066544, 8.251236, 8.426239, 8.540939, 
    8.573318, 8.630997, 8.69133, 8.657227, 8.53717, 8.460938, 8.415619, 
    8.354874, 8.368423, 8.424927, 8.535019, 8.684509, 8.86647, 8.931, 
    8.984253, 9.012039, 9.074997, 8.877075, 8.560211, 8.171356, 7.6698, 
    7.127533, 6.979172, 6.474609, 6.311081, 5.766724, 5.219925, 4.712173, 
    4.399994, 4.198502, 4.0513, 4.018097, 4.011002, 3.912308, 3.740311, 
    3.658844, 3.786972, 4.072464, 4.482224, 5.07605, 5.919983, 6.719193, 
    7.445572, 8.255936, 8.485153, 8.516327, 8.377518,
  8.881363, 8.858566, 8.851685, 8.794632, 8.820236, 8.851089, 8.8759, 
    8.895615, 8.898422, 8.922775, 8.927063, 8.929611, 8.916397, 8.900894, 
    8.897507, 8.87616, 8.836838, 8.782349, 8.739975, 8.673691, 8.571808, 
    8.456451, 8.290298, 8.142838, 7.98645, 7.918823, 7.877594, 7.775589, 
    7.657166, 7.57428, 7.503189, 7.467194, 7.448303, 7.478134, 7.539322, 
    7.593811, 7.649994, 7.729492, 7.804489, 7.874863, 7.93782, 7.997711, 
    8.085022, 8.132156, 8.164642, 8.225388, 8.256393, 8.289658, 8.330536, 
    8.384705, 8.389587, 8.40535, 8.404816, 8.405731, 8.405731, 8.468811, 
    8.548309, 8.648117, 8.763855, 8.872452, 8.960297, 9.068161, 9.090439, 
    9.105789, 9.134567, 9.155014, 9.109894, 9.1194, 9.050842, 8.980927, 
    8.823242, 8.72818, 8.605286, 8.505478, 8.213669, 8.068817, 7.98111, 
    7.99733, 8.007675, 7.870499, 7.935165, 7.783142, 7.808792, 7.822647, 
    7.997528, 8.274933, 8.550903, 8.686707, 8.864899, 8.862686, 8.905914, 
    8.924088, 8.995911, 9.031448, 8.953125, 8.893875,
  8.57988, 8.525848, 8.583008, 8.607285, 8.588806, 8.561066, 8.524933, 
    8.46048, 8.430603, 8.427795, 8.380142, 8.316208, 8.231369, 8.155136, 
    8.099792, 8.091797, 8.047913, 7.947525, 7.885818, 7.862564, 7.86348, 
    7.840164, 7.773239, 7.713547, 7.670898, 7.634903, 7.582031, 7.541916, 
    7.524673, 7.506699, 7.526962, 7.572128, 7.597, 7.621689, 7.624557, 
    7.635162, 7.672455, 7.710403, 7.738998, 7.757034, 7.758926, 7.799927, 
    7.855011, 7.908661, 7.948441, 8.004807, 8.074417, 8.155731, 8.19368, 
    8.201813, 8.224609, 8.263275, 8.300201, 8.352341, 8.406448, 8.410477, 
    8.45372, 8.504166, 8.580673, 8.652344, 8.703323, 8.755463, 8.827805, 
    8.906708, 8.981308, 9.031311, 9.083389, 9.128571, 9.160156, 9.166733, 
    9.193878, 9.160675, 9.144455, 9.15007, 9.172989, 9.19577, 9.172333, 
    9.137238, 9.128906, 9.111191, 9.073181, 8.995239, 8.952988, 8.945114, 
    8.947266, 8.925186, 8.88913, 8.879883, 8.847855, 8.784958, 8.754044, 
    8.711075, 8.676941, 8.642776, 8.629684, 8.575455 ;
}
