netcdf CGMR_SRA1B_1_huss-change_2070-2099 {
dimensions:
	time = 12 ;
	latitude = 48 ;
	longitude = 96 ;
	bounds = 2 ;
data:
 specific_humidity_anomaly =
  0.0001414621, 0.0001357719, 0.0001307651, 0.0001265212, 0.0001230245, 
    0.000120354, 0.0001184149, 0.0001170956, 0.0001164918, 0.0001163805, 
    0.0001171594, 0.000118415, 0.0001203859, 0.0001226112, 0.0001250272, 
    0.0001274749, 0.0001300181, 0.0001325294, 0.0001351202, 0.0001375839, 
    0.0001397138, 0.0001418436, 0.0001434967, 0.0001448318, 0.0001458173, 
    0.000146612, 0.0001471842, 0.0001475339, 0.0001477087, 0.0001477246, 
    0.0001476769, 0.0001476451, 0.0001478198, 0.0001481854, 0.0001485828, 
    0.0001491549, 0.0001501246, 0.0001515074, 0.0001535102, 0.0001558467, 
    0.000158517, 0.0001611237, 0.0001641437, 0.0001675928, 0.000170867, 
    0.0001739823, 0.0001770659, 0.0001804038, 0.0001835032, 0.0001863166, 
    0.000188367, 0.0001899406, 0.00019002, 0.0001891617, 0.0001887485, 
    0.0001870636, 0.000184902, 0.0001819615, 0.0001783217, 0.0001748248, 
    0.0001710419, 0.0001670683, 0.0001642073, 0.0001604084, 0.0001574521, 
    0.0001554334, 0.0001537486, 0.0001529697, 0.0001534784, 0.0001551791, 
    0.0001574202, 0.0001604243, 0.0001635078, 0.0001656695, 0.0001724565, 
    0.0001777494, 0.0001819932, 0.0001863007, 0.0001925471, 0.0001969975, 
    0.000200399, 0.0002030216, 0.0002043726, 0.0002048336, 0.0002041183, 
    0.0002024017, 0.0001994136, 0.0001953922, 0.0001907671, 0.0001851245, 
    0.0001793547, 0.0001730605, 0.0001668457, 0.0001603608, 0.0001538758, 
    0.0001475815,
  0.0001788144, 0.0001656695, 0.0001541937, 0.0001440211, 0.000134246, 
    0.0001249636, 0.0001163644, 0.0001081152, 0.0001003905, 9.357178e-005, 
    8.861269e-005, 8.54019e-005, 8.468665e-005, 8.554498e-005, 8.846959e-005, 
    9.328566e-005, 9.946869e-005, 0.0001064623, 0.0001136943, 0.0001200044, 
    0.0001242484, 0.0001264418, 0.0001262352, 0.0001236761, 0.0001188601, 
    0.0001124705, 0.000106351, 0.0001006449, 9.684602e-005, 9.45731e-005, 
    9.500227e-005, 9.764076e-005, 0.0001029972, 0.0001102768, 0.0001200045, 
    0.0001316711, 0.0001447204, 0.0001583103, 0.0001714392, 0.0001836145, 
    0.0001936598, 0.0002038483, 0.0002138776, 0.0002250039, 0.0002344932, 
    0.0002456987, 0.0002584303, 0.0002750242, 0.0002916498, 0.0003108823, 
    0.0003283027, 0.000346184, 0.0003631593, 0.0003758275, 0.0003859047, 
    0.0003880187, 0.0003866517, 0.0003843311, 0.000375303, 0.0003600918, 
    0.0003425602, 0.0003212297, 0.0002969586, 0.0002740386, 0.0002531852, 
    0.0002350969, 0.0002188685, 0.0002100154, 0.0002098088, 0.0002151175, 
    0.000225735, 0.0002373382, 0.0002515479, 0.0002701285, 0.0002878351, 
    0.0003059867, 0.0003220403, 0.0003354236, 0.0003451827, 0.000351191, 
    0.0003538611, 0.0003508254, 0.0003486638, 0.0003401919, 0.000336107, 
    0.0003273967, 0.0003178599, 0.0003063205, 0.0002942883, 0.0002807143, 
    0.0002664569, 0.000250928, 0.0002359076, 0.0002216342, 0.0002073291, 
    0.0001928332,
  0.0001355652, 0.0001207356, 0.0001100386, 0.000103474, 0.0001017416, 
    0.0001047457, 0.0001105631, 0.0001178746, 0.0001241847, 0.0001269981, 
    0.000126251, 0.0001225635, 0.0001159355, 0.0001090849, 0.0001030291, 
    0.0001006131, 0.000103188, 0.000109816, 0.0001171434, 0.0001240734, 
    0.0001281266, 0.0001286034, 0.0001253768, 0.0001180494, 0.0001086557, 
    0.0001010581, 9.652812e-005, 9.524068e-005, 9.714806e-005, 0.0001030926, 
    0.0001117552, 0.0001237238, 0.0001379493, 0.0001533512, 0.0001702948, 
    0.0001877948, 0.0002063597, 0.0002253537, 0.0002458895, 0.0002677285, 
    0.0002889319, 0.0003059867, 0.0003198627, 0.0003275875, 0.0003298763, 
    0.000331418, 0.0003292883, 0.0003252194, 0.0003250603, 0.0003186706, 
    0.0003102308, 0.0003036025, 0.0002992952, 0.0003003124, 0.0003006142, 
    0.0003056212, 0.0003170811, 0.0003313546, 0.0003481392, 0.0003645108, 
    0.0003763522, 0.0003782593, 0.0003734115, 0.0003680233, 0.0003527963, 
    0.0003322287, 0.0003095471, 0.0002934937, 0.0002810005, 0.0002802534, 
    0.0002857053, 0.0002964659, 0.0003055576, 0.0003112321, 0.000313346, 
    0.0003126308, 0.0003033006, 0.0002929374, 0.0002826694, 0.000272481, 
    0.0002632146, 0.0002530739, 0.0002538527, 0.0002598767, 0.0002712732, 
    0.0002803172, 0.0002880259, 0.0002944949, 0.0002936685, 0.0002871039, 
    0.0002770905, 0.0002581282, 0.000235383, 0.0002096021, 0.0001831534, 
    0.0001574203,
  0.0001617436, 0.0001313691, 0.000107257, 8.867623e-005, 7.500692e-005, 
    6.922119e-005, 7.336965e-005, 8.610124e-005, 0.0001037125, 0.0001216257, 
    0.0001338327, 0.0001377269, 0.0001361056, 0.0001329267, 0.0001297637, 
    0.0001337214, 0.000143719, 0.0001567526, 0.0001667821, 0.0001682763, 
    0.0001643344, 0.000154575, 0.0001404767, 0.0001233105, 0.0001101497, 
    0.0001017573, 0.0001014712, 0.0001085604, 0.0001200999, 0.0001318459, 
    0.0001423045, 0.000150077, 0.0001525724, 0.0001492187, 0.0001418118, 
    0.0001325135, 0.0001258854, 0.0001268231, 0.0001353585, 0.0001550837, 
    0.0001836622, 0.0002151653, 0.0002479716, 0.0002750241, 0.0002913319, 
    0.0003008846, 0.0002625943, 0.0002484482, 0.0002637866, 0.0002786799, 
    0.0002820813, 0.0002742929, 0.0002598607, 0.0002367974, 0.0002287391, 
    0.0002211733, 0.0002137981, 0.0002704624, 0.0003009797, 0.0003278577, 
    0.0003490929, 0.0003682141, 0.0003773377, 0.0003757799, 0.0003627146, 
    0.0003509048, 0.0003401601, 0.0003362501, 0.000338364, 0.0003398899, 
    0.0003389204, 0.0003344063, 0.0003262365, 0.0003173992, 0.000307465, 
    0.0002985641, 0.0002879306, 0.0002903148, 0.0003025059, 0.0003135526, 
    0.0003335795, 0.0003553075, 0.0003697078, 0.0003821536, 0.0004015923, 
    0.000411622, 0.0004096511, 0.000407696, 0.000398922, 0.0004001464, 
    0.0003906097, 0.0003643517, 0.000326904, 0.0002796494, 0.0002335712, 
    0.0001935167,
  0.0002244159, 0.0002168184, 0.0002165321, 0.0002129399, 0.0002059464, 
    0.0001921817, 0.0001844727, 0.000186857, 0.0001975539, 0.0002043727, 
    0.0002014958, 0.0001869682, 0.0001662416, 0.0001551632, 0.0001581196, 
    0.0001735372, 0.0001967752, 0.000217454, 0.0002306147, 0.0002277854, 
    0.0002169932, 0.0002012097, 0.0001768117, 0.0001486305, 0.0001248205, 
    0.0001105312, 0.000105445, 0.0001085126, 0.0001102927, 0.0001120095, 
    0.0001144891, 0.0001245185, 0.0001433377, 0.0001665438, 0.0001898611, 
    0.0002085213, 0.0002193932, 0.0002261802, 0.0002395157, 0.0002585416, 
    0.0002810482, 0.0002994699, 0.0003040794, 0.0003000104, 0.0002896949, 
    0.0002780919, 0.0002406917, 0.000209745, 0.0001632851, 0.0001195909, 
    9.412807e-005, 8.180947e-005, 8.166651e-005, 8.859648e-005, 0.0001002632, 
    0.0001197974, 0.0001458011, 0.0001701517, 0.0002065978, 0.000237783, 
    0.0002578259, 0.0002588753, 0.0002498154, 0.0002340479, 0.0002207758, 
    0.0002068363, 0.0001790845, 0.0001565616, 0.0001619181, 0.0001774472, 
    0.0002475423, 0.0002447448, 0.0002354623, 0.0002030374, 0.0001679901, 
    0.000149902, 0.0002296928, 0.0002413911, 0.000254679, 0.000270081, 
    0.0002811435, 0.0002804124, 0.0002759141, 0.0002701445, 0.0002687934, 
    0.000267013, 0.0002663934, 0.0002714796, 0.0002869291, 0.0003099602, 
    0.0003393018, 0.0003371402, 0.0003393337, 0.0003209276, 0.0002791884, 
    0.0002434575,
  0.0001352313, 0.0001262508, 0.0001706127, 0.000199652, 0.0002229855, 
    0.0002364005, 0.000255474, 0.0002849107, 0.0003161276, 0.0003335797, 
    0.0003383481, 0.0003205939, 0.0002901399, 0.0002560776, 0.000240517, 
    0.0002425198, 0.0002409304, 0.0002287549, 0.0002058034, 0.0001767164, 
    0.0001847271, 0.0002173587, 0.0002313142, 0.0002262439, 0.0002137983, 
    0.0002006692, 0.0002065661, 0.0002260528, 0.00024821, 0.0002559506, 
    0.0002455397, 0.0002220635, 0.0002026878, 0.0002028947, 0.000210969, 
    0.0002126537, 0.000200431, 0.0001796408, 0.0001649066, 0.0001717093, 
    0.0002006853, 0.0002195999, 0.0002176128, 0.000194629, 0.0001490593, 
    0.0001217686, 0.0001258217, 0.0001212442, 8.961395e-005, 5.664839e-005, 
    3.821077e-005, 5.302462e-005, 7.920293e-005, 9.454135e-005, 
    9.164866e-005, 9.044027e-005, 9.738631e-005, 0.0001157604, 0.0001377268, 
    0.0001379494, 0.0001224519, 0.0001135671, 0.0001157606, 0.0001253129, 
    0.0001267276, 0.0001190985, 0.00010589, 0.0001136782, 0.0001255993, 
    0.000128492, 0.0001163008, 9.323796e-005, 9.915046e-005, 0.0001068912, 
    0.0001198612, 0.000122007, 0.0001389189, 0.000171137, 0.000300074, 
    0.0003375851, 0.0003217859, 0.000313902, 0.0002902353, 0.0002766135, 
    0.000280587, 0.0002883754, 0.0002952099, 0.0002947175, 0.0003005667, 
    0.0003219766, 0.0003483614, 0.0003621103, 0.0003595355, 0.0003201487, 
    0.000246366, 0.0001738868,
  0.0002482892, 0.000269461, 0.0002928101, 0.0003148399, 0.0003308298, 
    0.0003483456, 0.0003539722, 0.0003488702, 0.0003322763, 0.0003124715, 
    0.0003077034, 0.0003126941, 0.0003115817, 0.0003174786, 0.0003304642, 
    0.0003216271, 0.0002878509, 0.0002408505, 0.0001686735, 0.0001085284, 
    7.843995e-005, 8.314475e-005, 0.000111755, 0.000128953, 0.0001219434, 
    0.0001099908, 9.924592e-005, 0.0001046341, 0.0001211963, 0.0001420183, 
    0.0001783532, 0.0001709464, 0.0001623633, 0.0002166433, 0.0002196315, 
    0.0002292634, 0.0002436005, 0.0002050402, 0.0001781147, 0.0001545113, 
    9.409594e-005, 9.945268e-005, 0.0001186372, 0.0001094344, 6.388081e-005, 
    2.64491e-005, -6.182352e-006, -2.787844e-005, -4.316936e-005, 
    -4.440895e-005, -2.884818e-005, 6.596558e-006, 2.614711e-005, 
    1.886743e-005, -1.223525e-006, -1.430046e-006, 5.275453e-005, 
    0.0001166826, 0.0001580087, 0.0001930245, 0.0002239554, 0.0002595112, 
    0.0003009641, 0.000321198, 0.0003079739, 0.0002933347, 0.0002862937, 
    0.0002960847, 0.0003167796, 0.0003251876, 0.0003348989, 0.0003398899, 
    0.0003530192, 0.0003584865, 0.0003570244, 0.0003372994, 0.0003115342, 
    0.0003016638, 0.0003533368, 0.0003869063, 0.0002734826, 0.0001774156, 
    0.0001181446, 0.0001098316, 0.0001349451, 0.0001409214, 0.0001422884, 
    0.0001514435, 0.0001593432, 0.0001698972, 0.0001773043, 0.0001886368, 
    0.000208219, 0.0002309007, 0.0002442838, 0.0002470496,
  0.0002879305, 0.0002920949, 0.0002933822, 0.0002847833, 0.0002873901, 
    0.0003180986, 0.0003630642, 0.0003906572, 0.0003942016, 0.0004064725, 
    0.0004422513, 0.0004769808, 0.0004950052, 0.0004731978, 0.0004446513, 
    0.0004256892, 0.0004119403, 0.0004017199, 0.0003746992, 0.0003296381, 
    0.0002882008, 0.0002695087, 0.000271146, 0.0002832417, 0.0002876287, 
    0.0002686821, 0.0002201085, 0.0001813418, 0.0001667347, 0.0001751746, 
    0.0001836619, 0.000201846, 0.0002292166, 0.0002562851, 0.0002783467, 
    0.0003037304, 0.0003183214, 0.0003003287, 0.0002751038, 0.0002605449, 
    0.0002337936, 0.0002083941, 0.0002145772, 0.0002411697, 0.0002411217, 
    0.0001834566, 5.633058e-005, -3.263075e-005, -4.614145e-005, 
    -7.176353e-005, -0.0001129941, -0.0001379326, -0.0001431778, 
    -0.0001478349, -0.0001159506, -3.840122e-005, 5.579041e-005, 
    0.0001376793, 0.0001751431, 0.000222445, 0.0003086417, 0.0003890684, 
    0.0004478944, 0.0004895059, 0.0005038427, 0.0005033663, 0.0005121082, 
    0.0005253642, 0.0005287342, 0.0005443422, 0.0005956497, 0.0006395192, 
    0.0006594509, 0.0006589899, 0.000657957, 0.0006610872, 0.0006431113, 
    0.0005900552, 0.00053471, 0.0004867562, 0.0004451121, 0.0003938205, 
    0.0003007578, 0.0002744682, 0.0003077511, 0.0003380941, 0.0003571038, 
    0.0003686273, 0.0003638589, 0.0003500625, 0.0003302579, 0.0003183845, 
    0.0003161435, 0.0003228828, 0.0003087204, 0.0002942565,
  0.0003684368, 0.000349252, 0.0003379828, 0.00032452, 0.0003067658, 
    0.000300122, 0.0003238681, 0.0003512546, 0.0003682622, 0.000385317, 
    0.0004037227, 0.0004250691, 0.0004273425, 0.0004349239, 0.0004546177, 
    0.0004612301, 0.0004533459, 0.0004556668, 0.0004501194, 0.0004212386, 
    0.0003872081, 0.000347456, 0.0003185119, 0.0003163824, 0.0003281282, 
    0.0003426247, 0.0003473926, 0.000347266, 0.000337983, 0.0003223429, 
    0.0003023474, 0.0002698274, 0.0002450314, 0.0002434258, 0.0002449835, 
    0.0002509593, 0.0002844972, 0.0003521121, 0.0004013223, 0.0004109866, 
    0.0003892584, 0.0003786725, 0.0004229546, 0.0004315535, 0.0004265783, 
    0.0004090145, 0.0003248528, 0.0001491071, -2.950057e-005, -0.000143433, 
    -0.0002030851, -0.0002004784, -0.0001610913, -0.0001473585, 
    -0.0001379009, -7.929746e-005, 1.104688e-005, 6.56452e-005, 
    6.340398e-005, 0.000155862, 0.0003419877, 0.0004631202, 0.000525252, 
    0.0006192843, 0.000702254, 0.0007276535, 0.0007341383, 0.0007600146, 
    0.0007802485, 0.0008008, 0.0008247532, 0.000841077, 0.0008257702, 
    0.0007886561, 0.0007689153, 0.0007374757, 0.0006407094, 0.000584315, 
    0.0005956795, 0.0006134505, 0.0006149611, 0.0005804538, 0.0004840861, 
    0.0003490616, 0.0002828287, 0.0003037457, 0.0003505554, 0.0003895606, 
    0.0004048832, 0.0004125445, 0.0004344787, 0.0004416311, 0.0004262291, 
    0.0004103505, 0.0004041041, 0.0003974917,
  0.0004428397, 0.0004360368, 0.0004807957, 0.0005193879, 0.0005079275, 
    0.0004943698, 0.0005112342, 0.0005294336, 0.0005501756, 0.0005579004, 
    0.0005446603, 0.0005316585, 0.0005266997, 0.0005494445, 0.0005869078, 
    0.0006045033, 0.0006374205, 0.0007003783, 0.0006879009, 0.0005311333, 
    0.0004181713, 0.0003722515, 0.0003475673, 0.0003523189, 0.000390959, 
    0.000458193, 0.0004984061, 0.00048817, 0.0004726411, 0.0004796823, 
    0.0004913649, 0.0004638676, 0.0004443484, 0.0004200609, 0.0004036734, 
    0.0004153084, 0.0004803329, 0.0005812952, 0.0006240201, 0.0005939952, 
    0.0005562138, 0.0005760025, 0.0006090156, 0.0005703438, 0.0005485681, 
    0.0005683415, 0.0005600601, 0.0004211096, 0.0002226182, 0.0001336406, 
    0.0001152824, 0.0001467853, 0.0001606774, 0.0001678937, 0.0001677186, 
    0.0001794966, 0.0002223961, 0.0002531204, 0.0002681403, 0.0003431467, 
    0.000485213, 0.0005896715, 0.0006455253, 0.0007256339, 0.0008002748, 
    0.0007930584, 0.0007824888, 0.0008283765, 0.0008598953, 0.0008495483, 
    0.0008481811, 0.0008583535, 0.0008497229, 0.0008117827, 0.000766451, 
    0.0006606253, 0.0006225575, 0.0006636293, 0.0007266672, 0.000761556, 
    0.0007695509, 0.0006711315, 0.0005096756, 0.0003707889, 0.0003767489, 
    0.0004443647, 0.0005325796, 0.0005775304, 0.0005749236, 0.0005799462, 
    0.0005834908, 0.0005774032, 0.0005388903, 0.0004932731, 0.0004786504, 
    0.0004725782,
  0.0006270888, 0.0006902856, 0.0007845564, 0.0008260407, 0.0008344492, 
    0.0008420628, 0.0008454481, 0.0008438746, 0.0008608503, 0.0008776663, 
    0.0008917651, 0.0008891425, 0.0008838652, 0.000894737, 0.0008836747, 
    0.0008586245, 0.0008879025, 0.0009652451, 0.0009772773, 0.0008735657, 
    0.0008188877, 0.0008147554, 0.0007668328, 0.0006992649, 0.0006790152, 
    0.0007057977, 0.0007541645, 0.0007658945, 0.0007478227, 0.0007234723, 
    0.0007097078, 0.0006886311, 0.0006562858, 0.0006206026, 0.0005954891, 
    0.0005915794, 0.0006343038, 0.0006964831, 0.0007401616, 0.0007883534, 
    0.0008568112, 0.0009080875, 0.0008942434, 0.0008409177, 0.0008275025, 
    0.0008290755, 0.0007546567, 0.0006146254, 0.0004820018, 0.0004534069, 
    0.0004904568, 0.0005399375, 0.0005511423, 0.0005532247, 0.0005487748, 
    0.0005748891, 0.0005905931, 0.000638213, 0.0006754068, 0.0007035881, 
    0.0007681986, 0.0008348292, 0.000855031, 0.0008623111, 0.0008845483, 
    0.0008867886, 0.0008867891, 0.0008915416, 0.0008789371, 0.000843476, 
    0.0008206195, 0.0008169482, 0.0007936945, 0.0007626363, 0.0006994391, 
    0.0006791735, 0.0007243943, 0.0007335651, 0.00084311, 0.000938986, 
    0.0009242832, 0.0007686289, 0.0005745399, 0.000495004, 0.000530703, 
    0.0006288518, 0.0007156366, 0.0007835063, 0.0008113063, 0.0008147713, 
    0.0008031684, 0.0007800739, 0.0007418315, 0.0006964845, 0.0006568432, 
    0.0006244183,
  0.0008856445, 0.0009450424, 0.0009958893, 0.00104111, 0.001104417, 
    0.001176452, 0.001264698, 0.001318836, 0.001329564, 0.001321585, 
    0.001329517, 0.001346476, 0.001343106, 0.00129876, 0.001243289, 
    0.001207843, 0.001209401, 0.001228188, 0.001221735, 0.001271676, 
    0.001389216, 0.001397243, 0.001296106, 0.001213804, 0.001161447, 
    0.001134967, 0.001115655, 0.001058117, 0.0009701559, 0.0009144447, 
    0.000927892, 0.0009370162, 0.0008648708, 0.000791755, 0.0007812334, 
    0.0008051693, 0.0008580508, 0.0009098668, 0.0009262068, 0.0009793574, 
    0.001094275, 0.001139351, 0.001146584, 0.001133693, 0.001143405, 
    0.001151717, 0.001126143, 0.001032556, 0.0009090072, 0.0008837199, 
    0.0009470433, 0.001014548, 0.00101272, 0.000939779, 0.0009024758, 
    0.0009141732, 0.0009407653, 0.001000639, 0.001048069, 0.001057606, 
    0.001058862, 0.001077222, 0.001071435, 0.0010344, 0.001048881, 
    0.001048833, 0.001002517, 0.000957503, 0.0009225989, 0.0008431096, 
    0.0007771626, 0.0007516043, 0.0007522078, 0.0007321658, 0.0007265871, 
    0.0007715048, 0.0008392008, 0.0008315863, 0.000743595, 0.001043302, 
    0.001054015, 0.0009555966, 0.0009030011, 0.0009150808, 0.0009824731, 
    0.001048548, 0.001078795, 0.001065031, 0.001041268, 0.001041761, 
    0.001022131, 0.0009923289, 0.0009534028, 0.0009032716, 0.0008687642, 
    0.0008545546,
  0.001200149, 0.001256512, 0.00134239, 0.001436581, 0.001547429, 
    0.001698379, 0.001897936, 0.002064686, 0.002192289, 0.002269933, 
    0.002303677, 0.00228899, 0.00211682, 0.001897364, 0.001763755, 
    0.00171871, 0.001695026, 0.001672281, 0.001672583, 0.001697714, 
    0.001669612, 0.001574673, 0.001448835, 0.001359652, 0.001299044, 
    0.001282689, 0.001261803, 0.00121795, 0.001201214, 0.001197606, 
    0.001159539, 0.001157822, 0.001158362, 0.001128274, 0.001132311, 
    0.001139639, 0.001145313, 0.001130627, 0.001113938, 0.001242001, 
    0.001509983, 0.001581032, 0.001546079, 0.001554789, 0.001601249, 
    0.001627634, 0.001600565, 0.001457643, 0.001537736, 0.0015868, 
    0.001601789, 0.001561021, 0.001465129, 0.001302543, 0.001252348, 
    0.001247437, 0.001266001, 0.00127309, 0.001269323, 0.001262901, 
    0.001230031, 0.001216871, 0.001225135, 0.001244718, 0.001258148, 
    0.001207413, 0.001114668, 0.001055747, 0.001000084, 0.0009349966, 
    0.0009188317, 0.0009149527, 0.0009038271, 0.0008831481, 0.0008452078, 
    0.0008309344, 0.000929242, 0.0008518677, 0.0006326502, 0.001100379, 
    0.001172716, 0.001160667, 0.001267828, 0.001411785, 0.00144545, 
    0.001414169, 0.001355232, 0.00127223, 0.001243653, 0.001250774, 
    0.001252696, 0.001232145, 0.001189595, 0.001169982, 0.001172699, 
    0.00117146,
  0.00136407, 0.001396209, 0.001459993, 0.001525718, 0.001661188, 
    0.001943206, 0.002148198, 0.002426512, 0.002680778, 0.002750204, 
    0.002609489, 0.002376555, 0.002138613, 0.001948673, 0.001807369, 
    0.001743093, 0.001697588, 0.001619004, 0.001555219, 0.001511303, 
    0.001433642, 0.001391282, 0.001390838, 0.001364882, 0.001322396, 
    0.001335047, 0.001332536, 0.001291528, 0.001296328, 0.001339992, 
    0.001364723, 0.001352135, 0.001331153, 0.001256608, 0.001290496, 
    0.001327435, 0.001318676, 0.001381221, 0.001302353, 0.001963263, 
    0.00187009, 0.002306746, 0.002324866, 0.002240387, 0.002216322, 
    0.002095635, 0.001941855, 0.002112038, 0.00186208, 0.001845629, 
    0.001728645, 0.001627618, 0.001579745, 0.001527483, 0.001478306, 
    0.0014376, 0.00143922, 0.00146427, 0.001450713, 0.001422452, 0.001406335, 
    0.001390917, 0.00139381, 0.001399992, 0.001421737, 0.001391076, 
    0.001338767, 0.001304355, 0.001219049, 0.001139591, 0.001110377, 
    0.001096215, 0.001025627, 0.000959537, 0.0009318646, 0.0009319773, 
    0.0009695683, 0.0009478703, 0.001252409, 0.001802316, 0.001475191, 
    0.001493135, 0.001641144, 0.001831832, 0.001859981, 0.001768732, 
    0.001710795, 0.001672314, 0.001660155, 0.001603729, 0.001525385, 
    0.001514609, 0.001461934, 0.00139114, 0.001357808, 0.001345315,
  0.001501719, 0.001445785, 0.001450013, 0.00156846, 0.001847759, 
    0.002115614, 0.002460366, 0.002798857, 0.002856332, 0.002695701, 
    0.002238002, 0.002008436, 0.001933224, 0.001885111, 0.00182371, 
    0.00174961, 0.001659805, 0.001576295, 0.00148595, 0.001496012, 
    0.001481358, 0.001417779, 0.001369571, 0.001363976, 0.001364071, 
    0.001382366, 0.001426394, 0.001502767, 0.001536496, 0.001640636, 
    0.001683313, 0.001660028, 0.001639032, 0.00152548, 0.001520584, 
    0.001534319, 0.001370683, 0.001976696, 0.002177031, 0.002881398, 
    0.002987986, 0.0030313, 0.003050563, 0.002676724, 0.002496241, 
    0.00234041, 0.002129299, 0.00199855, 0.001831657, 0.001669135, 
    0.001543123, 0.001498253, 0.001518296, 0.001492658, 0.001489114, 
    0.00149989, 0.001538435, 0.001612615, 0.001610183, 0.001614554, 
    0.001598882, 0.001586054, 0.001620625, 0.001600805, 0.001582415, 
    0.001474252, 0.001384957, 0.001346142, 0.001257324, 0.001181872, 
    0.00110162, 0.001061581, 0.001051488, 0.001022115, 0.0009414507, 
    0.0009123152, 0.0009644497, 0.001526307, 0.001847774, 0.001951613, 
    0.002019118, 0.002324723, 0.002118903, 0.002363998, 0.002407565, 
    0.002238462, 0.002139949, 0.002064259, 0.001979875, 0.001901085, 
    0.001782781, 0.00174268, 0.001671774, 0.001624361, 0.001605526, 
    0.001571003,
  0.001549466, 0.001505867, 0.001488478, 0.001684807, 0.001958783, 
    0.001881582, 0.002520766, 0.003661901, 0.003375385, 0.002776368, 
    0.002492714, 0.002583678, 0.002648511, 0.002548978, 0.00238598, 
    0.002214859, 0.002130713, 0.002075369, 0.0020109, 0.001998121, 
    0.001985992, 0.001927437, 0.001876734, 0.001823869, 0.001816716, 
    0.001803429, 0.001849586, 0.001965173, 0.001934592, 0.001897476, 
    0.001955491, 0.002462052, 0.001939661, 0.001561021, 0.001340244, 
    0.00141204, 0.001874843, 0.001961324, 0.002142572, 0.003049198, 
    0.003480115, 0.002677296, 0.002230261, 0.002088051, 0.002194068, 
    0.002166301, 0.002050716, 0.001850635, 0.00172022, 0.001712495, 
    0.001686793, 0.001685379, 0.001758367, 0.001763214, 0.00173141, 
    0.001751596, 0.001795083, 0.001836091, 0.001819291, 0.001859821, 
    0.001870233, 0.001830878, 0.001804016, 0.001701289, 0.001599294, 
    0.001423182, 0.001305943, 0.00117672, 0.001065586, 0.001033003, 
    0.0009552157, 0.0009860024, 0.0009792, 0.0009534983, 0.0008646958, 
    0.0009041782, 0.001043557, 0.001423628, 0.002068868, 0.002601987, 
    0.003007711, 0.003293941, 0.003114508, 0.002805645, 0.002839897, 
    0.002671447, 0.002610411, 0.002466964, 0.002334592, 0.002284287, 
    0.002154746, 0.002014842, 0.001901085, 0.001832578, 0.001742949, 
    0.001633245,
  0.001558667, 0.001549099, 0.00164418, 0.001879738, 0.002353317, 
    0.002522896, 0.003469479, 0.003509837, 0.0029874, 0.002550442, 
    0.002723141, 0.002977069, 0.00306516, 0.002967186, 0.002778608, 
    0.002615102, 0.002537552, 0.002463005, 0.00240933, 0.002400333, 
    0.002333003, 0.002287052, 0.002232105, 0.002163997, 0.00212046, 
    0.002067755, 0.002047013, 0.002119857, 0.002169766, 0.002359327, 
    0.002808157, 0.002969455, 0.002744291, 0.00134684, 0.0002392931, 
    0.0008212081, 0.001353214, 0.001906838, 0.002868109, 0.003340227, 
    0.003279478, 0.002293061, 0.001928344, 0.002040623, 0.002207198, 
    0.002260715, 0.002233964, 0.00215624, 0.002138057, 0.002226223, 
    0.002278342, 0.002227464, 0.00218663, 0.002153807, 0.002128696, 
    0.002114216, 0.002111163, 0.002132953, 0.002105408, 0.002075178, 
    0.001989712, 0.001891993, 0.00177841, 0.001564962, 0.001401756, 
    0.001213214, 0.001167263, 0.001071339, 0.0009996546, 0.001035959, 
    0.0009666588, 0.001032525, 0.0009346958, 0.0009674542, 0.0009293072, 
    0.001024706, 0.001245418, 0.0006744061, 0.003124808, 0.003319563, 
    0.003555397, 0.003583528, 0.003438934, 0.003288046, 0.00313214, 
    0.002961559, 0.0027606, 0.002603101, 0.002514759, 0.002403528, 
    0.002277039, 0.002149501, 0.002013268, 0.001859044, 0.001716198, 
    0.00162091,
  0.001652907, 0.001764693, 0.002017639, 0.002427814, 0.003007744, 
    0.003988073, 0.003710539, 0.003340243, 0.00266342, 0.002693016, 
    0.003064489, 0.003286568, 0.003306676, 0.003026931, 0.002751254, 
    0.002594678, 0.002484767, 0.002436018, 0.002398854, 0.002375873, 
    0.00231269, 0.002292362, 0.002282777, 0.002276195, 0.00222991, 
    0.002243835, 0.002333989, 0.002506129, 0.00260132, 0.002818424, 
    0.003291626, 0.003277697, 0.002441342, 0.0004584938, 0.0002919994, 
    0.001240617, 0.001623199, 0.002593087, 0.003226073, 0.003338034, 
    0.002640406, 0.002349392, 0.002500739, 0.002777115, 0.002805136, 
    0.002740826, 0.002692873, 0.002691267, 0.002781961, 0.002799779, 
    0.002777988, 0.00270818, 0.00262014, 0.002549058, 0.002503315, 
    0.002479123, 0.002428675, 0.00241998, 0.002388969, 0.002274064, 
    0.002096776, 0.001866611, 0.001720538, 0.001500558, 0.001343742, 
    0.001214551, 0.00115439, 0.001103464, 0.001048102, 0.001094355, 
    0.00112589, 0.001103542, 0.0009533716, 0.001072548, 0.001013485, 
    0.001326544, 0.001930012, 0.000495147, 0.002851676, 0.003573384, 
    0.003761038, 0.003528023, 0.003474683, 0.003312731, 0.003146222, 
    0.002861023, 0.002693765, 0.002515696, 0.002349865, 0.002189826, 
    0.002080312, 0.001998996, 0.001912259, 0.001828843, 0.00173756, 
    0.001669056,
  0.002044931, 0.002145845, 0.002401237, 0.002707384, 0.003585115, 
    0.003557601, 0.003022717, 0.002888916, 0.002681906, 0.002558341, 
    0.003002772, 0.003401089, 0.002784537, 0.002779832, 0.002843633, 
    0.002658319, 0.002530782, 0.002584457, 0.002595473, 0.002589909, 
    0.002602659, 0.002625035, 0.002602641, 0.002576955, 0.002582453, 
    0.002645398, 0.00281232, 0.002986446, 0.003153484, 0.003379058, 
    0.00374667, 0.003584798, 0.002713218, 0.0008081747, 0.001175433, 
    0.001789377, 0.002423873, 0.003494054, 0.003250806, 0.003054507, 
    0.002712043, 0.002850596, 0.003122948, 0.00320185, 0.003195714, 
    0.003134822, 0.003165405, 0.003202217, 0.003263935, 0.00319659, 
    0.003097646, 0.003036102, 0.002979914, 0.002998987, 0.002910281, 
    0.002835432, 0.002818409, 0.002760347, 0.002691999, 0.002509944, 
    0.002309354, 0.002054406, 0.001879629, 0.00170855, 0.001585737, 
    0.001501448, 0.001394556, 0.001413073, 0.00137955, 0.001405539, 
    0.001370269, 0.001321155, 0.001330247, 0.001381331, 0.001336779, 
    0.001886064, 0.002241275, 0.0008514067, 0.003063741, 0.003659056, 
    0.003919648, 0.003622072, 0.003449805, 0.003353663, 0.003035591, 
    0.003187895, 0.002575668, 0.002575906, 0.002440024, 0.002200982, 
    0.002095588, 0.00203711, 0.002010329, 0.001991143, 0.001947241, 
    0.001956937,
  0.002516045, 0.002670065, 0.002822811, 0.002998494, 0.003111059, 
    0.003343723, 0.003130311, 0.002937872, 0.002777973, 0.002452103, 
    0.002589878, 0.00325246, 0.00276947, 0.00274029, 0.002958123, 
    0.002852488, 0.002755435, 0.002854189, 0.002903381, 0.002959887, 
    0.0029593, 0.003027344, 0.003076935, 0.003063791, 0.003068751, 
    0.003142344, 0.003307564, 0.003411515, 0.003556982, 0.003619051, 
    0.003640987, 0.003770828, 0.003769239, 0.003720665, 0.003768062, 
    0.003466165, 0.003382161, 0.00357623, 0.003498221, 0.002773983, 
    0.003104448, 0.003317229, 0.003386607, 0.003392536, 0.003412548, 
    0.003409784, 0.003538243, 0.003525972, 0.003407367, 0.003284583, 
    0.003239062, 0.003245212, 0.003247613, 0.003216811, 0.003173878, 
    0.003108438, 0.003087156, 0.003061136, 0.002949206, 0.002737934, 
    0.002535202, 0.002432251, 0.002320511, 0.002253642, 0.002115503, 
    0.001997231, 0.001874605, 0.001871918, 0.001845834, 0.0018047, 
    0.001754298, 0.001761451, 0.001760544, 0.001736782, 0.001805812, 
    0.002365412, 0.002004479, 0.0020857, 0.002679808, 0.003766509, 
    0.003622705, 0.003378915, 0.003309727, 0.003314132, 0.00320843, 
    0.002942707, 0.002699915, 0.002647894, 0.002549425, 0.002438117, 
    0.002387872, 0.002382753, 0.00238358, 0.002374393, 0.002415147, 
    0.002417451,
  0.002959361, 0.003058767, 0.003114909, 0.003047068, 0.002694222, 
    0.002713122, 0.002823178, 0.002830949, 0.002792373, 0.002598412, 
    0.002776656, 0.003257196, 0.003159685, 0.003092542, 0.003165452, 
    0.003057132, 0.003103146, 0.00315539, 0.003175799, 0.003212053, 
    0.003222194, 0.00325362, 0.003219018, 0.003270261, 0.003368679, 
    0.003469896, 0.003593668, 0.003641892, 0.003717439, 0.003713928, 
    0.003629144, 0.003516482, 0.003479352, 0.00344998, 0.003576327, 
    0.003762882, 0.00366025, 0.003800455, 0.003385814, 0.003061406, 
    0.00326249, 0.003422929, 0.00347268, 0.003459424, 0.003490591, 
    0.003507853, 0.003586546, 0.003471866, 0.003352944, 0.003246879, 
    0.003163576, 0.003079209, 0.00317378, 0.003140099, 0.003231462, 
    0.003214503, 0.003274631, 0.003329055, 0.003218364, 0.003073009, 
    0.002931181, 0.00281992, 0.00271821, 0.002727063, 0.00258681, 
    0.002453629, 0.002325883, 0.002260175, 0.002242691, 0.002272493, 
    0.002263624, 0.002292679, 0.002341188, 0.002439068, 0.002494714, 
    0.002883241, 0.002935106, 0.002585504, 0.002973856, 0.0035518, 
    0.003303638, 0.00302447, 0.003217444, 0.003330071, 0.003050026, 
    0.002740001, 0.002841074, 0.002899598, 0.0029353, 0.002882831, 
    0.002759712, 0.002745202, 0.002746835, 0.002760997, 0.002831854, 
    0.00285344,
  0.00331316, 0.003262045, 0.003260851, 0.003118277, 0.002677773, 
    0.002499371, 0.002585489, 0.002647159, 0.002756149, 0.002743196, 
    0.003014388, 0.003348669, 0.003241269, 0.003264714, 0.003244909, 
    0.003226662, 0.003240285, 0.003167473, 0.003196161, 0.003243241, 
    0.003354615, 0.00331839, 0.003302129, 0.003392823, 0.003369698, 
    0.003399435, 0.003553756, 0.003599802, 0.00366289, 0.003661666, 
    0.00362703, 0.003480276, 0.003366835, 0.003416047, 0.003383653, 
    0.003308425, 0.003291305, 0.003330851, 0.003037836, 0.002902526, 
    0.003083691, 0.003359651, 0.003355121, 0.003287014, 0.003304433, 
    0.003278367, 0.003362607, 0.003364692, 0.003309283, 0.003212452, 
    0.003227536, 0.003164848, 0.003251456, 0.003256287, 0.003302017, 
    0.00331297, 0.003376691, 0.003423342, 0.003342694, 0.003352946, 
    0.003287507, 0.003188277, 0.003080782, 0.003054334, 0.003012611, 
    0.002943022, 0.002881687, 0.002861599, 0.002824893, 0.00287733, 
    0.002889251, 0.002945755, 0.00305155, 0.003088478, 0.002952833, 
    0.002614243, 0.002571485, 0.00274941, 0.003073055, 0.003505833, 
    0.003221165, 0.002950493, 0.002850279, 0.003073135, 0.00304402, 
    0.00280229, 0.00300972, 0.003131151, 0.003085995, 0.003060341, 
    0.003074249, 0.00309852, 0.003066445, 0.00309418, 0.003107216, 0.003144233,
  0.003374895, 0.00334781, 0.003266685, 0.003030475, 0.002886772, 
    0.002746469, 0.002653407, 0.002452373, 0.002535723, 0.002990896, 
    0.003009859, 0.003315082, 0.003360892, 0.003394207, 0.003284868, 
    0.003251635, 0.003186911, 0.003170317, 0.003250092, 0.003229208, 
    0.003307996, 0.003336256, 0.003416954, 0.003497729, 0.003397625, 
    0.003404237, 0.003502561, 0.003276825, 0.003019873, 0.003411675, 
    0.003398484, 0.003400596, 0.003298234, 0.003283802, 0.003260087, 
    0.003322506, 0.003313906, 0.002941402, 0.002730955, 0.003026325, 
    0.003070705, 0.003281195, 0.003211481, 0.003188532, 0.003213024, 
    0.0031943, 0.003383717, 0.00350407, 0.003521299, 0.003473965, 
    0.003534636, 0.003587309, 0.003705502, 0.003788535, 0.00381284, 
    0.003808897, 0.003828162, 0.003774406, 0.003733635, 0.003743459, 
    0.003752008, 0.003711892, 0.003665194, 0.003575437, 0.003501829, 
    0.003498476, 0.003483152, 0.003411943, 0.003340896, 0.003420988, 
    0.003390757, 0.003395652, 0.003266048, 0.003167503, 0.003144709, 
    0.002948157, 0.002734039, 0.003204869, 0.003745683, 0.003539657, 
    0.002963798, 0.002618823, 0.002413256, 0.002150854, 0.003184954, 
    0.003006585, 0.003148111, 0.003280289, 0.003275475, 0.003274202, 
    0.00329911, 0.00330515, 0.003248993, 0.003351036, 0.003343312, 0.003290288,
  0.003217505, 0.003162449, 0.003095753, 0.002826437, 0.002860116, 
    0.002606312, 0.00230352, 0.002076815, 0.002673591, 0.003279526, 
    0.002704762, 0.003353901, 0.003348971, 0.003382079, 0.003321568, 
    0.003251743, 0.003184717, 0.003190169, 0.00322555, 0.003302624, 
    0.003303593, 0.00335657, 0.003414823, 0.003374213, 0.003356079, 
    0.003316212, 0.003303479, 0.002931928, 0.002846576, 0.003315829, 
    0.003014136, 0.002918988, 0.002654633, 0.002883196, 0.002984809, 
    0.003017457, 0.002894146, 0.002878621, 0.002911869, 0.003002547, 
    0.003094085, 0.003185416, 0.003215455, 0.003283644, 0.0033336, 
    0.003353914, 0.003408065, 0.003395589, 0.003397625, 0.003378376, 
    0.003364597, 0.003407924, 0.003477972, 0.003627826, 0.003698079, 
    0.003758796, 0.003784815, 0.003749417, 0.003699191, 0.003673077, 
    0.003677431, 0.003627254, 0.003597831, 0.003616747, 0.003571765, 
    0.003557587, 0.003580444, 0.003582478, 0.003525097, 0.003541119, 
    0.003487363, 0.003467577, 0.00332381, 0.003214311, 0.002960032, 
    0.002945803, 0.003661025, 0.004131177, 0.004045647, 0.002997635, 
    0.00239841, 0.001905868, 0.001599945, 0.001865593, 0.002619551, 
    0.003067717, 0.003085246, 0.00324014, 0.003297886, 0.003228234, 
    0.003219811, 0.003269974, 0.003237294, 0.003231494, 0.003234226, 
    0.003264794,
  0.003176292, 0.003348144, 0.003166595, 0.002551762, 0.002031897, 
    0.002117839, 0.002108509, 0.002304059, 0.002982805, 0.003482944, 
    0.0028666, 0.003179676, 0.003149275, 0.003304608, 0.003443129, 
    0.003491925, 0.003349766, 0.003186243, 0.003154518, 0.003302593, 
    0.003266923, 0.003242176, 0.003304513, 0.003337907, 0.003377231, 
    0.003316611, 0.00306306, 0.00264379, 0.003058417, 0.003107328, 
    0.002784872, 0.002476564, 0.002508894, 0.002971778, 0.002756787, 
    0.002756787, 0.002743371, 0.002833318, 0.002897803, 0.002987305, 
    0.003051661, 0.003049485, 0.003098186, 0.003210433, 0.003314653, 
    0.003395749, 0.003453018, 0.003434548, 0.003440285, 0.003460201, 
    0.00343674, 0.003408687, 0.003355248, 0.003342183, 0.003371317, 
    0.003455799, 0.003491433, 0.003566584, 0.00358448, 0.003571987, 
    0.003544919, 0.00351386, 0.003498888, 0.00348549, 0.003468037, 
    0.003450077, 0.003419876, 0.00346899, 0.003495932, 0.003515022, 
    0.003436407, 0.00338974, 0.003213245, 0.003117561, 0.002885867, 
    0.003028439, 0.003312299, 0.003502033, 0.003390707, 0.002256233, 
    0.002160977, 0.001498873, 0.001979746, 0.002906339, 0.00278333, 
    0.002740478, 0.002723439, 0.002850024, 0.002894402, 0.002936522, 
    0.00305899, 0.003047386, 0.003096072, 0.003250059, 0.003290892, 
    0.003292495,
  0.002736504, 0.002947744, 0.001568221, 0.00205326, 0.001736242, 
    0.002043881, 0.002192417, 0.002047395, 0.002441468, 0.003146536, 
    0.003349016, 0.002862611, 0.003006249, 0.003053876, 0.003301319, 
    0.003553582, 0.003681755, 0.003620116, 0.003442001, 0.003340865, 
    0.003306691, 0.003295025, 0.003251061, 0.003266383, 0.003269879, 
    0.003339244, 0.002872307, 0.002440737, 0.003005646, 0.002942117, 
    0.002900632, 0.002839899, 0.00304769, 0.003134044, 0.002948284, 
    0.002980281, 0.003021494, 0.003105562, 0.003150068, 0.003217684, 
    0.003227506, 0.003189279, 0.003155567, 0.003128992, 0.003162323, 
    0.003271947, 0.003314782, 0.003344648, 0.003399055, 0.003494231, 
    0.00354851, 0.003565202, 0.003572639, 0.003530838, 0.003418908, 
    0.003378328, 0.003316863, 0.003310665, 0.003273567, 0.003255446, 
    0.00317858, 0.003200356, 0.003238471, 0.003206236, 0.003245942, 
    0.00331324, 0.00338785, 0.003490368, 0.003548622, 0.003613153, 
    0.003465589, 0.003442414, 0.003398545, 0.003373925, 0.003506962, 
    0.003571794, 0.003232191, 0.003490192, 0.003283229, 0.001706964, 
    0.002259665, 0.00270419, 0.002897073, 0.002864823, 0.002691858, 
    0.002695132, 0.002721135, 0.002729114, 0.002760775, 0.002848323, 
    0.002938397, 0.003023101, 0.003282197, 0.003223689, 0.002093076, 
    0.002502487,
  0.001336334, 0.0016194, 0.001442112, 0.001733254, 0.001912783, 0.001909095, 
    0.001680086, 0.001868167, 0.002395771, 0.002743275, 0.003095753, 
    0.002889615, 0.002874246, 0.002768038, 0.003123805, 0.003329692, 
    0.003468769, 0.003590902, 0.003601456, 0.003536813, 0.003293594, 
    0.003073801, 0.003153928, 0.003123252, 0.003047546, 0.003009224, 
    0.002800656, 0.0027757, 0.002669254, 0.002649896, 0.002841633, 
    0.002976133, 0.002949048, 0.002776574, 0.003033971, 0.003092464, 
    0.00306681, 0.003126239, 0.003098885, 0.003064394, 0.003033526, 
    0.003057543, 0.003039153, 0.003047148, 0.00306139, 0.003124952, 
    0.003160588, 0.003187133, 0.003229825, 0.003263155, 0.003312239, 
    0.003399007, 0.003433466, 0.003482342, 0.003471294, 0.003432799, 
    0.00329593, 0.003158236, 0.003005583, 0.002933279, 0.002866777, 
    0.002817711, 0.002854204, 0.002869925, 0.00286161, 0.002951209, 
    0.003066842, 0.003283931, 0.003443718, 0.003552597, 0.003656132, 
    0.003628857, 0.003401009, 0.003265364, 0.003116798, 0.003102094, 
    0.003112092, 0.003411386, 0.003135282, 0.002951064, 0.003059784, 
    0.002879474, 0.002983112, 0.002909616, 0.002832921, 0.002783012, 
    0.002777195, 0.002766624, 0.002790799, 0.002752557, 0.002859639, 
    0.003157841, 0.003047434, 0.002327424, 0.001439442, 0.001284565,
  0.001904517, 0.001646215, 0.001498189, 0.00157302, 0.001466162, 0.00143159, 
    0.001327482, 0.00146411, 0.001970449, 0.002892556, 0.002770309, 
    0.002086431, 0.002049223, 0.002108444, 0.002738569, 0.002935313, 
    0.003061451, 0.003261804, 0.003511399, 0.003608277, 0.002961077, 
    0.002847319, 0.003260886, 0.003088731, 0.002847483, 0.002655935, 
    0.00232291, 0.002229466, 0.002017686, 0.001983911, 0.002601909, 
    0.002784649, 0.002776735, 0.002656791, 0.002829583, 0.00297424, 
    0.00311726, 0.003167184, 0.003158538, 0.003190583, 0.003167724, 
    0.003116146, 0.003030252, 0.003022654, 0.003006984, 0.002951305, 
    0.002910519, 0.002916718, 0.002930084, 0.002951115, 0.003010577, 
    0.003081199, 0.003119186, 0.003192252, 0.003230972, 0.003203301, 
    0.003098248, 0.003016885, 0.002917988, 0.002768882, 0.002632998, 
    0.002542146, 0.00252687, 0.002515156, 0.00247941, 0.002569262, 
    0.002571391, 0.002905671, 0.003259532, 0.003264571, 0.003343141, 
    0.003130168, 0.003046287, 0.002596997, 0.003075331, 0.00323493, 
    0.00318669, 0.002991628, 0.002952781, 0.002859766, 0.002853106, 
    0.002776002, 0.002725283, 0.002566717, 0.002592323, 0.002491155, 
    0.002536057, 0.002567909, 0.002569053, 0.002512024, 0.002657667, 
    0.002689868, 0.002031388, 0.001804366, 0.001834566, 0.001700797,
  0.0007848279, 0.0007950794, 0.0007628612, 0.0006462899, 0.0005062581, 
    0.0007338375, 0.0007117437, 0.0005971598, 0.0007066415, 0.001800931, 
    0.002862834, 0.002425, 0.001455593, 0.001229621, 0.001688717, 
    0.002651117, 0.002722801, 0.002604133, 0.002964621, 0.003142213, 
    0.002710007, 0.002912583, 0.003126365, 0.002923756, 0.002793374, 
    0.00250929, 0.002169067, 0.001874811, 0.001324588, 0.001793001, 
    0.002317252, 0.002498483, 0.002490217, 0.00249985, 0.002630856, 
    0.002617091, 0.002741273, 0.002839565, 0.002877012, 0.002858432, 
    0.002840362, 0.002861818, 0.002848294, 0.002815679, 0.002732022, 
    0.002735518, 0.002710944, 0.002702475, 0.002714744, 0.002747551, 
    0.002715046, 0.002712598, 0.002781771, 0.002822301, 0.002830932, 
    0.0028467, 0.002814705, 0.002663468, 0.002461002, 0.00223344, 
    0.002070553, 0.001992765, 0.001964661, 0.001965713, 0.001983452, 
    0.002014684, 0.002001476, 0.002200125, 0.002276976, 0.002195261, 
    0.002121748, 0.001814524, 0.001829622, 0.002575777, 0.002967281, 
    0.003018716, 0.00303575, 0.002933884, 0.002935155, 0.002794805, 
    0.002648115, 0.002526426, 0.002358386, 0.002216401, 0.002212904, 
    0.002094775, 0.002177347, 0.002161883, 0.002205386, 0.002192638, 
    0.002374616, 0.002449368, 0.001519361, 0.001196877, 0.0008007223, 
    0.0006467667,
  0.000416311, 0.0004365288, 0.0003874623, 0.0005865104, 0.000177193, 
    0.0004564286, 0.000593297, 0.0006363078, 0.0005228841, 0.001206572, 
    0.002394102, 0.001575247, 0.001246152, 0.0008402194, 0.0007738597, 
    0.001876036, 0.002510133, 0.002147038, 0.002268489, 0.002356306, 
    0.002267295, 0.002178731, 0.002148118, 0.002177014, 0.002425319, 
    0.002033295, 0.001757811, 0.001791124, 0.0009487462, 0.0009143651, 
    0.001695362, 0.001942887, 0.00197261, 0.001983131, 0.002004701, 
    0.002041496, 0.002157336, 0.00228497, 0.002385567, 0.002469124, 
    0.002542878, 0.002535183, 0.002493125, 0.002447874, 0.002309702, 
    0.002275909, 0.002246029, 0.002239496, 0.002276004, 0.002313865, 
    0.002325485, 0.002375537, 0.002459492, 0.002492887, 0.002538186, 
    0.002564874, 0.002536723, 0.002398695, 0.002203351, 0.001974072, 
    0.001756459, 0.001546429, 0.001427395, 0.001468833, 0.001534573, 
    0.001599818, 0.001626458, 0.001543313, 0.0009736679, 0.001020112, 
    0.001206157, 0.001325098, 0.001524176, 0.002131986, 0.002420248, 
    0.002663406, 0.002938094, 0.002973572, 0.002839405, 0.002714904, 
    0.002607408, 0.002377826, 0.00218992, 0.001970035, 0.001792857, 
    0.001706264, 0.001720013, 0.001701052, 0.001792875, 0.00182468, 
    0.001986042, 0.002087846, 0.0009180391, 0.0005478226, 0.0001676404, 
    9.26021e-005,
  0.0007143982, 0.0004766786, 0.0002790135, 0.0001753969, 0.0002688251, 
    0.0004674438, 0.000387033, 0.0005849365, 0.0005100886, 0.0008605332, 
    0.001726833, 0.0008282983, 0.001120568, 0.0012956, 0.0008546833, 
    0.0012146, 0.002255074, 0.001904438, 0.001069657, 0.001067655, 
    0.001171764, 0.001410802, 0.001434564, 0.001338163, 0.001804891, 
    0.001600852, 0.001309013, 0.001505326, 0.0009708391, 0.0007531322, 
    0.0008715629, 0.001105339, 0.001598373, 0.001593413, 0.001553724, 
    0.001633483, 0.001691498, 0.00168487, 0.001730853, 0.001795513, 
    0.001879849, 0.001933017, 0.001933414, 0.001953505, 0.001893248, 
    0.001819497, 0.00172432, 0.001630876, 0.001619687, 0.001713623, 
    0.001831942, 0.001944063, 0.002042148, 0.002137452, 0.00220936, 
    0.00224722, 0.002256249, 0.002220518, 0.002110353, 0.001901101, 
    0.001697825, 0.001525878, 0.001388771, 0.001322458, 0.001289699, 
    0.001311983, 0.001314606, 0.0006508334, 0.0005830596, 0.001060166, 
    0.00126128, 0.001612216, 0.001462935, 0.001694883, 0.002010566, 
    0.002199235, 0.00239326, 0.002559341, 0.002681682, 0.002656252, 
    0.002581388, 0.00244622, 0.002330491, 0.002136419, 0.00201357, 
    0.001871726, 0.001734447, 0.001683949, 0.00164566, 0.001648283, 
    0.001789283, 0.001826523, 0.0009732572, 0.0007441523, 0.0008521883, 
    0.0006917482,
  0.0006482606, 0.0007628924, 0.0005715536, 0.0003847764, 0.0007711579, 
    0.0009276704, 0.0004621986, 0.0006472273, 0.001108345, 0.0008418567, 
    0.0006584332, 0.0005904357, 0.0009342041, 0.001097378, 0.0009947792, 
    0.0009483825, 0.0009451224, 0.0008286792, 0.0007217096, 0.0005966828, 
    0.0008103698, 0.0009271952, 0.001012247, 0.0007856053, 0.001018032, 
    0.001359162, 0.001012819, 0.001118788, 0.0008395198, 0.0007915341, 
    0.0007450108, 0.0007200404, 0.001062012, 0.001366121, 0.001376229, 
    0.001425616, 0.001457468, 0.001508712, 0.001558875, 0.001523303, 
    0.001495106, 0.001554536, 0.001546429, 0.001517453, 0.001441175, 
    0.00135134, 0.001282961, 0.001162083, 0.001070037, 0.001069576, 
    0.001158554, 0.00130863, 0.001496584, 0.001686063, 0.00180122, 
    0.001885683, 0.001929298, 0.001901212, 0.001832612, 0.001731823, 
    0.001624345, 0.001482867, 0.001323698, 0.001242699, 0.001225596, 
    0.001126081, 0.0004230966, 0.0003988105, 0.0005768137, 0.0008985037, 
    0.0009954125, 0.001513703, 0.001502751, 0.001637712, 0.001311682, 
    0.001797403, 0.001987678, 0.002066945, 0.002159228, 0.002228464, 
    0.002267517, 0.002261907, 0.002178524, 0.00205957, 0.001984133, 
    0.001827143, 0.001704183, 0.001673475, 0.001589201, 0.001506121, 
    0.001508791, 0.001605001, 0.001659757, 0.0008906517, 0.0005822189, 
    0.000393661,
  0.0007739714, 0.0004282161, 0.0003294633, 0.0007559778, 0.001150242, 
    0.001497043, 0.0007576137, 0.0008169804, 0.001546714, 0.001069545, 
    0.000663647, 0.000654221, 0.0007846204, 0.000789071, 0.0009094246, 
    0.0009208526, 0.0007181808, 0.0009420402, 0.001065032, 0.0005788172, 
    0.0001071456, 0.000552734, 0.0004791422, 0.000373634, 0.0004241471, 
    0.0004972938, 0.000516399, 0.0008083822, 0.0007699173, 0.0007510348, 
    0.0008858524, 0.0009225531, 0.0009222829, 0.0007292423, 0.0008092867, 
    0.001178406, 0.001293896, 0.001355329, 0.001388531, 0.001419893, 
    0.001387578, 0.001351099, 0.001300301, 0.001262281, 0.001217507, 
    0.001130229, 0.001084675, 0.001034004, 0.0009673256, 0.0009019356, 
    0.0008767741, 0.0009007128, 0.0009915177, 0.001181808, 0.00131572, 
    0.001415633, 0.001475411, 0.001451889, 0.00145405, 0.0014386, 
    0.001411865, 0.001335523, 0.001193776, 0.001145788, 0.001158902, 
    0.0008706087, 0.000462899, 0.0003809142, 0.0004671426, 0.0005309274, 
    0.0006071888, 0.0007522106, 0.0006575421, 0.0007086433, 0.000960683, 
    0.001495154, 0.001651969, 0.001666815, 0.001701482, 0.001727548, 
    0.001761085, 0.001803318, 0.001789616, 0.00170617, 0.001625394, 
    0.001560147, 0.001457324, 0.001394573, 0.001472726, 0.001518423, 
    0.001458342, 0.001480657, 0.00149671, 0.001464889, 0.0009971145, 
    0.0009242222,
  0.0007947446, 0.0007274151, 0.0008920822, 0.001476652, 0.001635978, 
    0.00164739, 0.001413357, 0.001332265, 0.001491608, 0.001493483, 
    0.000854508, 0.0006485153, 0.0008024857, 0.0008097813, 0.0008422856, 
    0.0009086775, 0.0007660869, 0.0009276078, 0.0009507977, 0.0004981204, 
    0.0003539088, 0.0004444762, 0.0004303937, 0.0003567699, 0.000337935, 
    0.0002906327, 0.0002719087, 0.0004193626, 0.0007055287, 0.0006287261, 
    0.0006103201, 0.0006067597, 0.0008696559, 0.0006993306, 0.0008385978, 
    0.001014279, 0.0008059032, 0.000779391, 0.00114053, 0.001227599, 
    0.001244353, 0.001235896, 0.001221909, 0.001177261, 0.001113477, 
    0.001053205, 0.0009944737, 0.0009408626, 0.0009306418, 0.000905036, 
    0.0008688434, 0.0008340497, 0.0008118451, 0.0008774903, 0.000962859, 
    0.001056382, 0.001163878, 0.001185304, 0.001199387, 0.00117831, 
    0.001162732, 0.001185128, 0.00114091, 0.001045941, 0.0008386131, 
    0.0006320323, 0.0005075939, 0.0005362674, 0.0005177979, 0.0003096906, 
    0.0005232021, 0.0006930516, 0.0007401635, 0.0006955159, 0.0007340442, 
    0.0008879662, 0.001285234, 0.001406828, 0.001515816, 0.001578361, 
    0.001592761, 0.001484615, 0.001415903, 0.001404952, 0.001343409, 
    0.001296883, 0.001175163, 0.001045892, 0.001162241, 0.001309473, 
    0.001355439, 0.001354438, 0.001312477, 0.001426076, 0.001462267, 
    0.001084041,
  0.000972732, 0.001266002, 0.001378789, 0.001492085, 0.001581571, 
    0.00142703, 0.001086856, 0.0008555267, 0.0007467752, 0.0007377316, 
    0.0007437712, 0.0007968107, 0.0008289337, 0.0007832854, 0.0009685513, 
    0.000879463, 0.0009117131, 0.000911888, 0.0009331228, 0.0005321348, 
    0.0003544015, 0.0003371242, 0.0001567209, 0.0002297087, 0.0003235186, 
    0.0003444676, 0.0003351534, 0.0003013297, 0.0003151102, 0.0003472808, 
    0.0003169381, 0.0003198945, 0.0004011476, 0.0003149673, 0.0003616337, 
    0.0008342108, 0.0009206287, 0.0006848814, 0.0009393692, 0.001031922, 
    0.001067924, 0.001089143, 0.001076649, 0.001032796, 0.0009861621, 
    0.0009315005, 0.0008765212, 0.0008409331, 0.0008164234, 0.0008152951, 
    0.0008268664, 0.0008056154, 0.0007983991, 0.0008393596, 0.000866889, 
    0.0008795732, 0.0009318809, 0.0009796768, 0.001029061, 0.001063043, 
    0.001047672, 0.001037724, 0.0009974623, 0.0008140882, 0.000765038, 
    0.0007855734, 0.0007812022, 0.0006601014, 0.0005589325, 0.0006513281, 
    0.0006270574, 0.0006550951, 0.0008146132, 0.0007050997, 0.0005501115, 
    0.0006613892, 0.0009126035, 0.001366932, 0.001439283, 0.001512795, 
    0.001524716, 0.001401151, 0.001158505, 0.000987988, 0.001021668, 
    0.000997588, 0.0008468768, 0.0006521996, 0.0005810549, 0.0008033887, 
    0.001047689, 0.001148906, 0.001164116, 0.001262965, 0.00122946, 
    0.001031701,
  0.0009194701, 0.001227394, 0.001321951, 0.001297076, 0.001403982, 
    0.001169858, 0.0009120784, 0.0007169091, 0.0005755743, 0.0005186561, 
    0.0005911035, 0.0006692254, 0.0007249035, 0.0007623844, 0.0007791528, 
    0.0008614382, 0.0007905962, 0.001222563, 0.001185687, 0.0006284558, 
    0.0004868193, 0.0004523916, 0.0004037224, 0.0003504596, 0.0002570475, 
    0.0001982375, 0.0002142751, 0.0002000336, 0.000200574, 0.000210365, 
    0.0002008124, 0.0002224608, 0.0002186302, 0.0001954084, 0.0001817072, 
    0.0002226675, 0.0006865829, 0.0008057291, 0.0006422522, 0.0008889523, 
    0.0009239363, 0.0007916936, 0.0006913194, 0.0006555088, 0.0006360696, 
    0.000636118, 0.0006468464, 0.000661104, 0.0006670002, 0.0006827828, 
    0.0007298947, 0.0007511298, 0.0007762583, 0.0008470686, 0.0009055454, 
    0.0009157811, 0.0009147795, 0.0009344728, 0.0009881803, 0.001009749, 
    0.001011291, 0.001012022, 0.0009817593, 0.0007912167, 0.000802692, 
    0.0006801765, 0.0004884885, 0.000398652, 0.0004966418, 0.0007177512, 
    0.0009045447, 0.0007569315, 0.0007786436, 0.0008467038, 0.0008051717, 
    0.0007797242, 0.0007506054, 0.0008215744, 0.001205509, 0.001260996, 
    0.001126289, 0.0009056088, 0.0009218846, 0.0008482928, 0.0007950454, 
    0.0007407656, 0.0005554347, 0.0004096017, 0.000421348, 0.000557771, 
    0.0007950757, 0.0009680092, 0.001074678, 0.001163593, 0.001076078, 
    0.00088207,
  0.0009084553, 0.0009053557, 0.001064794, 0.001052873, 0.0009959224, 
    0.00094657, 0.0008297602, 0.0007191182, 0.0006354493, 0.0005191169, 
    0.0005128067, 0.0005250454, 0.0005075934, 0.0005573593, 0.0006578136, 
    0.0006433174, 0.0005545779, 0.0006084923, 0.0006223206, 0.0006151998, 
    0.0006690505, 0.0005459472, 0.000318607, 0.0002398337, 0.0002250358, 
    0.0001804992, 0.0001756035, 0.0001826448, 0.0001793547, 0.0001764301, 
    0.000188351, 0.00017465, 0.000148869, 0.0001453087, 0.0001598203, 
    0.0001162056, 0.000119925, 0.0005487285, 0.0006755355, 0.0005789283, 
    0.0005711399, 0.0005620322, 0.0005508743, 0.0005170032, 0.0004987086, 
    0.0005165106, 0.0005337086, 0.0005564219, 0.0005789921, 0.0006030574, 
    0.0006525209, 0.0007244758, 0.0007965416, 0.0008454649, 0.0009123012, 
    0.0009840489, 0.0009977017, 0.0009844615, 0.001025215, 0.001047214, 
    0.00105745, 0.001044733, 0.0009693136, 0.0008187783, 0.0008172514, 
    0.0005919142, 0.0004971509, 0.0005342963, 0.0006840071, 0.0007354739, 
    0.0005675638, 0.0005994482, 0.0006840074, 0.0008591812, 0.0007464095, 
    0.0007222499, 0.0006667301, 0.0006744707, 0.0007594589, 0.0008933387, 
    0.0009006825, 0.0008199543, 0.0006886646, 0.0006041534, 0.0006056, 
    0.0006524562, 0.0005413047, 0.0003276342, 0.0002264171, 0.0003521116, 
    0.0005029347, 0.0006719898, 0.0008345591, 0.0009512734, 0.001046975, 
    0.0009594597,
  0.0007172115, 0.0007326452, 0.0008561299, 0.0008652217, 0.0008538407, 
    0.0008459254, 0.0007817745, 0.0006382787, 0.0004992168, 0.0004290427, 
    0.0004088088, 0.0004414404, 0.0004712428, 0.0004814313, 0.000430648, 
    0.0003927393, 0.0003662272, 0.0003465498, 0.0002853079, 0.0003036503, 
    0.0004007819, 0.0004147373, 0.0003310048, 0.0002445383, 0.0002027834, 
    0.00017101, 0.0001716299, 0.0001820567, 0.0001745227, 0.0001567208, 
    0.0001625383, 0.0001346752, 0.0001084332, 0.0001101657, 0.0001137261, 
    8.937554e-005, 7.956856e-005, 0.0001500293, 0.0007328354, 0.0006311579, 
    0.000540813, 0.000533581, 0.0005598709, 0.0005527022, 0.00055577, 
    0.0005547847, 0.0005308315, 0.0005205795, 0.0005534494, 0.0005960313, 
    0.000639376, 0.0007353951, 0.000840236, 0.0008996339, 0.0009482875, 
    0.001022021, 0.00106899, 0.001064063, 0.001069832, 0.001071929, 
    0.001071707, 0.001018667, 0.0008556219, 0.0006964048, 0.0006093027, 
    0.0006095574, 0.0006464963, 0.0006978675, 0.0006202224, 0.0006520435, 
    0.0006000204, 0.0005966349, 0.0006011489, 0.0006140871, 0.0006672385, 
    0.0007166865, 0.0007015072, 0.0006063305, 0.0005401932, 0.0006386761, 
    0.0008689405, 0.0009114271, 0.000716019, 0.0006498818, 0.0006300139, 
    0.0005605873, 0.000373174, 0.0001021381, -6.957073e-005, -2.729194e-005, 
    0.000189669, 0.0004469384, 0.0006167241, 0.0006988994, 0.0007721256, 
    0.0008085719,
  0.0006020553, 0.0007322789, 0.0007575201, 0.0007032875, 0.0006466708, 
    0.00065829, 0.0006441597, 0.0005648298, 0.0004376573, 0.0003532096, 
    0.0002882165, 0.0002573493, 0.0002687458, 0.0003086571, 0.0003033644, 
    0.0002434893, 0.0002042456, 0.0002311392, 0.0002535982, 0.0002314729, 
    0.0002270861, 0.0002521201, 0.0002550605, 0.0002389752, 0.0002217297, 
    0.0001983171, 0.0001797999, 0.0001640641, 0.0001437987, 0.0001314326, 
    0.0001237397, 0.0001018846, 9.985012e-005, 9.778378e-005, 7.861496e-005, 
    4.695295e-005, 6.272031e-005, 0.0001843139, 0.0008502963, 0.0008711974, 
    0.000641918, 0.0005956013, 0.0004584634, 0.0005353454, 0.0005786421, 
    0.0005840305, 0.0005544033, 0.0005222326, 0.0005524957, 0.0006189351, 
    0.0006950384, 0.0008094478, 0.0009305484, 0.001008258, 0.001040651, 
    0.001067973, 0.001066273, 0.001076508, 0.001106422, 0.001103036, 
    0.001022228, 0.000995907, 0.0007929327, 0.0006355769, 0.0005927725, 
    0.0006433331, 0.0006835305, 0.0007076585, 0.0006964528, 0.0006663008, 
    0.0006148659, 0.0005692167, 0.0006107015, 0.0007458053, 0.0009384953, 
    0.001587359, 0.0008544765, 0.0006091915, 0.0004776006, 0.0005520983, 
    0.0007592999, 0.001026774, 0.0007530216, 0.0006181723, 0.0005380476, 
    0.0005254115, 0.0004068383, 0.000194964, 9.219162e-006, -3.307685e-005, 
    0.0001026634, 0.000345245, 0.0005012504, 0.00054566, 0.0004930031, 
    0.0005268743,
  0.0005224873, 0.0005757818, 0.0005804072, 0.0005319756, 0.000535409, 
    0.000582902, 0.000528622, 0.000390721, 0.0002896471, 0.0002851172, 
    0.0003023311, 0.0002882007, 0.0002715276, 0.0002715115, 0.0002665365, 
    0.0002282307, 0.0002002243, 0.0001957897, 0.0002099993, 0.000206741, 
    0.0002114618, 0.0002226834, 0.0002116684, 0.0001983965, 0.0001987779, 
    0.0001996681, 0.0001872385, 0.000142225, 0.0001166984, 0.0001096412, 
    9.14101e-005, 7.449827e-005, 7.836064e-005, 7.818578e-005, 5.701419e-005, 
    3.852877e-005, 6.643965e-005, 0.0001817707, 0.0008169495, 0.001068958, 
    0.001036994, 0.0008415862, 0.0003322605, 0.0003296062, 0.0005372686, 
    0.0005910876, 0.0006589417, 0.0007533233, 0.0008100991, 0.0008582596, 
    0.0009338225, 0.001011674, 0.001047485, 0.001100604, 0.001209116, 
    0.001072487, 0.00106462, 0.001015585, 0.001020337, 0.001030526, 
    0.001024008, 0.0008125305, 0.0006968979, 0.0006567641, 0.0007037008, 
    0.0007768953, 0.0007590456, 0.0006320956, 0.0005126004, 0.0004905863, 
    0.0005605225, 0.0006657923, 0.001176469, 0.001450587, 0.001617003, 
    0.00159181, 0.0007546429, 0.000556517, 0.0005278591, 0.0006479108, 
    0.001360862, 0.001188771, 0.0008831499, 0.0007056557, 0.0005710446, 
    0.0006164238, 0.0005727776, 0.0004384364, 0.0003261734, 0.0003157463, 
    0.0003637155, 0.0004381975, 0.0005096914, 0.0005435147, 0.0005459627, 
    0.0004976755,
  0.0004227646, 0.0004621996, 0.0004206819, 0.0003361863, 0.0003735072, 
    0.0006019277, 0.0004711791, 0.000350571, 0.0002357964, 0.000192865, 
    0.0002063437, 0.000236321, 0.0002455715, 0.0002404694, 0.0002327923, 
    0.0002385143, 0.0002363844, 0.0002137823, 0.0001839164, 0.0001621885, 
    0.0001702472, 0.0001979831, 0.0002006375, 0.0001879855, 0.000170581, 
    0.0001545275, 0.0001453881, 0.0001311307, 0.0001201793, 0.0001121207, 
    9.490689e-005, 6.982521e-005, 5.655322e-005, 5.48684e-005, 5.067224e-005, 
    4.20097e-005, 4.173948e-005, 6.140108e-005, 8.320843e-005, 9.93891e-005, 
    0.0001089417, 0.0001251224, 0.0001344208, 0.0001522386, 0.000208696, 
    0.0003278101, 0.0004924937, 0.001255274, 0.001375389, 0.001480071, 
    0.001573515, 0.001616637, 0.0009991012, 0.0009210749, 0.0008910341, 
    0.0008741064, 0.0008386616, 0.0007790568, 0.0007101222, 0.0006690823, 
    0.0006547295, 0.0006465915, 0.0006364031, 0.0006218119, 0.0005863193, 
    0.000564512, 0.0005269531, 0.0004629298, 0.0004158978, 0.0004171535, 
    0.0004846577, 0.0007919155, 0.0009341084, 0.001039601, 0.001017603, 
    0.0009270514, 0.0005889419, 0.0005181315, 0.0007149383, 0.0008643472, 
    0.001239459, 0.00130229, 0.0009432001, 0.0006375634, 0.0005826, 
    0.0005712828, 0.0005570895, 0.0005517965, 0.0005424186, 0.0005668332, 
    0.0005445648, 0.0004450968, 0.000283767, 0.0002134964, 0.0003411458, 
    0.0004093978,
  0.0002432829, 0.0003104853, 0.0002579698, 0.0003649876, 0.0003463749, 
    0.0003565475, 0.0006961189, 0.0003532413, 0.0003058754, 0.0002571426, 
    0.0002426152, 0.0002551719, 0.0002590025, 0.0002297089, 0.0001821045, 
    0.0001455153, 0.0001414462, 0.0001495205, 0.0001682921, 0.000183821, 
    0.0001850451, 0.0001800064, 0.0001633808, 0.0001508241, 0.000142686, 
    0.0001291597, 0.0001169844, 0.0001032515, 9.007493e-005, 7.489556e-005, 
    6.715492e-005, 5.962086e-005, 5.507507e-005, 5.39465e-005, 5.491608e-005, 
    5.712541e-005, 6.443693e-005, 5.941425e-005, 5.900099e-005, 
    5.847646e-005, 6.119446e-005, 8.347865e-005, 0.000100915, 0.0001191143, 
    0.0001317823, 0.0001381719, 0.0001521115, 0.0002012574, 0.0002939069, 
    0.0004192516, 0.0005655134, 0.001170381, 0.0007175289, 0.0006649497, 
    0.0005936944, 0.0005405906, 0.0005129341, 0.0004993284, 0.0004853889, 
    0.0004654729, 0.0004647894, 0.0004719897, 0.0004881545, 0.0004675393, 
    0.000420253, 0.0003655916, 0.0003178919, 0.0002902194, 0.0002704147, 
    0.0002636118, 0.0002625787, 0.0002733711, 0.0002972765, 0.0003318155, 
    0.0004304413, 0.0004270079, 0.0003920082, 0.0002764387, 0.000263135, 
    0.0003177488, 0.000554578, 0.0007499857, 0.0004110499, 0.0003114864, 
    0.0002668226, 0.0002757711, 0.0003425919, 0.0003552756, 0.0004862789, 
    0.000635227, 0.0007679628, 0.0009168785, 0.0006573361, 0.0004016883, 
    0.0002209351, 0.0001748567,
  0.0003111209, 0.0002533442, 0.0002193772, 0.0001622841, 5.375571e-005, 
    0.0002930487, 0.0002741341, 0.0002566181, 0.0002666479, 0.0003065909, 
    0.0003824396, 0.0007659119, 0.0009064202, 0.0008818947, 0.0003570243, 
    0.0002520248, 0.000180213, 0.0001542573, 0.0001606945, 0.0001698975, 
    0.0001677359, 0.0001561646, 0.0001390779, 0.0001265689, 0.0001165235, 
    0.0001133605, 0.000101821, 8.56244e-005, 7.542007e-005, 6.920533e-005, 
    6.891922e-005, 6.775891e-005, 6.324484e-005, 5.612408e-005, 
    6.051097e-005, 6.294285e-005, 6.829931e-005, 8.30018e-005, 8.255675e-005, 
    8.484558e-005, 8.646683e-005, 9.126699e-005, 0.0001047297, 0.0001163168, 
    0.0001300656, 0.0001243754, 0.0001242641, 0.0001346274, 0.0001678947, 
    0.0002439026, 0.0003533526, 0.0004737541, 0.0005406862, 0.0004015768, 
    0.0003638749, 0.0003298605, 0.0003161276, 0.0003233755, 0.0003320539, 
    0.0003236456, 0.0003121698, 0.0002926513, 0.0002786322, 0.0002550924, 
    0.0002285802, 0.0002091253, 0.0002027515, 0.0002078219, 0.0002208554, 
    0.0002902353, 0.0002275947, 0.0002194408, 0.000210222, 0.000252279, 
    0.0002079968, 0.0002495769, 0.0002033714, 0.0002051834, 0.000228612, 
    0.0003318791, 0.0003839657, 0.0003989541, 0.0002345248, 0.0001620138, 
    0.000114187, 9.471609e-005, 0.0001136784, 0.0001804356, 0.0002947811, 
    0.0004440152, 0.0008412363, 0.001064889, 0.001357619, 0.001107264, 
    0.0007289732, 0.0004865015,
  0.0006943229, 0.0005198962, 0.0003628735, 0.0002800948, 0.0001883353, 
    0.0002218091, 0.0003615539, 0.0005246643, 0.0006664118, 0.0007853666, 
    0.0008946103, 0.001048247, 0.001169141, 0.001053318, 0.0007240776, 
    0.0003891313, 0.0003500307, 0.0002934778, 0.0002597494, 0.000198476, 
    0.000178719, 0.0001594388, 0.0001431628, 0.0001285239, 0.0001161102, 
    0.0001041575, 9.468432e-005, 8.692776e-005, 8.398724e-005, 8.579924e-005, 
    8.606946e-005, 9.040868e-005, 9.191867e-005, 9.059942e-005, 
    8.811986e-005, 0.0001032197, 9.957983e-005, 9.559029e-005, 8.36058e-005, 
    8.047458e-005, 8.86126e-005, 8.818343e-005, 9.366707e-005, 0.0001034581, 
    0.0001174454, 0.0001320366, 0.0001431628, 0.0001529697, 0.0001635555, 
    0.0001806899, 0.0002013369, 0.0002209667, 0.0002329989, 0.0002372904, 
    0.0002442999, 0.0002460324, 0.0002505465, 0.0002591455, 0.0002686345, 
    0.0002768679, 0.0002793793, 0.0002762639, 0.0002744043, 0.0001992706, 
    0.0001780196, 0.0001616799, 0.0001537326, 0.000156244, 0.0001650178, 
    0.0002251152, 0.0001794342, 0.0001707557, 0.0001915459, 0.0001415415, 
    0.0001343254, 0.0001362804, 0.0001520955, 0.0002173745, 0.0002516591, 
    0.0002882325, 0.000325537, 0.0002392614, 0.0002053265, 0.0001642708, 
    0.0001265053, 9.555851e-005, 7.346504e-005, 7.349682e-005, 0.0001067165, 
    0.000178258, 0.0002839569, 0.0004718309, 0.0006487532, 0.0008752032, 
    0.001163785, 0.001058038,
  0.0009675984, 0.0008187774, 0.0006281375, 0.0005332949, 0.0005695981, 
    0.0008259615, 0.00110852, 0.00101037, 0.0009666447, 0.0008609457, 
    0.000765753, 0.0006896181, 0.0006188397, 0.0005415285, 0.0004710996, 
    0.0004147056, 0.0003626351, 0.0003218813, 0.000290585, 0.0002635007, 
    0.0002445543, 0.0002252265, 0.0002075994, 0.0001931194, 0.0001846477, 
    0.0001503789, 0.0001403335, 0.0001248045, 0.0001167619, 0.0001109444, 
    0.0001067642, 0.00011886, 0.0001161102, 0.0001169844, 0.0001183195, 
    0.0001191937, 0.000120513, 0.0001222296, 0.0001238509, 0.0001238191, 
    0.0001219117, 0.0001190507, 0.0001165553, 0.0001139803, 0.0001117869, 
    0.0001095934, 0.0001076066, 0.000107702, 0.0001112782, 0.0001180811, 
    0.0001284603, 0.0001430515, 0.0001585328, 0.0001727744, 0.0001817866, 
    0.0001837098, 0.0001802289, 0.0001740301, 0.000168308, 0.0001661146, 
    0.0001683557, 0.0001716459, 0.0001745387, 0.0001766367, 0.0001842185, 
    0.0001426064, 0.0001341028, 0.0001274907, 0.0001241687, 0.0001234376, 
    0.0001245184, 0.0001245661, 0.0001274271, 0.0001307332, 0.0001339439, 
    0.0001597408, 0.0001622044, 0.0001768116, 0.0001364235, 0.0001348181, 
    0.000133022, 0.0001284285, 0.0001228972, 0.0001180811, 0.0001132492, 
    0.0001062238, 9.918246e-005, 9.975469e-005, 0.0001150294, 0.0001545592, 
    0.0002148791, 0.0002930804, 0.0004231774, 0.0005304659, 0.0006519957, 
    0.0008000854,
  0.0005092149, 0.0005382064, 0.0005644007, 0.0005956652, 0.000465632, 
    0.0004477029, 0.0004235432, 0.0004604503, 0.0004332865, 0.0004078075, 
    0.0003857935, 0.0003671808, 0.0003516995, 0.0003371084, 0.0003217225, 
    0.0003066067, 0.000289377, 0.0002701605, 0.0002493545, 0.0002290094, 
    0.0002100471, 0.0001933419, 0.000179164, 0.0001695478, 0.0001695955, 
    0.0001382354, 0.0001369003, 0.0001505379, 0.000153526, 0.0001516028, 
    0.0001498861, 0.0001441005, 0.0001365506, 0.0001285874, 0.0001201474, 
    0.0001110398, 0.0001025362, 9.59241e-005, 9.069479e-005, 8.724567e-005, 
    8.579926e-005, 8.600589e-005, 8.819933e-005, 9.206171e-005, 
    9.690956e-005, 0.0001024091, 0.0001079722, 0.0001137419, 0.0001199408, 
    0.0001264258, 0.0001314167, 0.0001350724, 0.0001361532, 0.0001342141, 
    0.0001297795, 0.0001241369, 0.0001189394, 0.0001154426, 0.0001147592, 
    0.0001179381, 0.0001252178, 0.0001347228, 0.0001456582, 0.0001553698, 
    0.0001621409, 0.0001614574, 0.0001584533, 0.0001524452, 0.0001436078, 
    0.0001365029, 0.0001375043, 0.0001001679, 0.0001019163, 0.000100152, 
    0.0001032038, 0.0001072887, 0.0001103564, 0.0001120094, 0.0001131061, 
    0.0001122478, 0.0001094503, 0.0001056674, 0.0001016461, 9.824471e-005, 
    9.660755e-005, 9.772017e-005, 0.0001025362, 0.000112073, 0.0001286987, 
    0.0001530015, 0.000187143, 0.0002306783, 0.0003200217, 0.0003660047, 
    0.0004192037, 0.0004677618,
  0.0003039046, 0.0003164613, 0.0003248536, 0.0003298922, 0.0003279849, 
    0.0003263636, 0.0003246788, 0.0003169222, 0.000307608, 0.000298866, 
    0.0002908233, 0.0002838456, 0.0002766613, 0.0002686504, 0.0002598607, 
    0.0002496882, 0.0002381805, 0.0002259576, 0.0002137823, 0.0002015912, 
    0.0001901789, 0.0001802766, 0.0001719637, 0.0001653834, 0.0001607103, 
    0.0001570387, 0.0001557512, 0.0001537326, 0.000151571, 0.0001510464, 
    0.0001504743, 0.000148408, 0.0001451973, 0.0001417323, 0.0001375043, 
    0.000133626, 0.0001293981, 0.0001254244, 0.0001217528, 0.0001192414, 
    0.000117795, 0.0001170957, 0.0001170321, 0.0001175407, 0.0001184149, 
    0.000119305, 0.0001198295, 0.0001199408, 0.0001197818, 0.0001191779, 
    0.0001178586, 0.0001158241, 0.0001137737, 0.0001117869, 0.0001103723, 
    0.000109959, 0.0001103723, 0.0001121207, 0.000115236, 0.0001190507, 
    0.0001241369, 0.0001298908, 0.0001349612, 0.0001389666, 0.0001414938, 
    0.0001424634, 0.0001419071, 0.0001398408, 0.0001367891, 0.0001333081, 
    0.0001297636, 0.0001248681, 0.0001238826, 0.0001231197, 0.0001233104, 
    0.0001257582, 0.0001266483, 0.0001261556, 0.0001285556, 0.0001321001, 
    0.0001321955, 0.0001337691, 0.0001351837, 0.0001371228, 0.0001399679, 
    0.0001441005, 0.0001500928, 0.0001581672, 0.0001688484, 0.0001832648, 
    0.0002003832, 0.0002235257, 0.0002388163, 0.0002548698, 0.00027264, 
    0.0002890432,
  0.0002266888, 0.000230567, 0.0002335711, 0.0002361301, 0.0002378309, 
    0.0002398018, 0.0002406442, 0.0002407237, 0.0002403263, 0.000239468, 
    0.0002381487, 0.0002365275, 0.0002339208, 0.000230567, 0.0002269271, 
    0.0002233668, 0.0002194567, 0.0002150221, 0.0002109055, 0.0002064868, 
    0.0002023701, 0.0001983011, 0.0001944387, 0.000190465, 0.0001866185, 
    0.0001830899, 0.0001796408, 0.0001765096, 0.000173426, 0.0001708511, 
    0.0001685941, 0.000166337, 0.0001642548, 0.0001624906, 0.0001604084, 
    0.0001582944, 0.0001567685, 0.0001555446, 0.0001541936, 0.0001529061, 
    0.0001516505, 0.0001506332, 0.0001495842, 0.000148408, 0.0001473589, 
    0.0001462781, 0.0001452926, 0.0001444025, 0.0001435283, 0.0001428131, 
    0.0001423204, 0.0001418117, 0.0001409693, 0.0001405084, 0.0001400315, 
    0.0001398408, 0.0001395229, 0.0001393799, 0.0001394275, 0.0001393798, 
    0.0001396183, 0.0001401905, 0.0001405878, 0.0001412236, 0.0001418912, 
    0.0001423204, 0.0001425747, 0.0001432899, 0.0001438939, 0.0001442118, 
    0.0001447999, 0.0001452926, 0.0001461509, 0.0001473112, 0.0001485828, 
    0.000149918, 0.0001513962, 0.0001530333, 0.0001552268, 0.000157754, 
    0.0001603925, 0.0001633807, 0.0001666232, 0.0001702153, 0.0001740459, 
    0.0001778289, 0.000181866, 0.0001862688, 0.000190767, 0.0001957738, 
    0.0002008601, 0.0002057715, 0.0002104286, 0.0002148314, 0.00021836, 
    0.0002225085,
  8.114483e-005, 7.7648e-005, 7.451675e-005, 7.162393e-005, 6.898544e-005, 
    6.660129e-005, 6.445551e-005, 6.262763e-005, 6.100637e-005, 
    5.955997e-005, 5.839966e-005, 5.757312e-005, 5.682607e-005, 
    5.631744e-005, 5.603133e-005, 5.587241e-005, 5.574526e-005, 
    5.566579e-005, 5.547504e-005, 5.541148e-005, 5.542737e-005, 
    5.545915e-005, 5.558632e-005, 5.582473e-005, 5.612672e-005, 
    5.657178e-005, 5.730292e-005, 5.814534e-005, 5.943279e-005, 
    6.092688e-005, 6.285014e-005, 6.510718e-005, 6.784104e-005, 
    7.100408e-005, 7.459625e-005, 7.8554e-005, 8.28773e-005, 8.764566e-005, 
    9.281142e-005, 9.812019e-005, 0.0001034926, 0.0001091987, 0.0001147142, 
    0.000120325, 0.0001259357, 0.0001313081, 0.000136299, 0.0001409561, 
    0.0001451364, 0.0001487762, 0.0001518757, 0.0001540691, 0.0001554361, 
    0.0001566123, 0.0001562308, 0.0001562467, 0.0001547367, 0.0001530201, 
    0.0001506518, 0.0001478384, 0.0001453589, 0.0001423389, 0.0001398117, 
    0.000136601, 0.0001339466, 0.0001314035, 0.0001292418, 0.0001277159, 
    0.0001269689, 0.0001268577, 0.000127096, 0.000127414, 0.0001277477, 
    0.0001272391, 0.0001290352, 0.0001303862, 0.0001303862, 0.0001305451, 
    0.0001319121, 0.0001319916, 0.000131467, 0.0001305293, 0.0001291782, 
    0.0001272391, 0.0001252364, 0.0001228522, 0.0001199594, 0.0001168282, 
    0.0001132837, 0.000109469, 0.0001054317, 0.0001012197, 9.705534e-005, 
    9.292271e-005, 8.874244e-005, 8.489596e-005,
  9.918518e-005, 9.222334e-005, 8.570656e-005, 7.971426e-005, 7.419885e-005, 
    6.938282e-005, 6.491644e-005, 6.081564e-005, 5.704863e-005, 
    5.402866e-005, 5.172391e-005, 5.027752e-005, 4.932383e-005, 
    4.951458e-005, 5.013446e-005, 5.145372e-005, 5.285245e-005, 
    5.477569e-005, 5.652409e-005, 5.79864e-005, 5.868575e-005, 5.833608e-005, 
    5.695324e-005, 5.487105e-005, 5.212129e-005, 4.870397e-005, 
    4.563632e-005, 4.323623e-005, 4.228255e-005, 4.26958e-005, 4.503231e-005, 
    4.965761e-005, 5.638106e-005, 6.526614e-005, 7.626516e-005, 
    8.982324e-005, 0.000105686, 0.0001237105, 0.0001436264, 0.0001642575, 
    0.000184682, 0.0002052655, 0.000224625, 0.0002450018, 0.0002634554, 
    0.0002804785, 0.0002992182, 0.0003181487, 0.0003357122, 0.0003518294, 
    0.0003656258, 0.0003781824, 0.000385367, 0.000392599, 0.0003914069, 
    0.0003997039, 0.0003949355, 0.0003841749, 0.0003693292, 0.0003483962, 
    0.0003270338, 0.0003032873, 0.0002787142, 0.000255826, 0.0002341776, 
    0.0002149611, 0.0002005924, 0.0001900384, 0.0001859854, 0.0001846025, 
    0.0001876543, 0.0001908809, 0.0001960466, 0.0002011647, 0.0002057583, 
    0.0002101292, 0.0002120206, 0.0002135306, 0.0002112894, 0.0002083807, 
    0.0002045184, 0.0001956651, 0.0001938531, 0.0001847137, 0.0001833786, 
    0.0001786262, 0.0001763691, 0.0001717915, 0.0001656403, 0.0001583287, 
    0.0001498729, 0.000141099, 0.0001324366, 0.0001238853, 0.0001152069, 
    0.00010691,
  9.778643e-005, 8.828149e-005, 8.098585e-005, 7.586781e-005, 7.32452e-005, 
    7.186236e-005, 7.068619e-005, 6.935102e-005, 6.769798e-005, 
    6.532967e-005, 6.227792e-005, 5.855858e-005, 5.464851e-005, 
    5.113582e-005, 4.8545e-005, 4.730522e-005, 4.852911e-005, 5.094512e-005, 
    5.374257e-005, 5.609496e-005, 5.768442e-005, 5.811357e-005, 
    5.611086e-005, 5.216897e-005, 4.708271e-005, 4.202824e-005, 
    3.849964e-005, 3.714861e-005, 3.799103e-005, 4.110635e-005, 
    4.566809e-005, 5.121529e-005, 5.784335e-005, 6.561579e-005, 
    7.464393e-005, 8.562706e-005, 9.877188e-005, 0.0001152705, 0.0001356155, 
    0.0001600772, 0.0001875749, 0.0002155969, 0.000245288, 0.0002690821, 
    0.0002884099, 0.0003084212, 0.0003225675, 0.0003381284, 0.0003555646, 
    0.0003703149, 0.0003834596, 0.0003999264, 0.0004136115, 0.000421988, 
    0.0004215904, 0.0004118312, 0.0003970334, 0.0003811707, 0.000365133, 
    0.0003489525, 0.0003369681, 0.0003269067, 0.0003176082, 0.0003083736, 
    0.0003019203, 0.0003005058, 0.0002959758, 0.0002948631, 0.0002929717, 
    0.0002899835, 0.0002885688, 0.0002881716, 0.0002868681, 0.0002872973, 
    0.0002866774, 0.0002876311, 0.0002803673, 0.0002770771, 0.0002738188, 
    0.0002649496, 0.0002574315, 0.0002532194, 0.0002561281, 0.000260213, 
    0.0002660941, 0.0002666821, 0.0002646794, 0.0002648542, 0.0002550791, 
    0.0002366097, 0.0002178539, 0.0001920253, 0.0001681992, 0.0001466145, 
    0.0001270006, 0.0001105498,
  9.511615e-005, 9.204852e-005, 9.034778e-005, 8.670788e-005, 8.187594e-005, 
    7.553402e-005, 7.125837e-005, 6.893776e-005, 6.885828e-005, 
    6.933515e-005, 6.928747e-005, 6.912851e-005, 6.92239e-005, 6.989145e-005, 
    7.249814e-005, 7.717113e-005, 8.217798e-005, 8.559533e-005, 
    8.360852e-005, 7.969839e-005, 7.370618e-005, 6.359725e-005, 
    5.108819e-005, 3.981893e-005, 3.250744e-005, 3.094977e-005, 
    3.265048e-005, 3.78003e-005, 4.557277e-005, 5.406047e-005, 6.04183e-005, 
    6.493235e-005, 6.6188e-005, 6.41535e-005, 5.936921e-005, 5.40287e-005, 
    5.196242e-005, 5.390152e-005, 6.292964e-005, 7.955538e-005, 0.0001057496, 
    0.0001396686, 0.0001837759, 0.0002322226, 0.0002787779, 0.0003202945, 
    0.0003616683, 0.0003820771, 0.0004447018, 0.0004371359, 0.0004412046, 
    0.0004443675, 0.0004533003, 0.0004543494, 0.0004449559, 0.0004295697, 
    0.0003984321, 0.0003646248, 0.0003475699, 0.0003327718, 0.0003251424, 
    0.0003288616, 0.0003321043, 0.0003373495, 0.0003439139, 0.0003522745, 
    0.0003619861, 0.000371952, 0.0003781032, 0.0003782621, 0.0003745745, 
    0.0003735413, 0.0003710458, 0.0003716022, 0.0003715865, 0.0003721745, 
    0.000367867, 0.0003676604, 0.0003673585, 0.0003751151, 0.0004370719, 
    0.0004629166, 0.0004811636, 0.000498886, 0.0005118243, 0.0005204552, 
    0.0005055621, 0.0004873787, 0.000451997, 0.0003306419, 0.0002783648, 
    0.0002260079, 0.0001814554, 0.0001460582, 0.0001181951, 0.0001018078,
  0.0001750499, 0.000176083, 0.0001751293, 0.0001639077, 0.0001495074, 
    0.0001363307, 0.0001309265, 0.0001360764, 0.0001460582, 0.0001469642, 
    0.0001372049, 0.0001224706, 0.00010478, 9.165116e-005, 8.834506e-005, 
    9.36221e-005, 0.0001060675, 0.0001163354, 0.0001170982, 0.0001060038, 
    0.0001001864, 9.279541e-005, 7.81407e-005, 6.038649e-005, 4.501641e-005, 
    3.705325e-005, 3.540024e-005, 3.562277e-005, 3.697377e-005, 
    3.832483e-005, 3.791155e-005, 3.964407e-005, 4.48098e-005, 5.229615e-005, 
    6.292967e-005, 7.157624e-005, 7.585189e-005, 7.558172e-005, 
    7.616982e-005, 8.303617e-005, 9.688025e-005, 0.0001203885, 0.0001479337, 
    0.0001771479, 0.0002058059, 0.0002273114, 0.000300681, 0.000242332, 
    0.0001906746, 0.0001524324, 0.0001383813, 0.0001407494, 0.0001676907, 
    0.0002015617, 0.0002326355, 0.0002599587, 0.0002994724, 0.0003518451, 
    0.0003996559, 0.000436547, 0.0004550961, 0.0004573851, 0.0004303481, 
    0.0003753849, 0.0003194835, 0.0002779192, 0.0002583372, 0.0002811777, 
    0.0003078487, 0.0003455349, 0.0004439384, 0.0005328525, 0.0005190878, 
    0.0004528393, 0.0003833801, 0.0003381122, 0.0003794227, 0.0003674697, 
    0.0003668499, 0.0003694727, 0.0003825062, 0.0004057598, 0.0004407279, 
    0.0004693381, 0.0005023035, 0.0005422465, 0.0005773415, 0.0006037266, 
    0.0006244374, 0.0006368191, 0.0006413014, 0.000447467, 0.0003624629, 
    0.0002870433, 0.000222066, 0.0001866371,
  0.0003907867, 0.0003522108, 0.000285676, 0.0002535055, 0.0002115757, 
    0.0001946003, 0.0002093188, 0.000255572, 0.0002966436, 0.0003236325, 
    0.0003276856, 0.0003080083, 0.0002663803, 0.0002130857, 0.0001636057, 
    0.0001301636, 0.0001143484, 0.0001094689, 0.0001094849, 0.0001024436, 
    9.424181e-005, 9.700749e-005, 0.0001018395, 9.842229e-005, 9.875605e-005, 
    0.0001030157, 0.0001157313, 0.0001331836, 0.0001526704, 0.0001608562, 
    0.0001458199, 0.0001187831, 9.516376e-005, 8.073152e-005, 7.930095e-005, 
    7.69645e-005, 6.633101e-005, 4.682847e-005, 3.398571e-005, 4.822714e-005, 
    7.774332e-005, 0.0001191011, 0.0001476796, 0.0001587899, 0.0001575185, 
    0.0001095803, 0.000121024, 0.0001108511, 6.903242e-005, 3.986596e-005, 
    3.004307e-005, 4.183664e-005, 6.054481e-005, 7.192511e-005, 
    8.406863e-005, 0.0001111529, 0.0001525106, 0.0002011321, 0.0002343995, 
    0.0002545856, 0.0002715769, 0.0002902215, 0.0003010298, 0.0002932095, 
    0.0002837521, 0.000273834, 0.0002833391, 0.0003061157, 0.0003384454, 
    0.0003719828, 0.0003712834, 0.0003253485, 0.0002830373, 0.0002688747, 
    0.000249404, 0.0002237661, 0.0001982076, 0.0001992725, 0.000318689, 
    0.0003682962, 0.0004195082, 0.0004495012, 0.0004603891, 0.0004633453, 
    0.0004907632, 0.0005393689, 0.0005848911, 0.0006110219, 0.0006336239, 
    0.0006594686, 0.0006806878, 0.0006920206, 0.0006800042, 0.000632464, 
    0.0005585542, 0.0004785722,
  0.0006196524, 0.000678367, 0.000720615, 0.0007083444, 0.0006783195, 
    0.0006480564, 0.0006315892, 0.0006270912, 0.0005969231, 0.0005707925, 
    0.0005760854, 0.0005965417, 0.0006144072, 0.0006265824, 0.0006007536, 
    0.0005489695, 0.0005043691, 0.0004732953, 0.0004493261, 0.0004190311, 
    0.0003630028, 0.000285628, 0.0002354011, 0.0002206352, 0.000202738, 
    0.0002079196, 0.0001918343, 0.0001993843, 0.0002078242, 0.0002121155, 
    0.0002068703, 0.0001925651, 0.0001866368, 0.000262693, 0.0002577339, 
    0.0002545386, 0.0003986068, 0.0002626763, 0.0002398512, 0.0002292814, 
    0.0002203172, 0.0002289158, 0.0002305054, 0.0001973019, 0.0001302105, 
    4.522246e-005, -3.329664e-005, -9.387126e-005, -0.0001149946, 
    -0.0001149317, -7.746788e-005, -1.177518e-005, 3.420748e-005, 
    4.108972e-005, 2.074498e-005, 2.686447e-005, 9.153946e-005, 0.0001644953, 
    0.0002103511, 0.0002488003, 0.0002922718, 0.0003335658, 0.0003713476, 
    0.0003988133, 0.0004176483, 0.0004330184, 0.0004606275, 0.0004653325, 
    0.0004611043, 0.0004457501, 0.0004236568, 0.0004097805, 0.0003993856, 
    0.0003913585, 0.0003734133, 0.0003521624, 0.0003233296, 0.0003169402, 
    0.0004143105, 0.0005269716, 0.000457814, 0.0003702345, 0.0003226621, 
    0.0003365858, 0.0003814083, 0.0004216693, 0.0004584016, 0.000480829, 
    0.0004924005, 0.0004966762, 0.0004868056, 0.0004940217, 0.0005161627, 
    0.0005327251, 0.0005421822, 0.000571047,
  0.0004264538, 0.000401404, 0.0003853822, 0.0003823785, 0.000382839, 
    0.0003829978, 0.0003833636, 0.0003878295, 0.0003849526, 0.0003942675, 
    0.0004259297, 0.000488284, 0.0005428661, 0.0005598096, 0.0005513537, 
    0.0005418486, 0.0005402118, 0.0005299598, 0.0005108698, 0.0004678434, 
    0.0004218447, 0.000384588, 0.0003604435, 0.0003424035, 0.0003198648, 
    0.0002904441, 0.0002477034, 0.0002004965, 0.0001568189, 0.0001388416, 
    0.0001370939, 0.0001621759, 0.0002100663, 0.0002657766, 0.0003048293, 
    0.0003358875, 0.0003843815, 0.0003868295, 0.0003835871, 0.0003797086, 
    0.0003584735, 0.0003350293, 0.0003328994, 0.0003250157, 0.0002786829, 
    0.0001871935, 5.468074e-005, -4.679011e-005, -8.68924e-005, -0.000129601, 
    -0.0001611197, -0.0001536966, -0.0001283609, -0.0001019598, 
    -7.60844e-005, -2.485607e-005, 5.49024e-005, 0.0001243302, 0.0001715692, 
    0.0002447958, 0.0003400999, 0.0004164255, 0.0004487708, 0.0004893178, 
    0.0005676304, 0.0006389492, 0.0006895261, 0.0007100618, 0.0007086946, 
    0.000693833, 0.000701224, 0.000702925, 0.0006810538, 0.0006607566, 
    0.0006434158, 0.0006253594, 0.0006046486, 0.0005713021, 0.0005387976, 
    0.0005209479, 0.0005173874, 0.0004877918, 0.0003977325, 0.0003496832, 
    0.000375194, 0.0003957937, 0.0004351162, 0.0004784607, 0.000492353, 
    0.000497916, 0.000489492, 0.0004715309, 0.0004561925, 0.0004515992, 
    0.0004463696, 0.0004418555,
  0.0004424755, 0.0004085409, 0.0003847783, 0.0003662771, 0.0003502867, 
    0.0003277962, 0.0003271452, 0.0003403532, 0.0003536581, 0.0003628763, 
    0.0003981148, 0.000436977, 0.0004697358, 0.0004912256, 0.0005255258, 
    0.0005490812, 0.00055501, 0.000557553, 0.0005556145, 0.000521536, 
    0.0004759664, 0.0004302533, 0.0004053628, 0.0004074452, 0.0004015001, 
    0.0003816797, 0.0003574565, 0.0003305152, 0.0003068801, 0.0002805111, 
    0.0002397094, 0.0001846505, 0.0001445487, 0.0001315633, 0.0001464565, 
    0.0001506051, 0.0001781345, 0.0002593077, 0.0003627338, 0.0004420793, 
    0.0004663342, 0.0004767133, 0.0004922906, 0.0004725335, 0.0004267893, 
    0.0003867988, 0.0003115223, 0.0001665158, 1.165457e-005, -0.0001149615, 
    -0.0001923204, -0.00021702, -0.0001935121, -0.0001581311, -0.0001322548, 
    -6.583147e-005, 3.37637e-005, 0.0001011086, 0.0001135389, 0.0002055047, 
    0.0003621145, 0.0004541436, 0.0004941183, 0.0005841772, 0.0007302007, 
    0.0008130269, 0.0008446099, 0.0008793077, 0.0009211898, 0.0009481949, 
    0.0009618956, 0.000957239, 0.0009394051, 0.0009237807, 0.0009038015, 
    0.0008462952, 0.0007397849, 0.0006670831, 0.0006502667, 0.0006598677, 
    0.000662935, 0.0006543831, 0.0005902164, 0.0004659849, 0.0003836667, 
    0.0003874023, 0.0004474195, 0.0004831501, 0.0004677484, 0.000469306, 
    0.0005168309, 0.0005243807, 0.0005027801, 0.0004801615, 0.0004681135, 
    0.0004655388,
  0.0005026534, 0.000505276, 0.0005280846, 0.0005198671, 0.0005052919, 
    0.0005105692, 0.0005348083, 0.0005329642, 0.0005139704, 0.0005112207, 
    0.0005235709, 0.0005372721, 0.0005571879, 0.0005856389, 0.0006343084, 
    0.0006824844, 0.0007357313, 0.0007865941, 0.000768045, 0.0006290469, 
    0.0005299761, 0.0004881895, 0.0004541753, 0.0004356741, 0.0004330198, 
    0.0004517911, 0.0004571159, 0.0004514572, 0.000438917, 0.0004264871, 
    0.0004120865, 0.0003814897, 0.0003526574, 0.0003370331, 0.0003212173, 
    0.0003295937, 0.0003642915, 0.0004203361, 0.0004850426, 0.0005224105, 
    0.0005412139, 0.0005674721, 0.0005992125, 0.0005879593, 0.0005911062, 
    0.0006011836, 0.0005399575, 0.0003810115, 0.0002061557, 0.000105225, 
    6.517069e-005, 6.240513e-005, 8.136733e-005, 9.794533e-005, 0.0001010937, 
    0.0001203576, 0.0001630187, 0.0002183476, 0.00026805, 0.0003757039, 
    0.0005027801, 0.0005694898, 0.0006326227, 0.0007603038, 0.0008746972, 
    0.0008971877, 0.0009079962, 0.0009746263, 0.001023343, 0.001013838, 
    0.0009970539, 0.0009981347, 0.00101546, 0.00099672, 0.0009204098, 
    0.0007878812, 0.0007291189, 0.0008444018, 0.0008685458, 0.0007783286, 
    0.000750402, 0.0006778119, 0.0005879286, 0.0004582601, 0.000418222, 
    0.0005051815, 0.0006118175, 0.0006441944, 0.0005926322, 0.0005784864, 
    0.0005951757, 0.0005945242, 0.0005687433, 0.0005559479, 0.0005373191, 
    0.0005139546,
  0.0007580956, 0.0007850518, 0.0008013924, 0.0008157925, 0.0008249315, 
    0.0008438146, 0.0008533513, 0.0008379025, 0.0008184314, 0.000841192, 
    0.000883806, 0.0009010993, 0.0009042937, 0.0009274525, 0.00095673, 
    0.0009751837, 0.001039954, 0.00110323, 0.001078451, 0.0009646458, 
    0.0009154356, 0.0009094439, 0.0008503003, 0.0007491312, 0.0006953916, 
    0.000705834, 0.0006930232, 0.0006644446, 0.0006317971, 0.0006083529, 
    0.000581014, 0.0005712709, 0.0005840017, 0.0005530068, 0.0005185325, 
    0.0005257321, 0.000555343, 0.0005771192, 0.0006126435, 0.0006714379, 
    0.0007252567, 0.0007581105, 0.0007463004, 0.0007284824, 0.0007275767, 
    0.0007316615, 0.0006492962, 0.0005114744, 0.0003740187, 0.0003251107, 
    0.0003593946, 0.0004079053, 0.0004541269, 0.0004986469, 0.0005221236, 
    0.0005399575, 0.0005592853, 0.000587116, 0.000636294, 0.0006817682, 
    0.0007215044, 0.000778852, 0.0008514905, 0.0009168973, 0.0009725909, 
    0.000998531, 0.001011263, 0.001021626, 0.001039047, 0.001034771, 
    0.001012471, 0.000996083, 0.0009679184, 0.0009427583, 0.0008750618, 
    0.0008253753, 0.0009022267, 0.0009748167, 0.0009550275, 0.001004381, 
    0.0008915928, 0.0006443369, 0.0004962804, 0.000460708, 0.0005469997, 
    0.0006834068, 0.0007866104, 0.0008295742, 0.0008349936, 0.0008583427, 
    0.0008534472, 0.0008162218, 0.0007830183, 0.0007592561, 0.0007510697, 
    0.0007401342,
  0.00100373, 0.001030639, 0.001042909, 0.001074953, 0.001103913, 
    0.001142902, 0.001231038, 0.001312274, 0.001318712, 0.001322987, 
    0.001332111, 0.001367603, 0.001414731, 0.001426843, 0.001414095, 
    0.001407309, 0.001450113, 0.001483427, 0.001471348, 0.001532956, 
    0.001652179, 0.001628799, 0.001446409, 0.001275065, 0.001192191, 
    0.001152089, 0.001109015, 0.001020689, 0.0009178193, 0.0008453401, 
    0.0008403324, 0.0008687521, 0.0008749035, 0.0008420972, 0.0008058725, 
    0.000795478, 0.0007870859, 0.0008001663, 0.0008320026, 0.0008802749, 
    0.0009580795, 0.0009670118, 0.0009595891, 0.0009987056, 0.001075176, 
    0.001123478, 0.001108489, 0.001040476, 0.0008997461, 0.0008555762, 
    0.0009245574, 0.0009837328, 0.0009869281, 0.0009549959, 0.0009026546, 
    0.0009148465, 0.0009474456, 0.0009950502, 0.001045626, 0.001042606, 
    0.001031162, 0.001074221, 0.001125274, 0.001132363, 0.001180477, 
    0.00124655, 0.001230656, 0.00119502, 0.001190934, 0.001146541, 
    0.001080181, 0.001005318, 0.0009699687, 0.0009624185, 0.0009245574, 
    0.0009210287, 0.0009814757, 0.0009445697, 0.0008660979, 0.001164868, 
    0.00108007, 0.000800183, 0.0006737728, 0.0007612575, 0.0009289766, 
    0.001064112, 0.001111128, 0.001094853, 0.001090244, 0.001083933, 
    0.001068643, 0.001066878, 0.001056038, 0.001038061, 0.001020911, 
    0.0009996286,
  0.001323241, 0.001365266, 0.001424616, 0.001499305, 0.001578285, 
    0.001721559, 0.001926011, 0.002073258, 0.002170184, 0.002268014, 
    0.002383044, 0.002418917, 0.002304492, 0.002152573, 0.002050958, 
    0.002030263, 0.002051705, 0.002051451, 0.002047351, 0.002066853, 
    0.00201564, 0.001829546, 0.001591048, 0.00143657, 0.001346861, 
    0.001296316, 0.001274969, 0.001212488, 0.001148384, 0.001118455, 
    0.001111128, 0.001127054, 0.001152914, 0.001137831, 0.001142759, 
    0.001145953, 0.001109888, 0.001088399, 0.001065033, 0.001157445, 
    0.001450112, 0.001512563, 0.001434059, 0.001436967, 0.001513817, 
    0.001549041, 0.001472985, 0.001513294, 0.001559134, 0.001630277, 
    0.001694158, 0.001625366, 0.0015262, 0.001415574, 0.00134187, 0.0013488, 
    0.001349262, 0.001314134, 0.001307522, 0.001293376, 0.001303946, 
    0.001355127, 0.001388458, 0.001415732, 0.001472206, 0.001474225, 
    0.001447887, 0.001416623, 0.001352838, 0.001287511, 0.001237109, 
    0.00117903, 0.001137386, 0.001066528, 0.0009548059, 0.0009127175, 
    0.0009252094, 0.0007887231, 0.0008023605, 0.001301037, 0.001244993, 
    0.001128915, 0.001217766, 0.00134853, 0.001408851, 0.001454085, 
    0.00144466, 0.001404971, 0.00139866, 0.001390364, 0.001375502, 
    0.001367523, 0.001332587, 0.001321399, 0.001351216, 0.001327374,
  0.00139809, 0.001415669, 0.00149244, 0.001614558, 0.001853071, 0.002160472, 
    0.002320325, 0.002579374, 0.002839791, 0.002851314, 0.00258058, 
    0.002300424, 0.002089789, 0.001989097, 0.001966272, 0.002017152, 
    0.00207593, 0.002044681, 0.00197306, 0.0018693, 0.001718, 0.001596374, 
    0.001497987, 0.001414158, 0.001362072, 0.001324751, 0.001296095, 
    0.001275034, 0.001296317, 0.001363026, 0.00140742, 0.001398503, 
    0.001377729, 0.001317695, 0.001369733, 0.001429704, 0.001398264, 
    0.001391668, 0.001398153, 0.001872876, 0.002041995, 0.002308243, 
    0.002268666, 0.002102123, 0.002076088, 0.002064675, 0.00205374, 
    0.002086452, 0.001956036, 0.001992896, 0.001952191, 0.001870841, 
    0.001786807, 0.001767844, 0.00175082, 0.001712451, 0.001631818, 
    0.001598679, 0.001589761, 0.001558783, 0.00157064, 0.001623298, 
    0.001634727, 0.001628337, 0.001639272, 0.001642101, 0.001654834, 
    0.001634615, 0.001516201, 0.001397373, 0.001303119, 0.001217669, 
    0.001136702, 0.00105038, 0.0009584939, 0.0009929361, 0.001025504, 
    0.001240574, 0.001578079, 0.001764253, 0.001510337, 0.001532415, 
    0.00169956, 0.001775363, 0.0017842, 0.001812619, 0.001798473, 
    0.001777477, 0.001804386, 0.001814337, 0.001774219, 0.001759739, 
    0.001688881, 0.001566635, 0.001495014, 0.001435728,
  0.001358797, 0.001365363, 0.001477865, 0.001674894, 0.001892299, 
    0.00218104, 0.002588179, 0.002730022, 0.002649135, 0.002468701, 
    0.002016404, 0.00194135, 0.001960694, 0.001975778, 0.002007154, 
    0.002052087, 0.002093159, 0.002036955, 0.001891075, 0.001757766, 
    0.001612952, 0.00153143, 0.00149681, 0.001443676, 0.001372149, 
    0.001357859, 0.001353504, 0.001420992, 0.001537977, 0.001675623, 
    0.001709719, 0.001765413, 0.001737867, 0.001572247, 0.001602398, 
    0.001587537, 0.001434091, 0.002035667, 0.002203118, 0.002740275, 
    0.002755263, 0.002790628, 0.002951116, 0.002699918, 0.002562525, 
    0.002599465, 0.002506434, 0.002351987, 0.002228089, 0.002083528, 
    0.001995789, 0.001975158, 0.00195715, 0.001898419, 0.001857539, 
    0.001798857, 0.001735659, 0.001812382, 0.001896877, 0.001894398, 
    0.001842326, 0.001830357, 0.0018398, 0.001811921, 0.001766907, 
    0.001709607, 0.001686958, 0.001617419, 0.001450381, 0.001286351, 
    0.00117272, 0.001085823, 0.001076588, 0.001055228, 0.0009481618, 
    0.001038713, 0.001184243, 0.001955894, 0.002168849, 0.001947151, 
    0.00172043, 0.001872415, 0.002000477, 0.00215305, 0.002210763, 
    0.002099437, 0.002061306, 0.002111136, 0.002167912, 0.002157738, 
    0.002024208, 0.001872207, 0.001738407, 0.001603796, 0.001481598, 
    0.001411377,
  0.001435617, 0.001481981, 0.00148187, 0.001693855, 0.00208893, 0.001936503, 
    0.002438566, 0.002749731, 0.002428249, 0.00220577, 0.002218551, 
    0.002477839, 0.002604264, 0.002558312, 0.002592629, 0.002582536, 
    0.002578086, 0.002462263, 0.002268031, 0.002118925, 0.001995121, 
    0.001882843, 0.001828292, 0.001722991, 0.001682093, 0.001704379, 
    0.001760041, 0.001854901, 0.00186706, 0.00185962, 0.001925504, 
    0.002264821, 0.001786347, 0.0013591, 0.001211392, 0.00134249, 
    0.001880601, 0.00226784, 0.002613675, 0.003189487, 0.002966087, 
    0.002636863, 0.002409158, 0.002432205, 0.002550954, 0.002699203, 
    0.002634495, 0.002421129, 0.00239282, 0.002399114, 0.002352178, 
    0.002337935, 0.002271161, 0.002147186, 0.002067139, 0.002018645, 
    0.001997807, 0.002034906, 0.001998634, 0.001942844, 0.00184487, 
    0.001821758, 0.001836812, 0.001780989, 0.00176225, 0.001695, 0.001582927, 
    0.001384977, 0.001249317, 0.001149943, 0.001068865, 0.001082344, 
    0.001036662, 0.001025283, 0.0009456174, 0.001083313, 0.001222057, 
    0.001625349, 0.002330719, 0.002528718, 0.00255259, 0.002538143, 
    0.002305812, 0.002464059, 0.002538875, 0.002470639, 0.002558853, 
    0.00261337, 0.002538525, 0.002380261, 0.002149711, 0.001901328, 
    0.00176117, 0.001639465, 0.001565587, 0.001493839,
  0.001610791, 0.00163182, 0.00170077, 0.002051579, 0.002444986, 0.002316811, 
    0.002817173, 0.002772796, 0.002392136, 0.002359821, 0.002548918, 
    0.002839344, 0.002937287, 0.002951767, 0.002992744, 0.002953263, 
    0.002906453, 0.002800517, 0.002619268, 0.002481097, 0.00231875, 
    0.00220674, 0.002147771, 0.002041247, 0.00199795, 0.00196899, 0.00190708, 
    0.00202416, 0.002171806, 0.002418568, 0.00274002, 0.002740578, 
    0.002434765, 0.001500688, 0.0009024963, 0.001136989, 0.001856807, 
    0.00260595, 0.003334478, 0.003405366, 0.002831906, 0.002539271, 
    0.002192022, 0.002357343, 0.002555532, 0.002846515, 0.002956918, 
    0.002851013, 0.002792694, 0.002845401, 0.00291316, 0.00280595, 
    0.002643729, 0.002479251, 0.002410255, 0.002329385, 0.002196345, 
    0.002102187, 0.001914408, 0.00183012, 0.001773773, 0.001787458, 
    0.001779271, 0.001633057, 0.00157943, 0.001454245, 0.001397341, 
    0.001236872, 0.001184736, 0.001170813, 0.00101484, 0.001093645, 
    0.0009845924, 0.001044055, 0.0009848941, 0.001191317, 0.001404145, 
    0.0008744267, 0.002783555, 0.003020797, 0.003007002, 0.002984257, 
    0.002730482, 0.002701335, 0.002793329, 0.002835736, 0.002854621, 
    0.002686378, 0.002507372, 0.002301091, 0.002132483, 0.002021634, 
    0.001903123, 0.001736072, 0.001682952, 0.001636364,
  0.00187607, 0.001943829, 0.002206377, 0.002630729, 0.00246762, 0.0022532, 
    0.002721298, 0.00277424, 0.002616996, 0.002397031, 0.002815453, 
    0.003173288, 0.003148368, 0.002979325, 0.002992518, 0.002942307, 
    0.002863519, 0.002769232, 0.002608489, 0.002462704, 0.002281446, 
    0.002240278, 0.002250243, 0.002232252, 0.002225338, 0.002251088, 
    0.002275866, 0.002516286, 0.002732772, 0.002952654, 0.003286537, 
    0.003261807, 0.002442695, 0.001756687, 0.001650733, 0.001743414, 
    0.002378037, 0.003262762, 0.00341015, 0.003325749, 0.002626961, 
    0.002703652, 0.002732515, 0.002873722, 0.002935154, 0.003152911, 
    0.003282102, 0.003200864, 0.003155533, 0.003123123, 0.003158251, 
    0.003103193, 0.002963431, 0.002823927, 0.002741113, 0.002613004, 
    0.002399428, 0.002309561, 0.002143096, 0.002043184, 0.001968844, 
    0.0018219, 0.00174338, 0.001594052, 0.001510765, 0.00134071, 0.001285776, 
    0.001266452, 0.001247837, 0.001230053, 0.001161706, 0.001157255, 
    0.001051127, 0.00114945, 0.001061728, 0.001547355, 0.002067251, 
    0.0007204562, 0.002801945, 0.003275063, 0.003506485, 0.003167503, 
    0.00288892, 0.002747951, 0.002627024, 0.002808427, 0.002834478, 
    0.002517859, 0.00233512, 0.00225649, 0.002154909, 0.002012048, 
    0.001919432, 0.001903854, 0.001882302, 0.001847637,
  0.002309325, 0.002364941, 0.002593791, 0.002940976, 0.002678841, 
    0.002671022, 0.002689365, 0.002499932, 0.00247725, 0.002415325, 
    0.00298354, 0.003345331, 0.002928736, 0.003012549, 0.003129689, 
    0.003032541, 0.002985684, 0.002892749, 0.002727747, 0.002650244, 
    0.002536949, 0.002587017, 0.002595266, 0.002565259, 0.002575638, 
    0.002703065, 0.002858419, 0.00308601, 0.003239855, 0.003356902, 
    0.003673365, 0.003710985, 0.002939736, 0.001756178, 0.002537904, 
    0.002702906, 0.003349006, 0.003776154, 0.003558479, 0.003315704, 
    0.003118467, 0.002996715, 0.003213741, 0.003231796, 0.003241681, 
    0.003368378, 0.003346825, 0.003250964, 0.003266335, 0.003212849, 
    0.003236802, 0.003289333, 0.003207574, 0.003106562, 0.002928449, 
    0.002822734, 0.002709975, 0.002628962, 0.002481492, 0.002306303, 
    0.002132829, 0.001882903, 0.001783388, 0.00166858, 0.001614828, 
    0.001544446, 0.00144404, 0.001435616, 0.001402905, 0.001406547, 
    0.001391872, 0.00133502, 0.001344382, 0.001415336, 0.001387917, 
    0.002011635, 0.002295242, 0.001265433, 0.002857131, 0.003344522, 
    0.003660535, 0.003331551, 0.003108708, 0.00295129, 0.002633637, 
    0.00301951, 0.002774414, 0.00258158, 0.002466727, 0.002382105, 
    0.002301902, 0.002211748, 0.002214704, 0.002197983, 0.002190021, 
    0.002205501,
  0.002714796, 0.00283507, 0.002947889, 0.003070261, 0.002842428, 
    0.002311392, 0.002612704, 0.002611003, 0.002713524, 0.002546709, 
    0.00285325, 0.00328983, 0.002894007, 0.002929037, 0.00323024, 
    0.003170412, 0.003167583, 0.003064219, 0.002944978, 0.00298365, 
    0.002883228, 0.00289968, 0.002900489, 0.002912935, 0.002960667, 
    0.003106054, 0.003255924, 0.003338385, 0.003435295, 0.00351561, 
    0.003633881, 0.003822967, 0.003808264, 0.003982957, 0.004048396, 
    0.004010996, 0.003922416, 0.003822885, 0.003653813, 0.003363863, 
    0.003347477, 0.003435533, 0.003496649, 0.003382128, 0.00337938, 
    0.003404301, 0.003325323, 0.003287015, 0.003249297, 0.003136573, 
    0.003142899, 0.003178187, 0.003119312, 0.003124271, 0.003048278, 
    0.003027694, 0.00300293, 0.002886774, 0.002780423, 0.002534786, 
    0.002311118, 0.002150392, 0.002171358, 0.00212992, 0.001993991, 
    0.001945879, 0.001861399, 0.001829086, 0.001818547, 0.001769164, 
    0.001732638, 0.00174909, 0.001812302, 0.001815083, 0.001869585, 
    0.002462978, 0.002095178, 0.002282909, 0.002570982, 0.003339611, 
    0.003408194, 0.003183316, 0.003002627, 0.003028221, 0.002939608, 
    0.00294851, 0.002799287, 0.002667379, 0.002651056, 0.002702696, 
    0.002664568, 0.002669988, 0.00265306, 0.00262747, 0.002705736, 0.002697884,
  0.003157714, 0.003228635, 0.003113635, 0.003012052, 0.002967837, 
    0.002685089, 0.002936158, 0.003047024, 0.002842427, 0.002765357, 
    0.002858307, 0.003274586, 0.00322544, 0.00316841, 0.003248757, 
    0.003195114, 0.003256196, 0.003227061, 0.003230987, 0.003243098, 
    0.003172271, 0.00316631, 0.003159825, 0.003196446, 0.003270006, 
    0.003353197, 0.00338467, 0.003375627, 0.003411232, 0.003454942, 
    0.003467973, 0.00346327, 0.003567271, 0.003522638, 0.003651414, 
    0.003689241, 0.003465684, 0.003674636, 0.003443781, 0.003352152, 
    0.00338928, 0.003559545, 0.003516294, 0.003353471, 0.003280532, 
    0.00327217, 0.003264541, 0.003337273, 0.003328755, 0.00310491, 
    0.003001153, 0.003071006, 0.003089542, 0.003040697, 0.003030382, 
    0.003074424, 0.003120504, 0.00308444, 0.003019542, 0.002841443, 
    0.00272239, 0.002579212, 0.002511185, 0.002571821, 0.002497783, 
    0.002401259, 0.002327142, 0.002283718, 0.002294907, 0.002318527, 
    0.002346534, 0.002396443, 0.0024306, 0.002484499, 0.002597811, 
    0.002879399, 0.002688539, 0.00228197, 0.002813549, 0.003292767, 
    0.003146743, 0.002873169, 0.002900871, 0.002938479, 0.002761891, 
    0.002733979, 0.002928574, 0.003019411, 0.002985097, 0.003007269, 
    0.003018633, 0.003021304, 0.003033815, 0.003081467, 0.003147842, 
    0.003123682,
  0.003427442, 0.003335031, 0.003220432, 0.003050502, 0.002902415, 
    0.002997669, 0.003051966, 0.003008177, 0.002821591, 0.002702953, 
    0.002908725, 0.00329485, 0.003282135, 0.003214933, 0.003225725, 
    0.003206939, 0.003344491, 0.003347574, 0.003384957, 0.003305802, 
    0.003331775, 0.003366219, 0.003361514, 0.003380237, 0.003380189, 
    0.003285473, 0.003278717, 0.00332831, 0.003465449, 0.003390236, 
    0.003310969, 0.003257262, 0.003292801, 0.003407577, 0.003345905, 
    0.003203044, 0.003070977, 0.003250331, 0.003207749, 0.002940848, 
    0.003047707, 0.003358208, 0.00344725, 0.003275955, 0.003161894, 
    0.003072582, 0.003049996, 0.003162498, 0.00323523, 0.003076429, 
    0.003061535, 0.003138816, 0.003120601, 0.003049806, 0.003103022, 
    0.003205778, 0.003225503, 0.003230017, 0.003194096, 0.003150465, 
    0.0030887, 0.002964243, 0.002867602, 0.002894815, 0.002881989, 
    0.002852837, 0.002850041, 0.002860326, 0.002851283, 0.002883866, 
    0.00292589, 0.002951704, 0.003041795, 0.003101604, 0.002999369, 
    0.002604025, 0.002449738, 0.002501744, 0.002902161, 0.003198942, 
    0.002830397, 0.002717879, 0.002572777, 0.002817424, 0.002806872, 
    0.002546631, 0.002745343, 0.003080733, 0.003091812, 0.003082896, 
    0.003145408, 0.00323019, 0.003324158, 0.003420783, 0.003425661, 
    0.003404412,
  0.003309043, 0.003287571, 0.003157647, 0.002957424, 0.002898712, 
    0.002770983, 0.002676552, 0.00281857, 0.002645208, 0.002757487, 
    0.002743596, 0.003245402, 0.003381712, 0.003403218, 0.003386419, 
    0.003394017, 0.003397642, 0.003361003, 0.003415331, 0.003349068, 
    0.003395019, 0.003410485, 0.003388898, 0.003373832, 0.003373515, 
    0.003339659, 0.003399359, 0.003242115, 0.003028091, 0.003303817, 
    0.003263351, 0.003269278, 0.003354331, 0.003259836, 0.003241558, 
    0.003391095, 0.003411392, 0.002970045, 0.002630061, 0.002810974, 
    0.002886076, 0.003213359, 0.003270168, 0.00316954, 0.003122602, 
    0.003046038, 0.003031287, 0.003011897, 0.00307069, 0.003088256, 
    0.003110906, 0.003101874, 0.003119009, 0.003219767, 0.003266957, 
    0.003343584, 0.003347605, 0.003336495, 0.00339823, 0.003437219, 
    0.003444785, 0.003376435, 0.003352705, 0.003322728, 0.003255844, 
    0.003279671, 0.003305307, 0.003247801, 0.003250552, 0.003338447, 
    0.003260262, 0.003243892, 0.003265731, 0.003221687, 0.00314296, 
    0.002821909, 0.002665491, 0.002699997, 0.002924714, 0.002982935, 
    0.002782729, 0.002711281, 0.002485389, 0.002133435, 0.002925906, 
    0.002819858, 0.002878904, 0.00301183, 0.003129708, 0.003152227, 
    0.003109027, 0.003195953, 0.003213406, 0.003324954, 0.003375547, 
    0.003300395,
  0.003004344, 0.002982076, 0.002919389, 0.002772683, 0.002848437, 0.0021568, 
    0.002164796, 0.002134118, 0.002606729, 0.002977516, 0.002529641, 
    0.003148986, 0.003339021, 0.003350861, 0.003440157, 0.003483152, 
    0.003445117, 0.003378885, 0.003381014, 0.003363086, 0.003306026, 
    0.003315752, 0.003428955, 0.003370589, 0.003343998, 0.003351593, 
    0.003406733, 0.002956327, 0.002791533, 0.003250284, 0.003041331, 
    0.002808413, 0.002729369, 0.003007144, 0.003066575, 0.003009001, 
    0.002897548, 0.002728926, 0.002743499, 0.00302121, 0.003027314, 
    0.003049806, 0.002919644, 0.002863679, 0.002843795, 0.002745487, 
    0.002731021, 0.00267075, 0.002657671, 0.002656145, 0.002673564, 
    0.002704812, 0.002763607, 0.002887106, 0.002928464, 0.003018428, 
    0.00308609, 0.003120581, 0.003173048, 0.00316879, 0.003259897, 
    0.003305515, 0.003317293, 0.003415251, 0.003410753, 0.003429094, 
    0.003452381, 0.003467735, 0.003458913, 0.003493739, 0.003392776, 
    0.003400849, 0.003317244, 0.003269227, 0.003097201, 0.002800213, 
    0.003243322, 0.003512209, 0.003340852, 0.002941356, 0.002426961, 
    0.001965749, 0.001740603, 0.001731524, 0.00249742, 0.002966769, 
    0.002926461, 0.002986303, 0.003007047, 0.003043905, 0.003040934, 
    0.003113095, 0.003097311, 0.003099838, 0.003067223, 0.00306212,
  0.002917498, 0.0031875, 0.003085788, 0.002175316, 0.0009505786, 
    0.0009483201, 0.001281869, 0.001259314, 0.00237257, 0.002849391, 
    0.002491747, 0.002843063, 0.003008878, 0.003314719, 0.003532855, 
    0.003597228, 0.003550449, 0.003462186, 0.003417078, 0.0033501, 
    0.00328625, 0.003216585, 0.003237486, 0.003327275, 0.003458884, 
    0.003419291, 0.003119519, 0.00251532, 0.003101921, 0.00314579, 
    0.002904814, 0.002693386, 0.002771587, 0.003119133, 0.002993427, 
    0.003014566, 0.002918802, 0.002925079, 0.003060501, 0.003125113, 
    0.003090907, 0.003131583, 0.003135111, 0.003168076, 0.003137305, 
    0.003130645, 0.003129421, 0.003097028, 0.003017426, 0.002983013, 
    0.002965609, 0.00292155, 0.00287571, 0.002857096, 0.002888855, 
    0.002882909, 0.002889188, 0.002929831, 0.002956996, 0.002980297, 
    0.003018586, 0.003100317, 0.003155025, 0.003208352, 0.003287982, 
    0.003376912, 0.003391346, 0.003441636, 0.00344472, 0.003477924, 
    0.003431082, 0.003415981, 0.003175369, 0.003077397, 0.002817869, 
    0.002623623, 0.003219655, 0.003809186, 0.003228873, 0.002350667, 
    0.002130414, 0.001570228, 0.001898481, 0.002734581, 0.002641996, 
    0.002657253, 0.002718369, 0.002873197, 0.002894307, 0.002948428, 
    0.003039615, 0.003027819, 0.003051091, 0.003168551, 0.003137732, 
    0.003133554,
  0.002435228, 0.002785858, 0.001158, 0.001301116, 0.00049771, 0.0008138688, 
    0.001186818, 0.001416337, 0.001989797, 0.00275493, 0.002590197, 
    0.002100407, 0.0025843, 0.002929594, 0.003368761, 0.003602171, 
    0.003729645, 0.003659217, 0.003597179, 0.003577169, 0.00354816, 
    0.003417015, 0.003273996, 0.003330534, 0.003406778, 0.003340339, 
    0.002807381, 0.002435304, 0.003044287, 0.002986655, 0.003018061, 
    0.003053222, 0.003239395, 0.003284296, 0.003079271, 0.003190503, 
    0.003252095, 0.003301432, 0.003354503, 0.003395701, 0.003353931, 
    0.003323732, 0.003322445, 0.003320266, 0.003314702, 0.00337828, 
    0.003397005, 0.00341665, 0.003382174, 0.003438901, 0.003478877, 
    0.003466224, 0.003502004, 0.003437772, 0.003337719, 0.003215918, 
    0.003128402, 0.00309108, 0.003005488, 0.002982283, 0.002927668, 
    0.002975559, 0.002998162, 0.002971807, 0.00304443, 0.00317971, 
    0.003272582, 0.003396193, 0.003460551, 0.003503688, 0.003340388, 
    0.003366612, 0.00333662, 0.003259024, 0.003300747, 0.002919374, 
    0.002905116, 0.003338323, 0.002611465, 0.001633408, 0.002042597, 
    0.002498644, 0.002710439, 0.002636099, 0.002588036, 0.002576608, 
    0.002689792, 0.002754452, 0.002803057, 0.002887188, 0.002921995, 
    0.0030447, 0.003168473, 0.003067797, 0.001964159, 0.002166258,
  0.001532017, 0.0013454, 0.001219943, 0.001407531, 0.001815004, 0.001896209, 
    0.001474367, 0.001905079, 0.002150286, 0.002459592, 0.002287168, 
    0.001876516, 0.002030199, 0.002216231, 0.002913462, 0.003278751, 
    0.00347748, 0.003690882, 0.003867054, 0.00412987, 0.003792206, 
    0.00346354, 0.003517691, 0.003390536, 0.00321296, 0.003026025, 0.0028018, 
    0.002872311, 0.002689123, 0.002724266, 0.00291721, 0.002952861, 
    0.002980549, 0.003030112, 0.00320344, 0.003277017, 0.003269562, 
    0.003272392, 0.003259817, 0.003247101, 0.003202805, 0.003183939, 
    0.003191391, 0.003219478, 0.003198974, 0.003230238, 0.003270848, 
    0.003330104, 0.003388453, 0.003408417, 0.00340155, 0.003449759, 
    0.003484312, 0.003503529, 0.003460536, 0.003395589, 0.00328045, 
    0.003173957, 0.003056604, 0.002925476, 0.002820905, 0.002769645, 
    0.002748154, 0.002774095, 0.002737269, 0.002836308, 0.003050342, 
    0.003243797, 0.003414409, 0.003520172, 0.00352467, 0.003493419, 
    0.00328695, 0.003110185, 0.00303353, 0.002727701, 0.002937208, 
    0.002892607, 0.002684103, 0.002691844, 0.002816917, 0.002744183, 
    0.002780089, 0.002686519, 0.002592819, 0.002592755, 0.002641696, 
    0.002632048, 0.002681639, 0.002701333, 0.002746997, 0.003028728, 
    0.002845082, 0.002291459, 0.00217295, 0.001858873,
  0.001789255, 0.001474668, 0.001509526, 0.001421645, 0.001134763, 
    0.00128023, 0.001322669, 0.001392511, 0.001819184, 0.00265759, 
    0.002501602, 0.001558546, 0.001266896, 0.00122716, 0.00244543, 
    0.002796541, 0.002997163, 0.00325432, 0.003575377, 0.003949787, 
    0.0035176, 0.00350172, 0.0036723, 0.003416017, 0.003054302, 0.002816759, 
    0.002267633, 0.002025481, 0.002143371, 0.002046254, 0.00260571, 
    0.002767198, 0.002728892, 0.002829807, 0.00298964, 0.003046831, 
    0.003071593, 0.003074439, 0.003079128, 0.003057351, 0.003038947, 
    0.003045257, 0.002988689, 0.002968965, 0.002946602, 0.002920836, 
    0.002874201, 0.002850153, 0.002907135, 0.002954802, 0.002983492, 
    0.003019001, 0.003018301, 0.00307476, 0.003104148, 0.003120933, 
    0.003078304, 0.00297955, 0.002862313, 0.002746839, 0.002613754, 
    0.002539032, 0.002513157, 0.002545152, 0.002509421, 0.002592804, 
    0.002644636, 0.002888395, 0.003284343, 0.003355805, 0.00343838, 
    0.003200231, 0.002923952, 0.002393836, 0.002955344, 0.003075426, 
    0.002920836, 0.002799784, 0.00269143, 0.002609874, 0.002601212, 
    0.00249731, 0.002469478, 0.002394519, 0.002381628, 0.002395028, 
    0.002407553, 0.002459209, 0.002475454, 0.002427787, 0.002519468, 
    0.002491109, 0.001942463, 0.001855678, 0.001880696, 0.001849687,
  0.0007034969, 0.0006766515, 0.0006054598, 0.0004452579, 0.0002637887, 
    0.0004874892, 0.0005294033, 0.000449724, 0.0006448459, 0.001686132, 
    0.002473739, 0.001962632, 0.000793254, 0.0005650874, 0.000980698, 
    0.002262325, 0.002604615, 0.002540147, 0.003068767, 0.003416047, 
    0.003225981, 0.003467706, 0.003698367, 0.003661253, 0.003374435, 
    0.002810274, 0.002352193, 0.00156433, 0.001320587, 0.00176996, 
    0.002289727, 0.002468573, 0.002383234, 0.002331164, 0.002522375, 
    0.002531387, 0.002596937, 0.002622241, 0.002626518, 0.002603406, 
    0.002568025, 0.002589656, 0.002635006, 0.002607871, 0.00255434, 
    0.002604965, 0.00263839, 0.002602563, 0.002618648, 0.00268148, 
    0.002710804, 0.002725588, 0.002719739, 0.002648483, 0.002616457, 
    0.002667032, 0.002665808, 0.002603614, 0.002460483, 0.002344674, 
    0.002162125, 0.00207995, 0.002024177, 0.002014989, 0.002045269, 
    0.002016166, 0.002012732, 0.002220554, 0.002243713, 0.002100345, 
    0.002236576, 0.00207124, 0.001895812, 0.002546202, 0.002879748, 
    0.002879636, 0.002821082, 0.002688172, 0.002668144, 0.002566085, 
    0.002413974, 0.002266984, 0.002110851, 0.002029152, 0.002018597, 
    0.002039992, 0.002087675, 0.00207477, 0.002112693, 0.002082208, 
    0.00218131, 0.002304351, 0.001576108, 0.001081518, 0.0006804499, 
    0.0006289515,
  0.0003055916, 0.000361922, 0.0003288293, 0.0004329069, -2.081867e-005, 
    0.000199829, 0.0002935757, 0.000353212, 0.0003344559, 0.0009524375, 
    0.001921896, 0.0009517549, 0.0005576159, 0.0004310159, 0.0001733811, 
    0.0009497683, 0.002441362, 0.002450788, 0.002659737, 0.002683022, 
    0.002683722, 0.002348569, 0.002917244, 0.00345418, 0.00309633, 
    0.002879623, 0.002234604, 0.002212449, 0.001278992, 0.001125657, 
    0.001751346, 0.002000176, 0.001976619, 0.001842994, 0.001813239, 
    0.001885369, 0.001970931, 0.002043838, 0.002067122, 0.002059398, 
    0.002080665, 0.002092299, 0.002147613, 0.002152715, 0.002100899, 
    0.002155337, 0.002179847, 0.002143196, 0.002148409, 0.002178768, 
    0.002186873, 0.002232395, 0.002326047, 0.002295226, 0.002271066, 
    0.002262786, 0.002249021, 0.002279744, 0.002221746, 0.002100026, 
    0.001906, 0.001704839, 0.001497431, 0.001472205, 0.001518251, 
    0.001583086, 0.001568716, 0.001386057, 0.0007974962, 0.0002098596, 
    0.001101098, 0.001502484, 0.001581226, 0.002234287, 0.002506164, 
    0.002625262, 0.002684562, 0.002645589, 0.00255836, 0.002416344, 
    0.002296975, 0.00217144, 0.002023492, 0.001872495, 0.001761377, 
    0.001799761, 0.001816037, 0.001758149, 0.001767782, 0.001713452, 
    0.001777556, 0.001843869, 0.0009309328, 0.0004843741, -3.90975e-005, 
    2.530729e-005,
  0.0005424686, 0.0003707435, 0.0001235195, 4.886277e-005, 9.201677e-005, 
    0.0002031352, 6.704638e-005, 8.759787e-005, 0.0001988444, 0.000615791, 
    0.001275097, 0.0003621918, 0.0004033591, 0.0005230457, 0.0001913894, 
    0.0003917716, 0.00196152, 0.001993898, 0.001435585, 0.001255389, 
    0.00140669, 0.001397598, 0.001770436, 0.001582641, 0.002430075, 
    0.002360092, 0.001857221, 0.002124725, 0.001142664, 0.0006346893, 
    0.000852921, 0.001168158, 0.001555081, 0.001572978, 0.00154796, 
    0.001570497, 0.001549135, 0.001618006, 0.001651956, 0.001655787, 
    0.001710339, 0.001763538, 0.001714439, 0.001666214, 0.00168095, 
    0.001709066, 0.0017355, 0.001763283, 0.001777462, 0.001806516, 
    0.001850385, 0.001889375, 0.001922849, 0.001923373, 0.001905556, 
    0.001945705, 0.002013193, 0.002031329, 0.002017659, 0.001945451, 
    0.001828768, 0.001679423, 0.001489785, 0.001396611, 0.001373771, 
    0.001425937, 0.001257152, 0.0002389615, 0.0003067218, 0.0009516426, 
    0.00130315, 0.001746942, 0.001579891, 0.001696907, 0.00200779, 
    0.002208903, 0.002279921, 0.002368437, 0.002453855, 0.002375351, 
    0.002255679, 0.002177559, 0.0020882, 0.00190031, 0.001824143, 
    0.001792942, 0.001749249, 0.001734497, 0.001674782, 0.001634536, 
    0.001667741, 0.001552108, 0.0007329336, 0.0006123255, 0.0006336085, 
    0.0003963024,
  0.0002854692, 0.0005244124, 0.0004572736, 0.0002862955, 0.0006679408, 
    0.0006671781, 0.0001342641, 0.0003220267, 0.0007511959, 0.0003016975, 
    0.0001605055, 0.0001681678, 0.0003225196, 0.0002660779, 0.0005221716, 
    0.0003349497, 0.0002286793, 0.0003368575, 0.0003035581, 0.0005030031, 
    0.001270871, 0.001240368, 0.001127373, 0.0008890019, 0.0009837493, 
    0.001527074, 0.001277959, 0.001436968, 0.001029701, 0.000933348, 
    0.001004588, 0.0009129078, 0.00112197, 0.00130029, 0.001358305, 
    0.001356176, 0.001367874, 0.001456947, 0.001441101, 0.001396706, 
    0.001350072, 0.001385247, 0.001375042, 0.00135651, 0.001342904, 
    0.001278133, 0.00127481, 0.001290927, 0.001279293, 0.001245564, 
    0.001303881, 0.001374914, 0.001419007, 0.001493965, 0.00156193, 
    0.001662336, 0.001712197, 0.001663163, 0.001700102, 0.001725915, 
    0.00165226, 0.001535371, 0.001394735, 0.001366315, 0.001291309, 
    0.001185483, 0.0003551841, 0.0001737475, 0.00034614, 0.0008640806, 
    0.001130742, 0.001561199, 0.001574089, 0.001548833, 0.001208627, 
    0.001730174, 0.00190581, 0.001914917, 0.001977462, 0.002032171, 
    0.002032839, 0.002073466, 0.002052691, 0.001923008, 0.001838306, 
    0.001739283, 0.001734164, 0.001771182, 0.001679105, 0.001590795, 
    0.001523434, 0.001480407, 0.00136851, 0.0005030832, 0.0002721336, 
    6.308872e-005,
  5.851965e-006, 7.937988e-005, 2.332008e-005, 0.0006184457, 0.0008933269, 
    0.00120764, 0.0002536494, 0.0003901678, 0.001289942, 0.000218173, 
    -4.813541e-006, 0.0002006555, 0.0003144129, 0.0004466402, 0.0005952385, 
    0.0005258112, 0.0004598969, 0.0007017483, 0.0006817691, 0.0001188302, 
    -0.0004370974, 0.0006356908, 0.0005265744, 0.0005153051, 0.0005694103, 
    0.0006795913, 0.0007132085, 0.0009689038, 0.0009652961, 0.0008779874, 
    0.0009950188, 0.001002871, 0.001080086, 0.0006267908, 0.0008836454, 
    0.001149116, 0.001234836, 0.001300258, 0.001314198, 0.001335353, 
    0.001264527, 0.001185516, 0.001120682, 0.001069659, 0.001066862, 
    0.001045262, 0.001030177, 0.001024867, 0.001021372, 0.001004047, 
    0.0009681396, 0.0009631813, 0.0010273, 0.001147049, 0.001301737, 
    0.001435999, 0.001456009, 0.001369718, 0.001374884, 0.001393416, 
    0.0013759, 0.001282646, 0.001211248, 0.001224504, 0.00113071, 
    0.0008729496, 0.0005248422, 0.00042922, 0.000564801, 0.0007169121, 
    0.0008371072, 0.001089259, 0.0009664265, 0.0008739037, 0.0008828514, 
    0.001339312, 0.001592431, 0.001625381, 0.001655756, 0.001641308, 
    0.001661065, 0.001698688, 0.001709766, 0.001717523, 0.001659492, 
    0.001586583, 0.001583452, 0.001532892, 0.001511036, 0.001536213, 
    0.001452656, 0.001438859, 0.001414843, 0.00118445, 0.0002241493, 
    2.610264e-005,
  0.0002326523, 0.0003863215, 0.0004216395, 0.001297921, 0.00140389, 
    0.00130652, 0.001110126, 0.001041764, 0.001221659, 0.001211566, 
    0.0005011121, 0.0002589095, 0.0006524909, 0.0008994604, 0.0009209509, 
    0.0008097989, 0.0009406274, 0.001052796, 0.0009891537, 0.0006642693, 
    0.0005131433, 0.0005651661, 0.0005112202, 0.0004421108, 0.0004490248, 
    0.0004802577, 0.0004955801, 0.0006019145, 0.0006948025, 0.0005956045, 
    0.0005361589, 0.0006804657, 0.0009784093, 0.0005786291, 0.001013154, 
    0.001080692, 0.000846229, 0.0008207189, 0.001118901, 0.001206337, 
    0.001204144, 0.00117051, 0.001140613, 0.001078655, 0.001040747, 
    0.001015951, 0.0009909654, 0.0009610835, 0.000950784, 0.0009458247, 
    0.0008921963, 0.0008520945, 0.0008339109, 0.0008836137, 0.0009901864, 
    0.001149625, 0.001232817, 0.001214379, 0.001186739, 0.001217987, 
    0.00120702, 0.00113071, 0.001081628, 0.001041955, 0.0008296845, 
    0.000746937, 0.0007672976, 0.0007300084, 0.0006454494, 0.0004676846, 
    0.000728738, 0.0008889232, 0.0009470498, 0.0009908075, 0.0009768037, 
    0.001027731, 0.001292358, 0.00136533, 0.001470218, 0.001498734, 
    0.0015262, 0.001464989, 0.001343539, 0.001350263, 0.001329123, 
    0.00130002, 0.001301387, 0.001235679, 0.001242275, 0.001319841, 
    0.001329774, 0.001257056, 0.001193955, 0.001251143, 0.001136924, 
    0.0004828973,
  0.0008443235, 0.001213283, 0.0012716, 0.001297762, 0.001267801, 
    0.001140709, 0.0009059464, 0.0008026627, 0.0007640871, 0.0007424224, 
    0.0007871022, 0.0008733144, 0.0008532072, 0.0009562999, 0.0009822724, 
    0.0009417878, 0.0009764379, 0.0009515791, 0.0009492105, 0.000584685, 
    0.0003891498, 0.0005514496, 0.0005175146, 0.0004515045, 0.000546999, 
    0.0005013339, 0.0005367948, 0.0003890547, 0.0003346951, 0.0003933777, 
    0.0003637343, 0.0004012616, 0.0005111406, 0.000406602, 0.0004048379, 
    0.0008409219, 0.0008949949, 0.0007666296, 0.0009034984, 0.0009896476, 
    0.001059568, 0.001061904, 0.001073396, 0.001090594, 0.001069009, 
    0.001008849, 0.0009669825, 0.0009248937, 0.000879372, 0.0008516195, 
    0.0008424162, 0.0008321642, 0.0007947795, 0.0008182717, 0.0009009391, 
    0.0009940495, 0.001071297, 0.001102149, 0.001109746, 0.001133382, 
    0.00116525, 0.001088829, 0.001014506, 0.0009091734, 0.0008835183, 
    0.0009313927, 0.0009140046, 0.0007406585, 0.0005898345, 0.0007032258, 
    0.0008133757, 0.0008519038, 0.0009810156, 0.0009565218, 0.0009287545, 
    0.001043974, 0.001196579, 0.001435442, 0.001476401, 0.001532032, 
    0.001521891, 0.001398343, 0.001140295, 0.0007944442, 0.0006412044, 
    0.0007387977, 0.0008109594, 0.0007641967, 0.0006830078, 0.0007940782, 
    0.001020323, 0.001037647, 0.0009624977, 0.001010706, 0.0008288738, 
    0.0006592316,
  0.0009780284, 0.001227811, 0.001259044, 0.001165966, 0.001227954, 
    0.001071361, 0.001039015, 0.0009601461, 0.0008312571, 0.0007340773, 
    0.0007348566, 0.0007363509, 0.0007979742, 0.0007465868, 0.0008382506, 
    0.0008820083, 0.0007973542, 0.001162007, 0.001121857, 0.0005920281, 
    0.0005008254, 0.0006940876, 0.0007129861, 0.0005776755, 0.0004145495, 
    0.0002752652, 0.0003236323, 0.0002728492, 0.0003190866, 0.0003610165, 
    0.0003215344, 0.0003495406, 0.0003335665, 0.0002763459, 0.000252218, 
    0.0002630422, 0.0006527926, 0.0007958286, 0.000662457, 0.0008758409, 
    0.0009594786, 0.0008621241, 0.0006944521, 0.0006558122, 0.0006487712, 
    0.0006623617, 0.0006872364, 0.0007026228, 0.0007321709, 0.000731424, 
    0.0007107607, 0.0007132404, 0.0007377025, 0.0007864833, 0.0008506021, 
    0.0009018779, 0.0009583198, 0.001004525, 0.001007163, 0.0009985953, 
    0.00101759, 0.0009801895, 0.000952072, 0.0008714553, 0.0009527553, 
    0.0007451882, 0.0005175145, 0.0004511389, 0.0004487548, 0.0006329883, 
    0.0008369633, 0.0007342368, 0.000793762, 0.0009277212, 0.0009338879, 
    0.0008533349, 0.000895837, 0.001005461, 0.001386089, 0.001492774, 
    0.001204288, 0.0008423841, 0.0007169759, 0.0005675191, 0.0004567346, 
    0.0002961676, 0.0002529491, 0.0003815521, 0.000452077, 0.0005934271, 
    0.0007278472, 0.0008380278, 0.0008579125, 0.0008881595, 0.0007412154, 
    0.0008442118,
  0.00102533, 0.001004318, 0.001082836, 0.001054035, 0.0009814447, 
    0.001005589, 0.000902592, 0.0009078211, 0.001023009, 0.0009433455, 
    0.0007871496, 0.0006917825, 0.0006481358, 0.0006330041, 0.000707549, 
    0.0006453702, 0.0005381458, 0.0005481272, 0.0005452823, 0.0005441222, 
    0.0005664539, 0.0005232525, 0.0003889113, 0.0003618748, 0.0003649584, 
    0.0002854377, 0.000262025, 0.000278603, 0.000288569, 0.00028779, 
    0.0002896657, 0.0002672542, 0.0002424587, 0.0002179811, 0.0002021501, 
    0.0001488239, 0.0001614441, 0.000570538, 0.0006147095, 0.0005423573, 
    0.0005682018, 0.0005449483, 0.0005599207, 0.0005535786, 0.000524285, 
    0.0005355859, 0.0005730337, 0.0005805839, 0.0005902953, 0.0005949368, 
    0.00060743, 0.0006501228, 0.0007091393, 0.0007611313, 0.0007884698, 
    0.0008048886, 0.0008317665, 0.0008792439, 0.0009143231, 0.000914562, 
    0.0009319982, 0.0009015445, 0.000902927, 0.0008382667, 0.0008291269, 
    0.000543518, 0.0004805119, 0.0005171648, 0.0005416584, 0.0005370013, 
    0.0004714363, 0.0005429141, 0.0006352296, 0.001121969, 0.0007205518, 
    0.0006131043, 0.0005822846, 0.000622959, 0.0007064691, 0.0009192972, 
    0.0008421764, 0.0007303266, 0.0006049662, 0.0004944031, 0.0004187454, 
    0.0003714599, 0.000202199, 5.517388e-005, 7.792376e-006, 0.0001868922, 
    0.0003917576, 0.0005680746, 0.0007245094, 0.0008226107, 0.0009271177, 
    0.0009237961,
  0.0009385776, 0.0009796964, 0.0009979911, 0.001010134, 0.0009813653, 
    0.0009235251, 0.0008416998, 0.0007577608, 0.0007241119, 0.0006924658, 
    0.0006465943, 0.000688127, 0.0006411903, 0.0005381139, 0.0004765067, 
    0.0004826895, 0.0004772692, 0.0004398692, 0.0003635914, 0.0003421179, 
    0.0004202713, 0.0004036933, 0.0003369521, 0.0003075629, 0.0002657443, 
    0.0002254675, 0.0002326042, 0.0002560009, 0.0002413144, 0.0002205083, 
    0.0002205878, 0.0001966187, 0.0001636535, 0.0001535922, 0.0001541962, 
    0.0001328657, 0.0001178613, 0.0001927565, 0.0005787403, 0.001091547, 
    0.0008431782, 0.0006523319, 0.0005772777, 0.0005638783, 0.0005650388, 
    0.0005441532, 0.0005715713, 0.0005958583, 0.0006030586, 0.0006247386, 
    0.0006430494, 0.0006669392, 0.0006814669, 0.0007010652, 0.0007318687, 
    0.000796766, 0.0008295253, 0.0008305265, 0.0008613463, 0.0008820407, 
    0.0008782577, 0.0008638892, 0.0007630694, 0.0006087015, 0.0004932752, 
    0.0004587523, 0.0005110933, 0.0004942768, 0.0003918682, 0.0004697673, 
    0.0004256915, 0.0004095427, 0.0004118474, 0.0004544448, 0.0004806709, 
    0.0005143991, 0.0005504003, 0.0005199939, 0.0004627577, 0.000544869, 
    0.0008729964, 0.0007929356, 0.0007725905, 0.0005937761, 0.0004797962, 
    0.0003399397, 0.0001350283, -0.0001357836, -0.0003028354, -0.0002012528, 
    7.933378e-005, 0.0003644349, 0.0005642138, 0.0006847898, 0.0007813657, 
    0.0008580564,
  0.0008346427, 0.0007686494, 0.0008418744, 0.0008360888, 0.0007486374, 
    0.0007138283, 0.0006606132, 0.0006172053, 0.0005649123, 0.0005558681, 
    0.0005293242, 0.0004770787, 0.0004292519, 0.000420796, 0.0004292678, 
    0.0004030417, 0.0003642114, 0.0003579966, 0.0003646087, 0.0003450584, 
    0.0003204853, 0.0003383666, 0.0003204216, 0.000274534, 0.0002200791, 
    0.000208953, 0.0002325565, 0.0002175996, 0.0001817414, 0.0001678656, 
    0.000169916, 0.0001467894, 0.0001314035, 0.0001277636, 0.0001192282, 
    9.060215e-005, 8.325881e-005, 0.0001615714, 0.0004987746, 0.001241926, 
    0.00114295, 0.0009171994, 0.0005359362, 0.0005532929, 0.0006181109, 
    0.0005807106, 0.0005713168, 0.0005789781, 0.0006052204, 0.0006496457, 
    0.0007192956, 0.0007892002, 0.0008324177, 0.0008412071, 0.0008410171, 
    0.0009090614, 0.0008978243, 0.0008513001, 0.0008771615, 0.000919282, 
    0.000887048, 0.000932696, 0.000726687, 0.0005442967, 0.0004642042, 
    0.0004662389, 0.0004996649, 0.0004941016, 0.0004943878, 0.0004784616, 
    0.0004258664, 0.0003504306, 0.000362415, 0.0004278689, 0.0005105048, 
    0.000816841, 0.000575482, 0.000472628, 0.0003674059, 0.000414756, 
    0.0005930137, 0.001130044, 0.001036679, 0.0005534037, 0.0003356319, 
    0.0003162569, 0.0002378493, 4.819501e-005, -0.0001447643, -0.0001539513, 
    3.738794e-005, 0.0003126664, 0.0005334732, 0.00063984, 0.0006907969, 
    0.0007246521,
  0.0005673757, 0.0006239759, 0.0005878636, 0.000684741, 0.0006625522, 
    0.0006442096, 0.0005712218, 0.0004082236, 0.0003566613, 0.0003898811, 
    0.0004193498, 0.0003925513, 0.0003544204, 0.0003639254, 0.0003864956, 
    0.0003435166, 0.000287361, 0.0002865663, 0.0003065935, 0.0003118226, 
    0.0002935121, 0.0002886484, 0.0002884894, 0.0002794136, 0.0002720703, 
    0.0002730716, 0.0002443025, 0.0001825361, 0.0001425614, 0.0001409084, 
    0.0001282087, 0.0001053046, 9.35267e-005, 9.649896e-005, 8.666021e-005, 
    7.074977e-005, 8.866291e-005, 0.0001746526, 0.0004921943, 0.000851952, 
    0.0008938342, 0.0008708669, 0.0004190792, 0.0004234186, 0.0007583968, 
    0.0006229589, 0.0007092662, 0.0008587225, 0.0009030844, 0.001018098, 
    0.001097237, 0.001097109, 0.0009723529, 0.0009502277, 0.0009023531, 
    0.0008885732, 0.0009172312, 0.0009019885, 0.0009407713, 0.0009181532, 
    0.0009088547, 0.0006908606, 0.0005555981, 0.0005074214, 0.0005236338, 
    0.0005343943, 0.0004885704, 0.0004001966, 0.0003438504, 0.0003294338, 
    0.0003292271, 0.0003466318, 0.0004455596, 0.0005226959, 0.0006021529, 
    0.0006351183, 0.0004293631, 0.0003555963, 0.0003213435, 0.0003902306, 
    0.0007157357, 0.001208992, 0.0008736961, 0.0003269706, 0.000175447, 
    0.0003420059, 0.0004242125, 0.0003305939, 0.0002096687, 0.0001986218, 
    0.0002869004, 0.0004115934, 0.0005156873, 0.0005963519, 0.000615505, 
    0.0006106563,
  0.000452871, 0.0004561772, 0.0004680504, 0.0004174263, 0.0004522356, 
    0.0008239935, 0.0004821809, 0.0003732076, 0.0002715142, 0.0002500884, 
    0.0002834033, 0.0003054174, 0.0002960871, 0.0002806377, 0.0002765685, 
    0.0002785235, 0.0002783805, 0.0002660939, 0.0002379923, 0.000214675, 
    0.0002106219, 0.0002371659, 0.0002425222, 0.0002239893, 0.000197207, 
    0.0001792143, 0.0001677226, 0.0001487445, 0.0001321982, 0.0001243781, 
    0.0001118849, 8.993447e-005, 7.553402e-005, 7.295911e-005, 7.35154e-005, 
    7.394457e-005, 8.419658e-005, 0.0001055112, 0.0001281292, 0.0001492371, 
    0.0001719346, 0.0002028336, 0.0002169639, 0.0002244503, 0.000253585, 
    0.0003526558, 0.0005064835, 0.001310256, 0.00142786, 0.001416257, 
    0.001356748, 0.001235138, 0.0006769688, 0.000628554, 0.0006388697, 
    0.0006848366, 0.0007270846, 0.0007257017, 0.0006882697, 0.0006494552, 
    0.0005771986, 0.0004986317, 0.0004509321, 0.0004433663, 0.0004401238, 
    0.0004181732, 0.0003685186, 0.0003148744, 0.000279954, 0.0002619774, 
    0.0002625655, 0.0003155262, 0.0003376515, 0.0003513526, 0.00035415, 
    0.0003613026, 0.0002921771, 0.0002677788, 0.0003053218, 0.0003697743, 
    0.0004919876, 0.0006220373, 0.0003818703, 0.0001853182, 0.0001914692, 
    0.0002796841, 0.0002787134, 0.000304447, 0.0003360454, 0.0004104329, 
    0.0004395195, 0.0003789142, 0.0002268506, 0.0002147867, 0.000374909, 
    0.0004378194,
  0.0001836163, 0.0002474166, 0.0002454463, 0.0004330664, 0.0004408552, 
    0.000442063, 0.0005716672, 0.0003342183, 0.0002700518, 0.0002409966, 
    0.0002539665, 0.0002898246, 0.0002971202, 0.0002826561, 0.0002579559, 
    0.0002429197, 0.0002428402, 0.0002441118, 0.0002338756, 0.0002198249, 
    0.0002069027, 0.0002020072, 0.0001922956, 0.0001747797, 0.0001625091, 
    0.000156199, 0.0001506199, 0.0001354248, 0.0001124889, 9.139678e-005, 
    8.591314e-005, 8.327464e-005, 7.742547e-005, 7.329286e-005, 
    7.184647e-005, 7.829964e-005, 9.428959e-005, 9.525915e-005, 
    9.886723e-005, 9.603798e-005, 0.0001024276, 0.0001272709, 0.0001401932, 
    0.0001479656, 0.00016359, 0.0001886398, 0.0002142141, 0.000244382, 
    0.0002792707, 0.0003019362, 0.0003364275, 0.0004672875, 0.0003947764, 
    0.000400276, 0.0004043769, 0.0004204623, 0.0004380575, 0.0004388998, 
    0.00042771, 0.0004065225, 0.0003966361, 0.000390771, 0.0003863683, 
    0.000363337, 0.0003088663, 0.0002515028, 0.0002073477, 0.0001841735, 
    0.0001758606, 0.0001695981, 0.0001632879, 0.0001596799, 0.000163876, 
    0.0001756539, 0.0002251496, 0.00023173, 0.000236101, 0.0001825998, 
    0.000173381, 0.0001976838, 0.0002744386, 0.0003093113, 0.0002010216, 
    0.0001430064, 0.0001196573, 0.0001170188, 0.0001162241, 0.0001689943, 
    0.0001982399, 0.000394363, 0.0006498203, 0.0005640539, 0.0005251272, 
    0.0002437297, 8.061971e-005, 0.0001077517,
  0.0001534962, 0.0001165573, 0.0001033335, 7.054233e-005, -8.194987e-005, 
    0.0001563899, 0.0001451204, 0.0001536558, 0.000202945, 0.0002885848, 
    0.0003840954, 0.0008053336, 0.000728054, 0.0005573622, 0.0003325332, 
    0.0002667616, 0.0002190462, 0.0001946162, 0.0001856675, 0.0001812806, 
    0.0001740168, 0.000165084, 0.0001556744, 0.0001493007, 0.0001410673, 
    0.0001387785, 0.0001207858, 0.0001004249, 8.799536e-005, 7.950765e-005, 
    7.661482e-005, 7.216434e-005, 6.415347e-005, 5.377432e-005, 
    5.523662e-005, 5.940099e-005, 6.885827e-005, 8.292496e-005, 
    8.314748e-005, 8.389453e-005, 8.78205e-005, 9.83268e-005, 0.0001147618, 
    0.0001262218, 0.0001387944, 0.0001422753, 0.0001500001, 0.0001600931, 
    0.0001792938, 0.0002224952, 0.0002732625, 0.0003286391, 0.0003839045, 
    0.0002854377, 0.0002601494, 0.0002397726, 0.0002366891, 0.0002463372, 
    0.0002524088, 0.0002475451, 0.0002398362, 0.0002292823, 0.0002133082, 
    0.0001890848, 0.0001668165, 0.0001516054, 0.0001444688, 0.0001407336, 
    0.0001427204, 0.0001767665, 0.0001505564, 0.0001495551, 0.0001464874, 
    0.0001692325, 0.0001469007, 0.0001755903, 0.0001505087, 0.0001540691, 
    0.0001606812, 0.0001907856, 0.0001778791, 0.0001555948, 9.544988e-005, 
    6.801594e-005, 5.077029e-005, 4.169445e-005, 3.894472e-005, 
    5.166035e-005, 8.869471e-005, 0.0001533855, 0.0002921133, 0.000463759, 
    0.0008135666, 0.0009645016, 0.0005743534, 0.0003065132,
  0.0005215672, 0.0003313567, 0.0002049468, 0.0001347882, 5.820813e-005, 
    9.901007e-005, 0.0002748361, 0.0004838021, 0.000772511, 0.0009979437, 
    0.001130314, 0.001146606, 0.0009846877, 0.0006482473, 0.0004847397, 
    0.0003078332, 0.0002954513, 0.0002533625, 0.0002350996, 0.0001963327, 
    0.000186351, 0.000176846, 0.0001680563, 0.0001558811, 0.0001409084, 
    0.0001249661, 0.0001099457, 9.799301e-005, 9.077688e-005, 8.851985e-005, 
    8.635819e-005, 8.726418e-005, 8.68827e-005, 8.527735e-005, 8.454621e-005, 
    0.0001009812, 9.808839e-005, 9.668966e-005, 8.28137e-005, 7.758439e-005, 
    8.540451e-005, 8.893311e-005, 9.991628e-005, 0.0001149367, 0.0001268894, 
    0.0001330088, 0.000137507, 0.0001441668, 0.0001562625, 0.0001703133, 
    0.0001823456, 0.0001850635, 0.0001756698, 0.000157995, 0.0001463761, 
    0.0001435151, 0.0001513193, 0.0001669119, 0.0001839509, 0.0001978745, 
    0.0002059649, 0.0002098431, 0.0002143254, 0.0001518279, 0.0001364421, 
    0.0001234085, 0.0001139353, 0.000111726, 0.0001155725, 0.0001529724, 
    0.0001317372, 0.0001334379, 0.000153481, 0.0001204044, 0.0001141419, 
    0.0001122187, 0.0001171142, 0.0001465509, 0.0001491259, 0.0001440715, 
    0.0001419098, 0.0001006951, 8.880603e-005, 8.411711e-005, 8.257529e-005, 
    7.059083e-005, 4.876756e-005, 3.191932e-005, 4.207595e-005, 7.81884e-005, 
    0.0001336287, 0.0002362916, 0.0003549765, 0.0005126188, 0.0007075341, 
    0.0008608688,
  0.0006382019, 0.0006297461, 0.000450789, 0.0004270901, 0.000623547, 
    0.0008769386, 0.0009365749, 0.000803728, 0.0007161808, 0.0006211151, 
    0.0005350142, 0.0004678439, 0.0004262478, 0.0003730486, 0.0003258099, 
    0.0002918751, 0.0002645363, 0.0002463848, 0.0002371182, 0.0002321432, 
    0.0002320637, 0.0002245774, 0.0002144049, 0.0002035012, 0.000196444, 
    0.0001501113, 0.0001354565, 0.0001187672, 0.0001080543, 0.0001008699, 
    9.59903e-005, 0.000113522, 0.0001046528, 0.0001025548, 0.000101617, 
    0.0001035243, 0.0001062582, 0.0001081338, 0.0001094212, 0.0001103431, 
    0.0001120756, 0.0001142055, 0.0001163831, 0.000117909, 0.0001173686, 
    0.0001148254, 0.0001116147, 0.0001093895, 0.000108706, 0.000111424, 
    0.0001166056, 0.0001228204, 0.0001281133, 0.0001319121, 0.0001335016, 
    0.0001328499, 0.0001300524, 0.000124998, 0.0001194507, 0.000115938, 
    0.0001142373, 0.0001151592, 0.0001182428, 0.0001237264, 0.0001362354, 
    0.0001043032, 0.0001017441, 9.943942e-005, 9.750028e-005, 9.726187e-005, 
    9.740492e-005, 9.810428e-005, 0.0001008223, 0.0001033972, 0.0001059085, 
    0.0001234403, 0.0001214217, 0.0001194507, 8.604032e-005, 7.284783e-005, 
    6.335876e-005, 5.547507e-005, 5.173981e-005, 5.339284e-005, 
    5.887648e-005, 5.922615e-005, 5.657176e-005, 5.674659e-005, 
    6.587012e-005, 9.001397e-005, 0.0001283517, 0.0001772593, 0.0002566686, 
    0.0003273357, 0.0004067928, 0.0005076597,
  0.0003076424, 0.0003225674, 0.0003368567, 0.0003868132, 0.0002726426, 
    0.0002618184, 0.0002496432, 0.000279366, 0.0002629946, 0.0002499134, 
    0.0002414733, 0.0002382308, 0.000238358, 0.0002394229, 0.0002415687, 
    0.0002417594, 0.0002391686, 0.0002334147, 0.0002244661, 0.0002126247, 
    0.0001987646, 0.0001845549, 0.0001724114, 0.000164035, 0.0001643688, 
    0.0001305133, 0.000126794, 0.00015755, 0.0001437536, 0.0001377612, 
    0.0001325955, 0.0001267463, 0.0001202136, 0.0001131246, 0.0001058767, 
    9.934406e-005, 9.319285e-005, 8.788407e-005, 8.451442e-005, 
    8.327464e-005, 8.348127e-005, 8.530915e-005, 8.877417e-005, 
    9.319285e-005, 9.823143e-005, 0.0001034449, 0.0001082927, 0.0001124889, 
    0.0001161764, 0.0001186719, 0.000119403, 0.0001180043, 0.0001138558, 
    0.0001070529, 9.856524e-005, 8.901259e-005, 8.046131e-005, 7.451673e-005, 
    7.106761e-005, 7.08133e-005, 7.375379e-005, 7.898311e-005, 8.63264e-005, 
    9.463926e-005, 0.0001015693, 0.0001051138, 0.0001051297, 0.0001017441, 
    9.62764e-005, 9.112656e-005, 9.39399e-005, 6.332695e-005, 6.280242e-005, 
    6.114938e-005, 6.396273e-005, 6.847679e-005, 7.229149e-005, 7.40558e-005, 
    7.467566e-005, 7.125836e-005, 6.428063e-005, 5.601544e-005, 4.79728e-005, 
    4.177392e-005, 3.830891e-005, 3.743471e-005, 4.115404e-005, 
    4.938742e-005, 6.191235e-005, 7.885595e-005, 0.000102062, 0.0001298617, 
    0.0001813283, 0.0002165506, 0.0002523452, 0.0002831967,
  0.0001765281, 0.0001819164, 0.0001863668, 0.0001894504, 0.0001876543, 
    0.0001882742, 0.0001898636, 0.0001884967, 0.000187241, 0.0001873364, 
    0.0001879563, 0.0001887828, 0.0001889894, 0.0001887351, 0.0001868119, 
    0.0001836171, 0.0001790077, 0.0001729678, 0.0001658629, 0.0001580428, 
    0.0001500637, 0.0001429111, 0.0001363625, 0.000131467, 0.0001283675, 
    0.0001258085, 0.0001249025, 0.0001256973, 0.0001260151, 0.0001264443, 
    0.0001268735, 0.0001270483, 0.0001261582, 0.0001246164, 0.000121819, 
    0.0001183222, 0.0001145552, 0.0001110901, 0.0001078, 0.000105082, 
    0.0001031429, 0.0001019508, 0.000101156, 0.0001006951, 0.0001006633, 
    0.0001010925, 0.0001016488, 0.0001013309, 0.0001007587, 9.970964e-005, 
    9.799301e-005, 9.562472e-005, 9.281139e-005, 8.998215e-005, 
    8.723239e-005, 8.503893e-005, 8.392632e-005, 8.414885e-005, 
    8.529325e-005, 8.783638e-005, 9.147624e-005, 9.521146e-005, 
    9.856522e-005, 0.000101013, 0.0001020938, 0.000101617, 9.940763e-005, 
    9.591083e-005, 9.171467e-005, 8.734365e-005, 8.341769e-005, 
    8.001626e-005, 7.890363e-005, 7.87129e-005, 8.022288e-005, 8.306801e-005, 
    8.540452e-005, 8.747081e-005, 9.036363e-005, 9.448031e-005, 
    9.565651e-005, 9.699166e-005, 9.632408e-005, 9.557704e-005, 
    9.508431e-005, 9.614925e-005, 9.810428e-005, 0.0001019826, 0.0001067668, 
    0.0001136174, 0.0001215965, 0.0001324843, 0.0001398911, 0.0001496504, 
    0.0001601408, 0.000169455,
  0.0001314511, 0.0001349956, 0.000135838, 0.0001378566, 0.000139605, 
    0.0001413534, 0.0001424502, 0.0001433085, 0.0001440714, 0.0001443098, 
    0.0001442463, 0.0001440078, 0.0001438012, 0.0001431495, 0.0001417031, 
    0.0001401931, 0.0001386037, 0.0001367122, 0.0001347095, 0.0001326273, 
    0.0001307358, 0.0001288285, 0.0001271437, 0.0001258721, 0.0001245211, 
    0.0001233926, 0.0001224548, 0.0001211514, 0.0001199911, 0.0001194507, 
    0.0001182586, 0.0001174639, 0.0001171142, 0.0001168122, 0.0001165102, 
    0.0001159221, 0.0001153181, 0.0001146982, 0.0001138717, 0.0001129498, 
    0.0001118372, 0.0001107564, 0.000109612, 0.0001084199, 0.0001072754, 
    0.0001061787, 0.0001049072, 0.0001036197, 0.0001024912, 0.0001013944, 
    0.00010025, 9.924868e-005, 9.824734e-005, 9.751617e-005, 9.638766e-005, 
    9.522736e-005, 9.4226e-005, 9.320875e-005, 9.230276e-005, 9.171465e-005, 
    9.119014e-005, 9.037951e-005, 8.952121e-005, 8.875827e-005, 
    8.810659e-005, 8.759797e-005, 8.708934e-005, 8.677145e-005, 8.63423e-005, 
    8.578598e-005, 8.54363e-005, 8.545219e-005, 8.530914e-005, 8.577009e-005, 
    8.615157e-005, 8.667608e-005, 8.734366e-005, 8.831322e-005, 8.95371e-005, 
    9.098351e-005, 9.266833e-005, 9.451211e-005, 9.648304e-005, 9.86288e-005, 
    0.0001008699, 0.0001032223, 0.0001055588, 0.0001079112, 0.0001103908, 
    0.0001128385, 0.0001157949, 0.0001185447, 0.0001207064, 0.0001233607, 
    0.0001257767, 0.0001286377,
  2.284739e-005, 2.084467e-005, 1.911216e-005, 1.74909e-005, 1.602861e-005, 
    1.472525e-005, 1.348547e-005, 1.243642e-005, 1.148274e-005, 
    1.079928e-005, 1.02112e-005, 9.734355e-006, 9.352883e-006, 9.130363e-006, 
    8.987307e-006, 8.907831e-006, 8.971416e-006, 9.209838e-006, 
    9.432362e-006, 9.750253e-006, 1.016351e-005, 1.062445e-005, 
    1.118076e-005, 1.188012e-005, 1.25318e-005, 1.326295e-005, 1.407357e-005, 
    1.499546e-005, 1.596503e-005, 1.707765e-005, 1.822204e-005, 
    1.944593e-005, 2.095593e-005, 2.249769e-005, 2.419841e-005, 2.59786e-005, 
    2.796543e-005, 3.003174e-005, 3.216161e-005, 3.427559e-005, 
    3.643726e-005, 3.86148e-005, 4.076057e-005, 4.279509e-005, 4.459117e-005, 
    4.632368e-005, 4.780186e-005, 4.885091e-005, 4.978871e-005, 
    5.029731e-005, 5.063112e-005, 5.026555e-005, 4.869199e-005, 
    4.784955e-005, 4.60217e-005, 4.457527e-005, 4.255668e-005, 4.025197e-005, 
    3.707306e-005, 3.42915e-005, 3.28133e-005, 3.058805e-005, 2.98887e-005, 
    2.81244e-005, 2.71866e-005, 2.669387e-005, 2.655083e-005, 2.666209e-005, 
    2.704357e-005, 2.814029e-005, 2.890323e-005, 2.977742e-005, 
    3.046089e-005, 3.01589e-005, 3.30517e-005, 3.464115e-005, 3.564251e-005, 
    3.65485e-005, 3.869427e-005, 4.004531e-005, 4.106258e-005, 4.18573e-005, 
    4.247719e-005, 4.281098e-005, 4.281098e-005, 4.233413e-005, 
    4.161887e-005, 4.052217e-005, 3.904395e-005, 3.740682e-005, 
    3.548358e-005, 3.340138e-005, 3.12874e-005, 2.925292e-005, 2.693229e-005, 
    2.489778e-005,
  3.179603e-005, 2.826744e-005, 2.539052e-005, 2.310169e-005, 2.121023e-005, 
    1.982741e-005, 1.882605e-005, 1.793595e-005, 1.699816e-005, 
    1.620343e-005, 1.54246e-005, 1.469346e-005, 1.410537e-005, 1.348547e-005, 
    1.281789e-005, 1.19278e-005, 1.122844e-005, 1.037014e-005, 9.654883e-006, 
    9.066789e-006, 8.589952e-006, 8.160798e-006, 8.113118e-006, 
    8.160805e-006, 8.415114e-006, 8.733008e-006, 9.003212e-006, 
    9.559524e-006, 1.024299e-005, 1.108539e-005, 1.213443e-005, 
    1.354905e-005, 1.54087e-005, 1.769754e-005, 2.079699e-005, 2.494548e-005, 
    3.017478e-005, 3.661209e-005, 4.425738e-005, 5.322193e-005, 
    6.285406e-005, 7.393256e-005, 8.434356e-005, 9.573987e-005, 0.0001053561, 
    0.0001123338, 0.0001222997, 0.0001296748, 0.0001355399, 0.000138083, 
    0.0001419613, 0.0001445998, 0.0001430899, 0.0001458078, 0.0001398155, 
    0.000145919, 0.0001432964, 0.0001389572, 0.0001336961, 0.0001260985, 
    0.0001172293, 0.0001071045, 9.513591e-005, 8.366004e-005, 7.34716e-005, 
    6.484083e-005, 5.778362e-005, 5.252258e-005, 4.900986e-005, 4.68323e-005, 
    4.786545e-005, 4.953438e-005, 5.250667e-005, 5.592399e-005, 
    6.012016e-005, 6.434813e-005, 6.773365e-005, 7.115098e-005, 
    7.245431e-005, 7.466368e-005, 7.68731e-005, 7.536306e-005, 7.809693e-005, 
    7.404381e-005, 7.60624e-005, 7.471137e-005, 7.388482e-005, 7.196158e-005, 
    6.922771e-005, 6.542896e-005, 6.067645e-005, 5.541537e-005, 
    5.026552e-005, 4.529055e-005, 4.025195e-005, 3.578558e-005,
  2.437326e-005, 1.9287e-005, 1.563125e-005, 1.302452e-005, 1.130791e-005, 
    1.008403e-005, 9.241608e-006, 8.876035e-006, 9.209834e-006, 
    1.038604e-005, 1.175297e-005, 1.307221e-005, 1.432788e-005, 
    1.548818e-005, 1.645775e-005, 1.701406e-005, 1.680744e-005, 1.57584e-005, 
    1.383515e-005, 1.13556e-005, 9.162144e-006, 7.668063e-006, 7.127644e-006, 
    7.270697e-006, 7.922376e-006, 8.431001e-006, 8.542269e-006, 
    8.589952e-006, 8.574058e-006, 8.494586e-006, 8.510473e-006, 
    9.289306e-006, 1.083109e-005, 1.323115e-005, 1.663259e-005, 
    2.094003e-005, 2.670977e-005, 3.42279e-005, 4.325602e-005, 5.477961e-005, 
    6.817869e-005, 8.203878e-005, 9.77903e-005, 0.0001102039, 0.0001201062, 
    0.0001315981, 0.0001402129, 0.0001442819, 0.000146237, 0.0001453469, 
    0.0001436143, 0.000144107, 0.000142756, 0.000137495, 0.0001362711, 
    0.0001382898, 0.0001404196, 0.0001429309, 0.0001449496, 0.0001438051, 
    0.000139609, 0.0001349837, 0.0001322179, 0.0001270521, 0.0001208215, 
    0.0001152744, 0.0001103788, 0.000106437, 0.0001005877, 9.539019e-005, 
    9.149607e-005, 8.78562e-005, 8.572632e-005, 8.574221e-005, 8.561506e-005, 
    8.580578e-005, 8.574221e-005, 8.803103e-005, 9.144837e-005, 
    9.278351e-005, 9.332394e-005, 9.198877e-005, 8.998608e-005, 
    8.667997e-005, 8.230898e-005, 7.954333e-005, 7.920954e-005, 
    8.075131e-005, 8.184803e-005, 8.078309e-005, 7.84625e-005, 7.078541e-005, 
    6.069237e-005, 4.983638e-005, 3.972743e-005, 3.114436e-005,
  1.017943e-005, 9.511874e-006, 1.181656e-005, 1.486832e-005, 1.704587e-005, 
    1.745913e-005, 1.682335e-005, 1.509083e-005, 1.291326e-005, 
    1.089467e-005, 9.909192e-006, 9.543604e-006, 1.032244e-005, 
    1.270663e-005, 1.660081e-005, 2.16394e-005, 2.794955e-005, 3.42279e-005, 
    3.850354e-005, 3.826513e-005, 3.400538e-005, 2.779061e-005, 
    2.128973e-005, 1.655313e-005, 1.408948e-005, 1.310401e-005, 1.22139e-005, 
    1.089464e-005, 9.098556e-006, 7.032264e-006, 5.411024e-006, 
    4.807029e-006, 5.713009e-006, 8.049516e-006, 1.097413e-005, 
    1.380336e-005, 1.580609e-005, 1.728429e-005, 1.917574e-005, 
    2.349906e-005, 3.042912e-005, 4.00612e-005, 5.603525e-005, 7.684124e-005, 
    0.0001007785, 0.000128594, 0.000325782, 0.0003373057, 0.0003322514, 
    0.0003245741, 0.0003057232, 0.0002931665, 0.0002834706, 0.0002746491, 
    0.0002693563, 0.000262776, 0.000268657, 0.0001943338, 0.0001895496, 
    0.0001865297, 0.0001820791, 0.0001748472, 0.0001662164, 0.0001634508, 
    0.0001598268, 0.0001574426, 0.0001560598, 0.0001541364, 0.0001494317, 
    0.0001459984, 0.0001454581, 0.0001441547, 0.0001441071, 0.0001452515, 
    0.0001510212, 0.0001560598, 0.0001582215, 0.0001624812, 0.0001662482, 
    0.0001733849, 0.0002080668, 0.0002135822, 0.0002231349, 0.0002316067, 
    0.0002389023, 0.0002431144, 0.0002455303, 0.0002440363, 0.0002666224, 
    0.0001668682, 0.0001369068, 0.0001046408, 7.447295e-005, 4.742041e-005, 
    2.731377e-005, 1.547231e-005,
  3.638957e-005, 2.349907e-005, 1.865119e-005, 1.696643e-005, 1.625114e-005, 
    1.604448e-005, 1.774519e-005, 2.136918e-005, 2.632829e-005, 
    3.305171e-005, 3.545178e-005, 3.324244e-005, 2.801312e-005, 
    2.198909e-005, 1.958899e-005, 2.337193e-005, 3.152582e-005, 
    4.300171e-005, 5.56856e-005, 6.267917e-005, 6.263156e-005, 5.482725e-005, 
    3.858301e-005, 2.235464e-005, 1.227751e-005, 9.432377e-006, 
    1.151458e-005, 1.397824e-005, 1.55677e-005, 1.528159e-005, 1.466169e-005, 
    1.575841e-005, 1.855587e-005, 2.299044e-005, 2.821976e-005, 
    3.282916e-005, 3.446631e-005, 3.343319e-005, 3.19073e-005, 3.336958e-005, 
    3.925058e-005, 4.754755e-005, 5.667104e-005, 6.887806e-005, 
    8.701376e-005, 0.0001140504, 0.0002931665, 0.0003072966, 0.0002735524, 
    0.0002395699, 0.0002088457, 0.0001953354, 0.0002030761, 0.0002259321, 
    0.0002485341, 0.0002787977, 0.0003278167, 0.0003788064, 0.0004147121, 
    0.0004513809, 0.0004788628, 0.0004979044, 0.0004993351, 0.0004861108, 
    0.000480786, 0.0004778455, 0.0004834721, 0.000519664, 0.0005511829, 
    0.0005689691, 0.0004648117, 0.0005700816, 0.0006002974, 0.00059839, 
    0.0005608788, 0.0005290578, 0.0003873578, 0.0003507367, 0.0003193289, 
    0.000300049, 0.0002951215, 0.0003017496, 0.0003326804, 0.0003699054, 
    0.0004154909, 0.0004610447, 0.0004931201, 0.0005077749, 0.0005021323, 
    0.0004913082, 0.0004894644, 0.0002696742, 0.0002073993, 0.0001472065, 
    9.283115e-005, 5.643265e-005,
  0.0006837754, 0.0005716712, 0.0002162686, 0.0001357467, 7.318554e-005, 
    3.627833e-005, 2.159172e-005, 2.496131e-005, 4.440051e-005, 
    7.614191e-005, 0.0001036554, 0.0001231264, 0.0001311848, 0.0001152902, 
    8.687071e-005, 6.225004e-005, 5.048804e-005, 4.835817e-005, 
    6.126455e-005, 7.823997e-005, 9.839423e-005, 0.0001093456, 9.605772e-005, 
    6.74476e-005, 4.726145e-005, 3.804261e-005, 4.01407e-005, 4.920061e-005, 
    5.810158e-005, 6.479316e-005, 6.010424e-005, 5.112385e-005, 
    4.277917e-005, 3.656442e-005, 3.664388e-005, 3.913933e-005, 
    4.247716e-005, 3.928237e-005, 3.281329e-005, 3.85989e-005, 5.074235e-005, 
    6.480905e-005, 7.688889e-005, 8.67754e-005, 0.0001967023, 0.0001223475, 
    0.0001213937, 6.538117e-005, 4.373281e-005, 3.370317e-005, 2.764747e-005, 
    2.901419e-005, 3.243168e-005, 3.478397e-005, 4.29221e-005, 6.477698e-005, 
    9.610527e-005, 0.0001441387, 0.0001892317, 0.0002308118, 0.0002741246, 
    0.0003110953, 0.0003496238, 0.000378107, 0.0003879773, 0.0003886924, 
    0.0003973073, 0.0004149345, 0.0004456905, 0.0005002725, 0.0005527721, 
    0.000609071, 0.0005588122, 0.0004817233, 0.0004288263, 0.0004098483, 
    0.0003956228, 0.0003945897, 0.0004137107, 0.0004310041, 0.0005110652, 
    0.0005391031, 0.0005823524, 0.0006520658, 0.0007246564, 0.0008012205, 
    0.0008600622, 0.0008855889, 0.0008948555, 0.0009282022, 0.000959896, 
    0.001016481, 0.001068408, 0.001054962, 0.0009903818, 0.0008460432,
  0.0009709587, 0.001004989, 0.001025413, 0.0009868373, 0.0009286315, 
    0.0008639721, 0.0008427373, 0.000825396, 0.0007804781, 0.0007396927, 
    0.0007279464, 0.0007503896, 0.0007590204, 0.0007579236, 0.0007332871, 
    0.0006862551, 0.0006385238, 0.0005753904, 0.0005455404, 0.0005485127, 
    0.0005443802, 0.0005345414, 0.0004857131, 0.0004303365, 0.0003643741, 
    0.0002814839, 0.0002161572, 0.0001634667, 0.0001343952, 0.0001287209, 
    0.0001368432, 0.0001332189, 0.0001472542, 0.0002248674, 0.0002503146, 
    0.0002967268, 0.0005563328, 0.0003583657, 0.0003159908, 0.0002960907, 
    0.0003106662, 0.0003093309, 0.0003034978, 0.000282787, 0.0002099264, 
    0.000106103, 1.110113e-005, -4.836055e-005, -7.042196e-005, 
    -7.816264e-005, -6.153737e-005, -3.057439e-005, -1.512491e-005, 
    -1.461618e-005, -2.758624e-005, -2.655317e-005, -3.283611e-006, 
    4.516332e-005, 9.179791e-005, 0.0001337121, 0.0001785029, 0.0002351508, 
    0.0003114445, 0.000385243, 0.0004351675, 0.00046435, 0.0005008755, 
    0.0005370677, 0.0005662027, 0.0005950197, 0.0006041115, 0.0006026013, 
    0.0005912366, 0.0005721154, 0.0005320294, 0.0004839324, 0.0004373617, 
    0.0004127254, 0.0004764465, 0.0006196725, 0.0006593135, 0.0005953219, 
    0.0005437441, 0.0005093005, 0.0005336511, 0.0005828447, 0.0006453739, 
    0.0007022447, 0.0007211752, 0.0007397085, 0.0007692089, 0.0008165112, 
    0.0008739859, 0.0009032001, 0.0009194603, 0.0009406637,
  0.0005235097, 0.000532395, 0.0005316958, 0.0005087443, 0.0004676569, 
    0.000446978, 0.000458708, 0.0004856014, 0.0004874768, 0.0004713277, 
    0.0004640324, 0.0004912913, 0.0005250038, 0.0005443792, 0.0005607507, 
    0.000576884, 0.0006000104, 0.0006032847, 0.0005612595, 0.0004986513, 
    0.0004390304, 0.0004020599, 0.0003757386, 0.000356172, 0.0003464289, 
    0.0003261634, 0.0002854576, 0.0002570697, 0.0002364698, 0.0002273303, 
    0.0002220692, 0.0002217195, 0.0002452596, 0.000280228, 0.0003266078, 
    0.0003579836, 0.0003752769, 0.0003768504, 0.0003766594, 0.0004070816, 
    0.0004407302, 0.0004553059, 0.0004440849, 0.0004185108, 0.0003516739, 
    0.0002357704, 9.798072e-005, -3.999099e-006, -5.829474e-005, 
    -0.000103801, -0.0001475271, -0.0001672362, -0.0001702881, -0.0001527565, 
    -0.0001216033, -7.528625e-005, -1.700083e-005, 4.478171e-005, 
    8.100504e-005, 0.0001036711, 0.0001471583, 0.0002077483, 0.0002584364, 
    0.0003173258, 0.0004083542, 0.0004984285, 0.0005764388, 0.0006237254, 
    0.0006562774, 0.0006851419, 0.0007300917, 0.0007811608, 0.0008201986, 
    0.0008304031, 0.0008141743, 0.00077412, 0.0007275804, 0.0006699944, 
    0.0005957033, 0.0005528196, 0.0005740705, 0.00055479, 0.0004562915, 
    0.0003741011, 0.0004053495, 0.0004500614, 0.0004985719, 0.0005295502, 
    0.0005291051, 0.0005240345, 0.0005215555, 0.0005126067, 0.0005059622, 
    0.0005071384, 0.0005129559, 0.0005186622,
  0.0004848698, 0.0004716143, 0.0004537329, 0.0004212605, 0.0003768187, 
    0.0003520073, 0.0003548367, 0.0003732112, 0.0003887084, 0.0003989441, 
    0.0004193215, 0.0004452453, 0.0004547182, 0.0004673703, 0.0004884307, 
    0.0005102218, 0.0005411534, 0.0005700332, 0.0005675377, 0.0005251472, 
    0.0004706606, 0.0004328, 0.00039683, 0.0003927136, 0.0004096413, 
    0.0004166192, 0.000410134, 0.0003866898, 0.0003667576, 0.0003382587, 
    0.0002971399, 0.0002582613, 0.0002166973, 0.0001836522, 0.0001787883, 
    0.0002082251, 0.0002377098, 0.0002708659, 0.0003262265, 0.0003936198, 
    0.0004595988, 0.0005145464, 0.0005705585, 0.0005557444, 0.0004941854, 
    0.0004327213, 0.0003661541, 0.0002601058, 0.0001125885, -1.563272e-005, 
    -9.098928e-005, -0.0001283097, -0.000140707, -0.0001436956, -0.000147908, 
    -0.0001298841, -5.978858e-005, 2.333988e-005, 4.308112e-005, 
    6.784452e-005, 0.0001608911, 0.0002612351, 0.0003140992, 0.0003658207, 
    0.0004821694, 0.0005884715, 0.0006405106, 0.0006646859, 0.0007085237, 
    0.0007815589, 0.0008669919, 0.0009311903, 0.0009573847, 0.0009567016, 
    0.0009251349, 0.0008687563, 0.0007986138, 0.0007628193, 0.0007288526, 
    0.0007008305, 0.0006664353, 0.0006246478, 0.0005509281, 0.0004480425, 
    0.0004087831, 0.0004024254, 0.0004358198, 0.0004592645, 0.000470724, 
    0.0004924042, 0.0005226512, 0.0005202354, 0.0004942953, 0.0004815641, 
    0.0004825653, 0.0004890184,
  0.0005094432, 0.000520363, 0.0005458575, 0.000532602, 0.0004993821, 
    0.0004882561, 0.0004997319, 0.0005079652, 0.0005145455, 0.0005315212, 
    0.0005445546, 0.0005540438, 0.0005565071, 0.00057245, 0.0006204196, 
    0.0006703609, 0.0007305052, 0.0007845149, 0.0007786178, 0.0006854446, 
    0.0006216434, 0.0005915873, 0.000531299, 0.0004994143, 0.0004904182, 
    0.0004986832, 0.0005092216, 0.0005110172, 0.0004897662, 0.000441256, 
    0.0003928896, 0.0003795535, 0.0003558868, 0.000316977, 0.0002964726, 
    0.0003217924, 0.0003560614, 0.0003837338, 0.0004231208, 0.0004663537, 
    0.0005103974, 0.0005708127, 0.0006218343, 0.0006309263, 0.0006260942, 
    0.0006024749, 0.0005435375, 0.0004558316, 0.0003210139, 0.0001943815, 
    0.0001431536, 0.0001238734, 9.442074e-005, 6.709807e-005, 3.273366e-005, 
    2.497714e-005, 6.078789e-005, 0.0001246519, 0.0001617023, 0.0001891367, 
    0.0002614888, 0.0003481777, 0.0004182886, 0.0005021961, 0.0006151274, 
    0.0006744773, 0.0006834418, 0.0007014503, 0.0007361639, 0.0007860572, 
    0.00082538, 0.0008400036, 0.0008590766, 0.0008676755, 0.0008491902, 
    0.0007592752, 0.0007371819, 0.0008078646, 0.0008157799, 0.000734495, 
    0.0007327786, 0.0006973017, 0.0006482196, 0.0005289628, 0.0004519057, 
    0.0005256729, 0.0006061615, 0.000653083, 0.0006524953, 0.0006441027, 
    0.0006414955, 0.0006447383, 0.0006297496, 0.0005848315, 0.0005420432, 
    0.000515833,
  0.0007602284, 0.0007659663, 0.0007852945, 0.0007907301, 0.0007906663, 
    0.0008018082, 0.0008069421, 0.0008070851, 0.0007917313, 0.0007793182, 
    0.0007842928, 0.0008079596, 0.0008416083, 0.0008732388, 0.0009099394, 
    0.0009683361, 0.001060016, 0.001138408, 0.001128077, 0.001035539, 
    0.001003718, 0.001020296, 0.0009832615, 0.0009162338, 0.0008609048, 
    0.0008332003, 0.0008319449, 0.0008205166, 0.0007796674, 0.000724752, 
    0.0006717434, 0.0006356151, 0.000621628, 0.0006009168, 0.0005711149, 
    0.0005483539, 0.0005533611, 0.0005859449, 0.0006355359, 0.0006900863, 
    0.0007511852, 0.0007969295, 0.0008009989, 0.0007942114, 0.0008096448, 
    0.0007908102, 0.0007013879, 0.0006187358, 0.0005366877, 0.0005052323, 
    0.0005230024, 0.0005335878, 0.0005102549, 0.0004749373, 0.000436727, 
    0.0004042219, 0.0003951471, 0.0004149349, 0.0004415899, 0.0004677372, 
    0.0005298369, 0.0005775839, 0.0006252681, 0.0006717439, 0.0007313327, 
    0.0007427135, 0.0007468136, 0.0007541254, 0.0007659825, 0.0007798276, 
    0.0008023335, 0.0008270182, 0.0008671521, 0.0008904692, 0.0008683596, 
    0.0008329949, 0.0008796449, 0.0008474896, 0.0008234098, 0.0008681538, 
    0.0008267476, 0.000665227, 0.0005513895, 0.0004655435, 0.0005452065, 
    0.0007073474, 0.0008041454, 0.0008387477, 0.0008565974, 0.0008582342, 
    0.0008367128, 0.0008304506, 0.000811568, 0.0007699081, 0.0007505328, 
    0.0007522656,
  0.0009662705, 0.0009600711, 0.001016068, 0.001068011, 0.001097734, 
    0.001141, 0.001208297, 0.001241055, 0.001242216, 0.001278186, 
    0.001335199, 0.00140841, 0.001461863, 0.001460687, 0.001469747, 
    0.001509467, 0.001562444, 0.00160687, 0.001604008, 0.001715525, 
    0.001859657, 0.001833097, 0.001646876, 0.001437592, 0.001303506, 
    0.001237908, 0.001197854, 0.001132019, 0.00105822, 0.001009646, 
    0.0009741224, 0.0009526326, 0.0009477208, 0.0009279647, 0.0009194291, 
    0.0009247698, 0.0009075403, 0.0009132624, 0.0009377403, 0.000977857, 
    0.00105687, 0.001120226, 0.001129953, 0.00114785, 0.001216133, 
    0.001241614, 0.001117158, 0.001037097, 0.0009595156, 0.0009275042, 
    0.001000317, 0.001063084, 0.001016449, 0.0009193979, 0.0008384306, 
    0.0007996168, 0.0007784609, 0.0007833876, 0.0007866621, 0.000785931, 
    0.0008106632, 0.000833408, 0.0008256836, 0.0008169413, 0.0008397661, 
    0.000885685, 0.0009232434, 0.0009363089, 0.0009321449, 0.0009466726, 
    0.0009591971, 0.0009583551, 0.0009557335, 0.0009608977, 0.000954397, 
    0.0009326544, 0.0009113229, 0.000772404, 0.0006374433, 0.001044424, 
    0.0009776512, 0.0007306812, 0.0005812724, 0.000593558, 0.0007524556, 
    0.000979193, 0.001105698, 0.001111913, 0.001123244, 0.001153922, 
    0.001129365, 0.001098942, 0.001068011, 0.001036684, 0.00103352, 
    0.001017912,
  0.001335041, 0.001308911, 0.001309101, 0.00136168, 0.001452962, 
    0.001660084, 0.001923935, 0.002084804, 0.002184749, 0.002307915, 
    0.002425901, 0.002402616, 0.002253637, 0.002087792, 0.001993315, 
    0.00197793, 0.002014692, 0.002068877, 0.002153596, 0.00222156, 
    0.002183668, 0.001983825, 0.00169251, 0.001477106, 0.001365256, 
    0.001322229, 0.001332323, 0.001304125, 0.001262912, 0.001263944, 
    0.001256792, 0.001277518, 0.001323644, 0.001308099, 0.00128502, 
    0.001307877, 0.001323676, 0.001323692, 0.001315284, 0.001455458, 
    0.001761572, 0.001812196, 0.001691922, 0.001634622, 0.00168302, 
    0.001713793, 0.001565417, 0.001599813, 0.001670131, 0.001665856, 
    0.001631475, 0.001510422, 0.001352652, 0.00122896, 0.001145847, 
    0.001101311, 0.001082349, 0.001080075, 0.001095796, 0.00110554, 
    0.001115171, 0.001154542, 0.00116616, 0.00115788, 0.001186077, 
    0.001223032, 0.001255616, 0.001295019, 0.001249243, 0.001200588, 
    0.001180004, 0.001138536, 0.001103838, 0.001049272, 0.0009430805, 
    0.000900913, 0.0008931719, 0.0005390393, 0.0004177643, 0.001182866, 
    0.001193532, 0.001038146, 0.001037844, 0.001180578, 0.001283431, 
    0.001438784, 0.001541273, 0.001489345, 0.00144632, 0.001463152, 
    0.001467268, 0.001489266, 0.001495099, 0.00147407, 0.001465217, 
    0.001408219,
  0.001441823, 0.001360602, 0.001329957, 0.001427723, 0.001709614, 
    0.002014282, 0.002193097, 0.002507253, 0.002652115, 0.002518952, 
    0.00219208, 0.001943552, 0.001788754, 0.001724906, 0.001742723, 
    0.001829441, 0.001962114, 0.002038964, 0.002006142, 0.001915957, 
    0.001812944, 0.001711997, 0.001571251, 0.001496418, 0.001466171, 
    0.001400447, 0.001363127, 0.001380165, 0.001430329, 0.00154558, 
    0.001565656, 0.001551703, 0.001515701, 0.001447258, 0.001537491, 
    0.001593983, 0.001593885, 0.001649405, 0.001713507, 0.002027567, 
    0.002276066, 0.002513085, 0.00246669, 0.002244706, 0.002148099, 
    0.002162785, 0.002124226, 0.002037375, 0.001936304, 0.001883326, 
    0.001700492, 0.00164311, 0.001607538, 0.00158012, 0.001547918, 
    0.001473054, 0.001459035, 0.001460497, 0.001484483, 0.001542562, 
    0.001521215, 0.001527906, 0.001532852, 0.001514427, 0.001562908, 
    0.001596844, 0.001610767, 0.001607111, 0.001491509, 0.001358328, 
    0.001263564, 0.001169659, 0.001040356, 0.0009066677, 0.0008217255, 
    0.0008592363, 0.0008044168, 0.0007577175, 0.0009288699, 0.001315332, 
    0.001300423, 0.001421317, 0.00173605, 0.001949783, 0.001964264, 
    0.00190984, 0.001885695, 0.001851936, 0.00184518, 0.001840934, 
    0.001823355, 0.001821605, 0.001782665, 0.001716273, 0.001657225, 
    0.001549364,
  0.001425675, 0.001345201, 0.001338033, 0.001480083, 0.001714321, 
    0.002010501, 0.002294981, 0.002290878, 0.002104516, 0.002019273, 
    0.001620255, 0.001737797, 0.001858898, 0.002010151, 0.002156571, 
    0.002233183, 0.002279643, 0.002205924, 0.00208956, 0.001959702, 
    0.001865352, 0.001809623, 0.001692306, 0.001636993, 0.001558948, 
    0.001461229, 0.001463836, 0.001523917, 0.001603628, 0.001706755, 
    0.001710124, 0.001784877, 0.001690288, 0.001624134, 0.001752706, 
    0.001704816, 0.001648881, 0.002076874, 0.00242765, 0.002750834, 
    0.002821648, 0.002874402, 0.002989764, 0.002694761, 0.002475972, 
    0.002496318, 0.002401555, 0.002220755, 0.002061172, 0.001888335, 
    0.001881866, 0.001981159, 0.00203296, 0.002013298, 0.001980189, 
    0.001921824, 0.001870739, 0.001831098, 0.001828809, 0.0018688, 
    0.001872487, 0.001897616, 0.00191758, 0.001899223, 0.001904721, 
    0.001836741, 0.00174673, 0.00162679, 0.001442746, 0.001323521, 
    0.001172841, 0.0009966176, 0.0009019338, 0.0008442048, 0.0007831836, 
    0.0008367952, 0.000944877, 0.001436639, 0.001623225, 0.001789183, 
    0.001772511, 0.002009802, 0.002274207, 0.002335019, 0.00222824, 
    0.002071806, 0.002074158, 0.002133699, 0.002145843, 0.002136258, 
    0.002100862, 0.002037585, 0.001919488, 0.001809196, 0.001742121, 
    0.001594539,
  0.001396509, 0.001417188, 0.001378787, 0.001555201, 0.001945825, 
    0.001988817, 0.002213471, 0.002212472, 0.002103627, 0.002057973, 
    0.002190216, 0.002519393, 0.002775216, 0.002949643, 0.003028591, 
    0.002987952, 0.00293221, 0.002791748, 0.002624203, 0.002452067, 
    0.00226634, 0.002105772, 0.00192664, 0.00183121, 0.001810499, 
    0.001748034, 0.001779758, 0.001814441, 0.001829159, 0.001871677, 
    0.001979712, 0.002346305, 0.002327229, 0.002245514, 0.00202253, 
    0.002125273, 0.002490133, 0.002663462, 0.003008453, 0.003422956, 
    0.003029454, 0.002795516, 0.002413346, 0.002296203, 0.002358987, 
    0.00242735, 0.002332873, 0.002203746, 0.002226203, 0.002383003, 
    0.002475128, 0.002538786, 0.002531125, 0.002445581, 0.002367634, 
    0.002227253, 0.002068291, 0.002012566, 0.00206651, 0.002147892, 
    0.002129707, 0.002162085, 0.00218758, 0.002129485, 0.002065986, 
    0.001898822, 0.00172864, 0.001531739, 0.001404743, 0.001271181, 
    0.001063772, 0.001002801, 0.0009221993, 0.0008850694, 0.0008039912, 
    0.0009559114, 0.001237468, 0.00148801, 0.002023913, 0.002390238, 
    0.002428447, 0.002595708, 0.002531779, 0.002521316, 0.002518155, 
    0.002465843, 0.002521046, 0.00260877, 0.002540599, 0.002443785, 
    0.002415238, 0.00229738, 0.002107727, 0.001913702, 0.001747494, 
    0.001551528,
  0.001402946, 0.001458101, 0.001556424, 0.001891417, 0.0022352, 0.002082184, 
    0.002367459, 0.002424967, 0.00232232, 0.002426187, 0.002661221, 
    0.00304517, 0.003263131, 0.003391448, 0.003450688, 0.003444567, 
    0.003372421, 0.003239449, 0.003009439, 0.002703341, 0.002423136, 
    0.002196385, 0.002010308, 0.001916101, 0.001931042, 0.001892419, 
    0.001899634, 0.001962926, 0.002191903, 0.002483265, 0.002728136, 
    0.00317794, 0.003146167, 0.002892645, 0.002325574, 0.002311875, 
    0.002795339, 0.003143051, 0.003463725, 0.003312789, 0.002774742, 
    0.002434677, 0.00215482, 0.00227638, 0.002533014, 0.002757542, 
    0.002767777, 0.002786756, 0.002883619, 0.002978031, 0.002946448, 
    0.002855627, 0.002817942, 0.002611088, 0.002388056, 0.002266891, 
    0.002198514, 0.002243781, 0.002277095, 0.0022585, 0.002137892, 
    0.00210302, 0.002063727, 0.001908008, 0.001760442, 0.001534836, 
    0.001435369, 0.001316653, 0.001260609, 0.001211668, 0.001043681, 
    0.001100202, 0.0009596152, 0.001010192, 0.0009682458, 0.001195475, 
    0.00152357, 0.0008130777, 0.002425044, 0.002751602, 0.002750723, 
    0.002867119, 0.002710875, 0.002690402, 0.002859887, 0.002852241, 
    0.002776645, 0.002680581, 0.002628572, 0.002498174, 0.002337146, 
    0.00214951, 0.001978789, 0.001745759, 0.00158513, 0.001408366,
  0.001711108, 0.001783588, 0.002050983, 0.002472122, 0.001785177, 
    0.001680879, 0.00244164, 0.002947801, 0.002748706, 0.002605177, 
    0.002987979, 0.003433265, 0.003357576, 0.003437512, 0.003515122, 
    0.003448479, 0.003206182, 0.003006751, 0.002770862, 0.002504738, 
    0.002232259, 0.002113175, 0.002084961, 0.002087155, 0.002090462, 
    0.002101857, 0.002221704, 0.002471821, 0.002748769, 0.00302236, 
    0.003366033, 0.003779196, 0.003845799, 0.002903151, 0.002854148, 
    0.003228562, 0.003267632, 0.003506275, 0.003213558, 0.00283959, 
    0.002475524, 0.002488097, 0.002662985, 0.002898734, 0.003079074, 
    0.003194196, 0.003163617, 0.003156813, 0.003219724, 0.003189253, 
    0.003073158, 0.002939356, 0.002901591, 0.002761243, 0.002642017, 
    0.002611134, 0.002606239, 0.002601057, 0.002418287, 0.002258085, 
    0.002146792, 0.00202984, 0.001958791, 0.001735106, 0.001543736, 
    0.001349011, 0.001287453, 0.001271766, 0.001184761, 0.001189831, 
    0.001172904, 0.001149921, 0.001074278, 0.001191405, 0.001149221, 
    0.00163159, 0.002126753, 0.0007390566, 0.002353549, 0.0029509, 
    0.00312558, 0.003025429, 0.00284199, 0.002778904, 0.002788456, 
    0.002840877, 0.002797976, 0.002560034, 0.002378216, 0.002264317, 
    0.002127543, 0.001943566, 0.001826817, 0.001745789, 0.001725795, 
    0.001654062,
  0.002135681, 0.002185449, 0.002461759, 0.002904726, 0.002293405, 
    0.002384691, 0.002609755, 0.002874892, 0.002831072, 0.002696269, 
    0.003149644, 0.003393512, 0.003124197, 0.003258474, 0.003414843, 
    0.003329489, 0.003084728, 0.002919093, 0.002743948, 0.002650457, 
    0.002485791, 0.0024736, 0.002400024, 0.002375817, 0.002418319, 
    0.00255773, 0.002791986, 0.003024155, 0.003226874, 0.003488181, 
    0.003882602, 0.004103411, 0.00435339, 0.003821143, 0.003893798, 
    0.003993696, 0.003831715, 0.003697705, 0.003170801, 0.002743157, 
    0.002845006, 0.002970798, 0.003141902, 0.003268454, 0.003365284, 
    0.00344746, 0.003395483, 0.003288386, 0.00325229, 0.003187472, 
    0.003067054, 0.002950341, 0.002919871, 0.002899494, 0.002880055, 
    0.002801346, 0.002779935, 0.00270593, 0.002521504, 0.002366787, 
    0.002261041, 0.002061326, 0.001930641, 0.001744932, 0.001637053, 
    0.00157373, 0.001476949, 0.001469031, 0.001386557, 0.001414134, 
    0.001400307, 0.001358995, 0.001433177, 0.001493959, 0.001489763, 
    0.002114432, 0.0023611, 0.001403197, 0.002497156, 0.003139488, 
    0.003374951, 0.003162393, 0.003126375, 0.002848951, 0.002664289, 
    0.002847664, 0.002723429, 0.002656212, 0.002429603, 0.002324969, 
    0.002256004, 0.002140656, 0.002091862, 0.002039535, 0.002102146, 
    0.002066921,
  0.002634389, 0.002605015, 0.002764568, 0.002875032, 0.002445499, 
    0.002226444, 0.002670566, 0.002715152, 0.002760389, 0.002675827, 
    0.002922734, 0.003308844, 0.003302995, 0.003340444, 0.003471285, 
    0.003291138, 0.003125388, 0.003046932, 0.003001649, 0.003031243, 
    0.002982432, 0.003003286, 0.002865193, 0.002868308, 0.002971767, 
    0.003119221, 0.00323409, 0.003357496, 0.003480569, 0.003564252, 
    0.003684858, 0.003840499, 0.004102202, 0.00442547, 0.004321439, 
    0.004294308, 0.004166326, 0.003639132, 0.003293745, 0.003090642, 
    0.003213698, 0.00336759, 0.00333715, 0.003242403, 0.003281759, 
    0.003380416, 0.003313148, 0.003206991, 0.003100814, 0.003045501, 
    0.002926832, 0.002820767, 0.002893344, 0.002926148, 0.002896443, 
    0.002887113, 0.002913196, 0.002786499, 0.002702115, 0.002532568, 
    0.002393777, 0.002272263, 0.002234783, 0.0021569, 0.002029968, 
    0.001976006, 0.001890302, 0.001893688, 0.001836372, 0.00182288, 
    0.001787785, 0.001815711, 0.001833909, 0.001832529, 0.00197367, 
    0.00253319, 0.002036741, 0.002219048, 0.002491724, 0.003156973, 
    0.003334448, 0.003061811, 0.002860347, 0.002819341, 0.002719617, 
    0.00273451, 0.002800867, 0.002807416, 0.00266327, 0.00273853, 
    0.002707649, 0.002655482, 0.002681978, 0.002647234, 0.00267319, 
    0.002633803,
  0.002929281, 0.002923861, 0.002962707, 0.002969669, 0.002779014, 
    0.002461236, 0.002714324, 0.002814542, 0.00267551, 0.002640588, 
    0.002841575, 0.003162786, 0.003426557, 0.003375202, 0.003302103, 
    0.003134431, 0.00313122, 0.003189299, 0.003286686, 0.00332577, 
    0.00329886, 0.003315948, 0.00322495, 0.003288036, 0.003345925, 
    0.003412332, 0.003452163, 0.003467105, 0.003515853, 0.003409011, 
    0.003333034, 0.003338341, 0.003392175, 0.003266068, 0.003486812, 
    0.0037149, 0.003724612, 0.003397182, 0.003259426, 0.003212729, 
    0.003244327, 0.00334133, 0.003195228, 0.003023615, 0.003004668, 
    0.00309708, 0.00301406, 0.002945015, 0.002959764, 0.002905961, 
    0.002889017, 0.002792921, 0.002857706, 0.002885858, 0.002905168, 
    0.002974007, 0.00300912, 0.002892658, 0.002881452, 0.002821008, 
    0.002725653, 0.002644625, 0.002608463, 0.002607733, 0.00249107, 
    0.002420211, 0.00237995, 0.002330104, 0.002327817, 0.00238548, 
    0.002382175, 0.00242641, 0.002392983, 0.00245076, 0.00266532, 
    0.002831914, 0.002476848, 0.002216254, 0.002536515, 0.003016433, 
    0.003149342, 0.00284512, 0.002881743, 0.002960928, 0.002592143, 
    0.002580317, 0.002954107, 0.003132366, 0.00303115, 0.003109811, 
    0.00307567, 0.003074748, 0.003035791, 0.003046583, 0.003047252, 
    0.002998902,
  0.003231516, 0.003167652, 0.003105519, 0.003043832, 0.002975138, 
    0.002992082, 0.003119953, 0.003060333, 0.002981893, 0.00276091, 
    0.002935385, 0.003214778, 0.003303183, 0.00327103, 0.003214922, 
    0.003155777, 0.003234964, 0.003219021, 0.003414892, 0.003449492, 
    0.00335527, 0.00329975, 0.003325405, 0.003383674, 0.003404988, 
    0.003360691, 0.003298813, 0.003281949, 0.003462065, 0.003499052, 
    0.003361436, 0.003308367, 0.003352331, 0.003325164, 0.003153043, 
    0.003208341, 0.003209533, 0.00318628, 0.003101166, 0.002973482, 
    0.003049156, 0.003132522, 0.003117772, 0.003091928, 0.002983971, 
    0.002965583, 0.002939131, 0.002928134, 0.002946524, 0.002915496, 
    0.002998691, 0.002929438, 0.003003713, 0.003018923, 0.002982158, 
    0.002966471, 0.002973957, 0.002976011, 0.002937974, 0.002924019, 
    0.002869278, 0.0028434, 0.002860505, 0.002810612, 0.002767887, 
    0.002813552, 0.002824249, 0.002823027, 0.002849221, 0.002880406, 
    0.002936497, 0.003000697, 0.00306607, 0.003115376, 0.00301883, 
    0.002581525, 0.002411472, 0.002402285, 0.002751898, 0.002998088, 
    0.002818799, 0.002657946, 0.00274368, 0.003070824, 0.002946114, 
    0.002617717, 0.002721572, 0.003062906, 0.003086381, 0.003098082, 
    0.003145557, 0.003240606, 0.003232056, 0.003338248, 0.003252052, 
    0.003241051,
  0.003148513, 0.003185501, 0.003130347, 0.002917454, 0.003087051, 
    0.002871204, 0.003039401, 0.003075274, 0.003150217, 0.002966984, 
    0.002827542, 0.003150597, 0.003295189, 0.003370911, 0.003359292, 
    0.003335308, 0.003350059, 0.00333127, 0.003384724, 0.00336495, 
    0.00339604, 0.003405893, 0.003465641, 0.003453372, 0.003529761, 
    0.003422838, 0.003299354, 0.003306091, 0.003175916, 0.003332602, 
    0.003277704, 0.003244117, 0.003285332, 0.00318202, 0.003228605, 
    0.003368812, 0.003267657, 0.002880374, 0.002613203, 0.002779778, 
    0.002981462, 0.003072521, 0.003074365, 0.003062712, 0.002976406, 
    0.002914593, 0.002907932, 0.002859185, 0.002911206, 0.002906691, 
    0.002933029, 0.002847342, 0.002921633, 0.002975944, 0.002952356, 
    0.003017843, 0.003106441, 0.003163964, 0.003120793, 0.003101783, 
    0.003085969, 0.003064144, 0.0030555, 0.003059965, 0.003094759, 
    0.003120301, 0.003134511, 0.003143204, 0.003168462, 0.003243737, 
    0.003265578, 0.003281232, 0.003289022, 0.003224252, 0.003094202, 
    0.002858585, 0.002823428, 0.00266243, 0.002844673, 0.00291663, 
    0.002798406, 0.002921971, 0.002786247, 0.002564725, 0.003162788, 
    0.002942681, 0.002924211, 0.00301829, 0.003052907, 0.003097827, 
    0.003148658, 0.003165774, 0.003112497, 0.003174167, 0.003119443, 
    0.003172785,
  0.003063351, 0.003114898, 0.003069995, 0.00238475, 0.002818322, 
    0.002317341, 0.002666973, 0.002579395, 0.00304234, 0.0030264, 
    0.002599421, 0.003327407, 0.003259968, 0.003315756, 0.003386583, 
    0.003522862, 0.003645759, 0.003669856, 0.003527552, 0.003434394, 
    0.003473606, 0.00343789, 0.003462002, 0.003355158, 0.003364362, 
    0.003361087, 0.003500974, 0.003424428, 0.003018467, 0.003200615, 
    0.003200967, 0.002949515, 0.002694726, 0.003034152, 0.003211711, 
    0.003158735, 0.003009932, 0.002783941, 0.002844008, 0.003072521, 
    0.003087398, 0.002978886, 0.002834737, 0.002790568, 0.002714654, 
    0.00261781, 0.002551481, 0.002475284, 0.002465429, 0.002425676, 
    0.002401771, 0.002394872, 0.002423262, 0.00247371, 0.002555916, 
    0.002706947, 0.002840145, 0.002943173, 0.003040843, 0.003090866, 
    0.003176106, 0.003192844, 0.003175106, 0.003249427, 0.003278531, 
    0.003277753, 0.003311194, 0.003325658, 0.003301974, 0.003312912, 
    0.003224507, 0.003217099, 0.003144778, 0.003087876, 0.00294554, 
    0.002678689, 0.003256234, 0.003382944, 0.003543288, 0.003589734, 
    0.002900245, 0.002556209, 0.002128358, 0.002139258, 0.002595132, 
    0.003002649, 0.003018115, 0.003063589, 0.003128089, 0.003123814, 
    0.003133779, 0.00310358, 0.003132127, 0.00313494, 0.003085269, 0.003114993,
  0.002969701, 0.003135879, 0.003075177, 0.002320567, 0.001844177, 
    0.002278494, 0.002104688, 0.00187366, 0.002907014, 0.003115759, 
    0.002896843, 0.00313906, 0.003051447, 0.003376236, 0.003539776, 
    0.003632709, 0.003647793, 0.003602305, 0.003545212, 0.003476562, 
    0.003352107, 0.003277307, 0.003301736, 0.003359595, 0.003423966, 
    0.003462099, 0.0032761, 0.002671679, 0.002980841, 0.003153663, 
    0.003087766, 0.002538116, 0.002542457, 0.003117202, 0.003049379, 
    0.00299011, 0.00293467, 0.002936719, 0.003034947, 0.003152281, 
    0.00310323, 0.003002459, 0.002978267, 0.003019307, 0.003000297, 
    0.002956556, 0.002926229, 0.00286966, 0.002782844, 0.002739975, 
    0.002688413, 0.002601184, 0.002512159, 0.002496965, 0.002516339, 
    0.00253972, 0.002642717, 0.002777424, 0.002865575, 0.002944969, 
    0.003002793, 0.003055835, 0.00311029, 0.003139663, 0.003166396, 
    0.003241086, 0.003242819, 0.003298001, 0.003298845, 0.003361883, 
    0.003310798, 0.003290294, 0.003040083, 0.002933731, 0.002661521, 
    0.002414441, 0.003198345, 0.004074374, 0.004128131, 0.003108289, 
    0.002376997, 0.001718466, 0.002057819, 0.002903197, 0.002767695, 
    0.002826156, 0.002789505, 0.002909236, 0.002985356, 0.003019577, 
    0.003114484, 0.003150119, 0.003175393, 0.003139773, 0.003089782, 
    0.003057852,
  0.003147576, 0.003315438, 0.002530487, 0.002419353, 0.002265588, 
    0.002315227, 0.002319487, 0.00231437, 0.002844294, 0.003175918, 
    0.002709639, 0.002683667, 0.002944732, 0.002986962, 0.003430406, 
    0.003575951, 0.003662657, 0.003624635, 0.00355977, 0.003485303, 
    0.003340982, 0.003320716, 0.00318593, 0.003301691, 0.003394945, 
    0.003440434, 0.002798947, 0.002237963, 0.002994305, 0.003085857, 
    0.003036998, 0.002871171, 0.003136149, 0.003211426, 0.003064893, 
    0.00312251, 0.003229195, 0.003315995, 0.003367702, 0.003452545, 
    0.003506524, 0.00343007, 0.003360756, 0.003356066, 0.003368797, 
    0.003357479, 0.003348103, 0.003419088, 0.003376633, 0.003358353, 
    0.003345065, 0.003269328, 0.003168065, 0.003071139, 0.002982907, 
    0.002902545, 0.00283175, 0.002797483, 0.00274271, 0.00278216, 0.00279966, 
    0.002821736, 0.002820276, 0.00285979, 0.0029731, 0.003074605, 
    0.003157511, 0.003312752, 0.00332159, 0.003412046, 0.003256137, 
    0.003231565, 0.003245058, 0.003152441, 0.00297175, 0.002738371, 
    0.002924785, 0.003392816, 0.003077229, 0.001887505, 0.002078925, 
    0.002588042, 0.002800297, 0.002679404, 0.002653942, 0.002663096, 
    0.002617098, 0.002672585, 0.002715038, 0.002819626, 0.002817782, 
    0.003018051, 0.003163377, 0.003149785, 0.002837904, 0.002919095,
  0.003253388, 0.003225858, 0.003065119, 0.002483075, 0.002426316, 
    0.002703089, 0.002415604, 0.002476432, 0.002522714, 0.00273227, 
    0.002016175, 0.001931773, 0.002289498, 0.002303864, 0.003090834, 
    0.003334658, 0.003379783, 0.003520036, 0.003568623, 0.003836226, 
    0.003710657, 0.003520288, 0.0032716, 0.003328981, 0.003230548, 
    0.003172802, 0.00294303, 0.003011361, 0.002820274, 0.002802044, 
    0.002954219, 0.002888765, 0.002936004, 0.002937643, 0.003192034, 
    0.003305219, 0.003286781, 0.00333262, 0.003343033, 0.003352774, 
    0.003344368, 0.003327059, 0.00336042, 0.003369655, 0.003367461, 
    0.00339024, 0.003402287, 0.003445648, 0.003436938, 0.003420535, 
    0.003376571, 0.003336914, 0.003264101, 0.003196709, 0.003116472, 
    0.003072921, 0.002952535, 0.002871808, 0.002771275, 0.002665782, 
    0.002617558, 0.002652081, 0.002628809, 0.002695631, 0.002746159, 
    0.002901543, 0.003148753, 0.003301149, 0.003348356, 0.003370784, 
    0.003284046, 0.003242005, 0.003149388, 0.003059221, 0.002648696, 
    0.002535799, 0.003145129, 0.002717073, 0.002500511, 0.002663414, 
    0.002846075, 0.002718996, 0.002722908, 0.002588153, 0.002545841, 
    0.002513194, 0.002499031, 0.002527514, 0.002528293, 0.002591856, 
    0.002533332, 0.002875939, 0.002877846, 0.002803794, 0.003129316, 
    0.003178495,
  0.002335415, 0.002298795, 0.002162659, 0.002061249, 0.001932042, 
    0.002000991, 0.001806108, 0.001945155, 0.002101162, 0.00232898, 
    0.00195668, 0.001143241, 0.001104999, 0.001271812, 0.002589758, 
    0.002880454, 0.003051543, 0.003172675, 0.003285782, 0.003619473, 
    0.003747646, 0.004169582, 0.003579924, 0.003388045, 0.003168223, 
    0.00300605, 0.002794048, 0.00277485, 0.002674159, 0.00228428, 
    0.002797736, 0.002873505, 0.002891025, 0.002935989, 0.003046567, 
    0.003167842, 0.003175123, 0.003209423, 0.003222534, 0.003216257, 
    0.003222235, 0.003175711, 0.003130587, 0.003091455, 0.003040591, 
    0.003047634, 0.003043611, 0.003057662, 0.003037684, 0.003030069, 
    0.002979556, 0.00295586, 0.002930459, 0.002928758, 0.002852973, 
    0.002820611, 0.002752185, 0.002672616, 0.002612313, 0.00254546, 
    0.002466129, 0.002467688, 0.002492564, 0.002557207, 0.002584737, 
    0.002656085, 0.002732158, 0.003030099, 0.003406309, 0.003384342, 
    0.003385087, 0.003136516, 0.002791221, 0.002241303, 0.002806386, 
    0.002892263, 0.002804922, 0.002827955, 0.002721889, 0.002618226, 
    0.00259219, 0.002502179, 0.002504198, 0.002353741, 0.002331966, 
    0.002285776, 0.002311621, 0.002365409, 0.002348098, 0.002327451, 
    0.00237415, 0.002443133, 0.002222962, 0.00193516, 0.002053843, 0.002114465,
  0.001101723, 0.001157243, 0.001121941, 0.0009424281, 0.0005460004, 
    0.0009297119, 0.000943651, 0.0009186179, 0.001196185, 0.00186627, 
    0.002269582, 0.001683354, 0.0005399934, 0.0004473762, 0.0009641256, 
    0.002119599, 0.002665307, 0.002685763, 0.003119555, 0.003282953, 
    0.003341655, 0.00423763, 0.003913665, 0.003673991, 0.003416687, 
    0.00302287, 0.002831153, 0.002768099, 0.002217841, 0.00191489, 
    0.00239489, 0.002564041, 0.002514703, 0.0024877, 0.002677767, 
    0.002758576, 0.002836362, 0.002869599, 0.002889879, 0.00289182, 
    0.002889324, 0.00285016, 0.002794163, 0.00275816, 0.002733905, 
    0.002752883, 0.002764201, 0.002784801, 0.002763248, 0.002739357, 
    0.002689241, 0.002635537, 0.002554077, 0.00248732, 0.002452097, 
    0.002422169, 0.002349815, 0.00228236, 0.002182287, 0.002129503, 
    0.002056737, 0.00204407, 0.002031703, 0.002047344, 0.002112018, 
    0.002085298, 0.002203682, 0.002466384, 0.00251518, 0.002756558, 
    0.002740745, 0.0023097, 0.001705929, 0.002452079, 0.002722112, 
    0.002713909, 0.0026503, 0.002461314, 0.002466449, 0.002402475, 
    0.002317502, 0.002265162, 0.002172671, 0.002047454, 0.002044465, 
    0.00196598, 0.001977821, 0.001966648, 0.001990966, 0.001928102, 
    0.002062031, 0.002356892, 0.001646622, 0.001327681, 0.001082379, 
    0.001006832,
  0.0006086095, 0.0007573669, 0.0006625082, 0.0007559201, 6.835372e-005, 
    0.0006041755, 0.0004962671, 0.0003808406, 0.0005705899, 0.00139277, 
    0.00217941, 0.0009303321, 0.0003047213, 5.926169e-005, -0.0002965543, 
    0.0006063692, 0.002561725, 0.00267378, 0.002748295, 0.002602239, 
    0.002643485, 0.002922655, 0.003987721, 0.004386003, 0.003453724, 
    0.003202021, 0.002762534, 0.00276409, 0.002045167, 0.001490587, 
    0.001851012, 0.002112254, 0.002106993, 0.002081737, 0.002126432, 
    0.002199436, 0.00227805, 0.002383686, 0.002482486, 0.002541009, 
    0.002522969, 0.002509951, 0.002470723, 0.002358842, 0.002288365, 
    0.002300572, 0.002298206, 0.002296856, 0.002300194, 0.002295631, 
    0.002276272, 0.002212473, 0.00213931, 0.002103786, 0.002073984, 
    0.002023995, 0.001956125, 0.00192494, 0.001812295, 0.00172025, 
    0.001634721, 0.001611641, 0.00158915, 0.001571285, 0.001638503, 
    0.001668259, 0.001841764, 0.001863905, 0.001407472, 0.001243726, 
    0.001910282, 0.001755711, 0.001469593, 0.002201961, 0.002236979, 
    0.002290765, 0.002369253, 0.00228026, 0.002250268, 0.002212264, 
    0.002125797, 0.002043081, 0.002007765, 0.001940438, 0.001822388, 
    0.001698983, 0.001676921, 0.001643463, 0.001625184, 0.001561956, 
    0.001642333, 0.001758221, 0.001003733, 0.0003717013, 1.110137e-005, 
    0.0001278152,
  0.000724338, 0.0006124398, 0.0003395784, 0.0003372263, 0.0003996759, 
    0.0005078542, 0.0001204878, 0.0002300967, 0.0002905915, 0.001008215, 
    0.001679193, 0.0006600441, 0.0006243447, 0.0004316396, -0.0001467797, 
    0.0002513155, 0.002305902, 0.002317997, 0.001764131, 0.001591564, 
    0.001918786, 0.001992727, 0.002497538, 0.002650556, 0.003409905, 
    0.00325719, 0.002754966, 0.002623884, 0.00174927, 0.0008978471, 
    0.0009155869, 0.001012607, 0.001499124, 0.001649233, 0.001658722, 
    0.001734635, 0.001772447, 0.001849425, 0.001950324, 0.002045914, 
    0.002061554, 0.002072426, 0.001999199, 0.001948003, 0.001888796, 
    0.001763738, 0.001730549, 0.001769792, 0.001810945, 0.001867657, 
    0.001942487, 0.001930154, 0.001880324, 0.001865224, 0.001789884, 
    0.001755059, 0.001738179, 0.001668877, 0.001582983, 0.001534263, 
    0.001468762, 0.00144357, 0.001436292, 0.001400384, 0.001429471, 
    0.001433479, 0.001579738, 0.001593472, 0.001118827, 0.001568485, 
    0.001784844, 0.002067339, 0.00196002, 0.001818495, 0.001821592, 
    0.001852048, 0.001893136, 0.001982717, 0.002134812, 0.002211488, 
    0.002182575, 0.00207454, 0.0019762, 0.001897887, 0.001894502, 
    0.001748844, 0.001644973, 0.001601931, 0.00147118, 0.00143931, 
    0.001463946, 0.001376288, 0.0009129914, 0.0007302985, 0.0007346692, 
    0.0005731008,
  0.0004820095, 0.000781876, 0.0007343516, 0.000417287, 0.0007039774, 
    0.0008112341, 0.0002586592, 0.0003172942, 0.0006400014, 0.0005245118, 
    0.0006748897, 0.0004907993, 0.0006976346, 0.0005889479, 0.0008540223, 
    0.0007522018, 0.0006536716, 0.0007078876, 0.0006574383, 0.0008866224, 
    0.001861311, 0.001896357, 0.001541256, 0.0009955941, 0.001274592, 
    0.001829266, 0.001974033, 0.002033146, 0.00145684, 0.001117189, 
    0.001134514, 0.0008445024, 0.0008428972, 0.001188414, 0.001307752, 
    0.001360062, 0.00139773, 0.001513219, 0.001579627, 0.00157106, 
    0.001567627, 0.001634129, 0.001607633, 0.001578851, 0.001555582, 
    0.001439647, 0.001382522, 0.001335459, 0.001311202, 0.001350095, 
    0.001452455, 0.001520547, 0.001525681, 0.001538079, 0.001514937, 
    0.001492493, 0.001449959, 0.001419283, 0.001410734, 0.001376384, 
    0.001316126, 0.001268697, 0.001253819, 0.001288977, 0.001245825, 
    0.001305589, 0.001141095, 0.001115361, 0.001014955, 0.001374905, 
    0.001692208, 0.001916848, 0.00191809, 0.001762385, 0.00144508, 
    0.001580806, 0.001635897, 0.001669228, 0.00178324, 0.001938609, 
    0.002015062, 0.002032355, 0.001976677, 0.001904594, 0.00187306, 
    0.001758077, 0.001689938, 0.001618905, 0.001445476, 0.001355355, 
    0.00123915, 0.001215483, 0.001290043, 0.0007603876, 0.0006111525, 
    0.0002684663,
  0.0005741506, 0.0004247255, 0.0002001352, 0.0007165498, 0.001043725, 
    0.001401464, 0.0007192679, 0.0005883598, 0.001548902, 0.0007611029, 
    0.000577345, 0.0005497513, 0.0006766384, 0.0007634703, 0.0003418191, 
    0.0003169603, 0.0002508545, 0.0002295398, 0.0002780505, 0.0002511735, 
    0.0002478343, 0.0009750277, 0.0007140387, 0.0007543158, 0.0007828146, 
    0.001022012, 0.000992289, 0.001192528, 0.001436288, 0.001402432, 
    0.001625465, 0.001424064, 0.0009294422, 0.0005825744, 0.000887895, 
    0.001034061, 0.001042866, 0.001171947, 0.001254948, 0.001282589, 
    0.001297625, 0.001319321, 0.001315141, 0.001280379, 0.00127728, 
    0.00128847, 0.001252802, 0.001185426, 0.001136024, 0.001114282, 
    0.001158929, 0.001207534, 0.001218184, 0.001227005, 0.00123988, 
    0.001191926, 0.001115569, 0.001104506, 0.001113438, 0.00106976, 
    0.001091074, 0.001061129, 0.001065373, 0.00112218, 0.001079537, 
    0.001050035, 0.001002017, 0.0008680574, 0.0008946331, 0.001157132, 
    0.001055518, 0.001261211, 0.001073925, 0.001005356, 0.001080203, 
    0.001323551, 0.001418761, 0.001398461, 0.001470893, 0.001527001, 
    0.001639995, 0.001808668, 0.0018825, 0.001837932, 0.001731674, 
    0.001673358, 0.001654952, 0.001490586, 0.001384569, 0.001349871, 
    0.001212191, 0.001197028, 0.001202513, 0.001172375, 0.0008664676, 
    0.0007269611,
  0.0005910466, 0.0006127269, 0.0006143004, 0.00142499, 0.001582186, 
    0.001595219, 0.001466362, 0.001443951, 0.001610096, 0.001441089, 
    0.0006076721, 0.0001118085, 0.0001136209, 0.000954777, 0.0008154144, 
    0.0005564918, 0.0009296006, 0.001302281, 0.001028671, 0.0009276618, 
    0.0007959912, 0.0009109408, 0.0007620882, 0.0007108918, 0.0008560568, 
    0.0007810504, 0.0006756217, 0.0009803365, 0.0009559216, 0.0008916445, 
    0.0009086991, 0.001135959, 0.001029927, 0.0005815094, 0.001015462, 
    0.001002605, 0.0007536467, 0.0008558016, 0.001039989, 0.001115997, 
    0.001152953, 0.001155767, 0.00119544, 0.001210745, 0.001212874, 
    0.001205627, 0.001202035, 0.001205168, 0.001170961, 0.001128983, 
    0.00112644, 0.001089184, 0.001049336, 0.001018437, 0.0009769518, 
    0.000964093, 0.0009426186, 0.0009322073, 0.0009101629, 0.0008877357, 
    0.0009154873, 0.0009375163, 0.0009735343, 0.0009780796, 0.0008709338, 
    0.0008600145, 0.0009295535, 0.0009345915, 0.001087434, 0.0007076175, 
    0.0008318336, 0.0009988695, 0.0009852001, 0.0009777779, 0.001004433, 
    0.001096891, 0.001333881, 0.001392118, 0.001476965, 0.001500837, 
    0.001603198, 0.001665759, 0.001640567, 0.001665203, 0.001540748, 
    0.001409491, 0.001361123, 0.001256458, 0.0011873, 0.001211349, 
    0.001216357, 0.001199238, 0.001067265, 0.001035873, 0.00100445, 
    0.0006884015,
  0.0008766404, 0.001160328, 0.001304999, 0.001426085, 0.0014522, 
    0.001354686, 0.001289533, 0.001327887, 0.00138692, 0.001343607, 
    0.001269156, 0.001204942, 0.001001301, 0.001191384, 0.001068281, 
    0.0007965793, 0.000665131, 0.0007503894, 0.001128664, 0.0007691137, 
    0.0005496413, 0.0009402186, 0.00100688, 0.0009964691, 0.0009674933, 
    0.00106205, 0.0008217881, 0.0006335168, 0.000669518, 0.0006613166, 
    0.0005466691, 0.0005887896, 0.0005988029, 0.0005488782, 0.0005690167, 
    0.0008442313, 0.0008853986, 0.0008379202, 0.0009450023, 0.0009861854, 
    0.001041324, 0.001069282, 0.001095731, 0.001092393, 0.001102009, 
    0.001121861, 0.001144209, 0.001140935, 0.001094793, 0.001084573, 
    0.001119446, 0.001075354, 0.001026176, 0.001009296, 0.0009685904, 
    0.0009253891, 0.0008759573, 0.0008202628, 0.0008236007, 0.0008560098, 
    0.0008639256, 0.0008814414, 0.000927249, 0.000893123, 0.00101365, 
    0.001038383, 0.001033599, 0.0008666741, 0.0008337086, 0.00114068, 
    0.001039512, 0.001185265, 0.001265835, 0.001225987, 0.001157179, 
    0.001250083, 0.001361074, 0.001486928, 0.001537092, 0.001616534, 
    0.001687043, 0.001665664, 0.00149742, 0.001184837, 0.0007860744, 
    0.0007065693, 0.0008045435, 0.0007779999, 0.0007309197, 0.0007813852, 
    0.0009873947, 0.001074307, 0.001000093, 0.0009813062, 0.0007620412, 
    0.0006308467,
  0.0009472594, 0.001171374, 0.001222872, 0.001136851, 0.001275785, 
    0.001167208, 0.001268838, 0.001324533, 0.001323865, 0.001229721, 
    0.001153602, 0.001315537, 0.001180607, 0.0009002755, 0.0009434605, 
    0.00100963, 0.0008957447, 0.0009367843, 0.00105148, 0.0006184008, 
    0.000511955, 0.0006629687, 0.000800807, 0.0008502391, 0.0008646715, 
    0.0007925581, 0.0007541885, 0.0007458439, 0.0006668638, 0.0006061147, 
    0.0004854908, 0.000444435, 0.0004816125, 0.0004767805, 0.00040721, 
    0.0003505299, 0.0006374579, 0.0007617222, 0.0007894901, 0.0009340348, 
    0.0009489919, 0.0008891963, 0.0007851664, 0.0007163906, 0.0007065837, 
    0.0007290114, 0.0007684296, 0.0008354727, 0.0009024371, 0.0009228936, 
    0.0009021033, 0.0008736365, 0.0008741599, 0.0008838405, 0.0008740812, 
    0.0008710138, 0.000860523, 0.0008240771, 0.0008137929, 0.0008165906, 
    0.0008250941, 0.0008291313, 0.0008578845, 0.0009120526, 0.001234935, 
    0.001185837, 0.0008993538, 0.0006752561, 0.000625792, 0.0007359728, 
    0.0009864869, 0.000936578, 0.0009220187, 0.001030244, 0.0009179024, 
    0.001134164, 0.001202097, 0.001216514, 0.001494907, 0.001571487, 
    0.001325249, 0.001026081, 0.0008252533, 0.0006090398, 0.0004935651, 
    0.0003705886, 0.0003383229, 0.0002804035, 0.0002922295, 0.0004553236, 
    0.0006053359, 0.0007428401, 0.0008142549, 0.0008726511, 0.0007997425, 
    0.0008516698,
  0.0008591879, 0.0009784605, 0.001002636, 0.001038892, 0.001003748, 
    0.001064386, 0.0009422211, 0.001090565, 0.001232218, 0.001193498, 
    0.001097479, 0.001010187, 0.0008397645, 0.0007123696, 0.0007032617, 
    0.0005347319, 0.0004316079, 0.0004406678, 0.0004846323, 0.0005063284, 
    0.0005376723, 0.0005164847, 0.0004562447, 0.0005427112, 0.0006175269, 
    0.000491197, 0.0004990805, 0.0005645026, 0.0004996845, 0.0004743966, 
    0.0005060424, 0.0004593919, 0.00045634, 0.0004038084, 0.0003607818, 
    0.0002507755, 0.0002124696, 0.0005534715, 0.0005790142, 0.0006271114, 
    0.0006480601, 0.0005702404, 0.0005602902, 0.0005449839, 0.0005468912, 
    0.0005646932, 0.0005925875, 0.0006298285, 0.0006829957, 0.0007088403, 
    0.0007148809, 0.0007344629, 0.000764647, 0.0007642494, 0.0007453826, 
    0.0007310305, 0.0007493091, 0.0007909364, 0.0008056075, 0.0008105664, 
    0.0008392083, 0.0008276533, 0.0008473783, 0.0008807252, 0.001103026, 
    0.0008184502, 0.0007533142, 0.0007471789, 0.000675224, 0.0006501102, 
    0.0007000198, 0.0007433961, 0.0008361568, 0.001032805, 0.000791954, 
    0.0007565886, 0.0007009099, 0.0006845385, 0.0007693678, 0.001030611, 
    0.0008980818, 0.0007586866, 0.0006530511, 0.0005063126, 0.0003883746, 
    0.0003874209, 0.000262999, 2.35308e-005, -0.0001113187, -2.297666e-005, 
    0.0002179691, 0.0004737289, 0.000662636, 0.0007645516, 0.0008874326, 
    0.0008153035,
  0.0007795403, 0.0008651004, 0.0008766875, 0.0009644094, 0.0009962786, 
    0.0009069827, 0.00086456, 0.0008322464, 0.0008421012, 0.0008112499, 
    0.0006756056, 0.0006749541, 0.0006050179, 0.0004653679, 0.0004019646, 
    0.0003409137, 0.0002616474, 0.0003042291, 0.0003192178, 0.0002882711, 
    0.0003997714, 0.0004526048, 0.0004275549, 0.0004333247, 0.0003628323, 
    0.0003069788, 0.0003705571, 0.0003975143, 0.0003693968, 0.0003569672, 
    0.0004078615, 0.0003587952, 0.0002927691, 0.0002730597, 0.0002351673, 
    0.0001433918, 0.0001113167, 0.0002366771, 0.0005151818, 0.0009728661, 
    0.0008687088, 0.0006413527, 0.0005591463, 0.0005479881, 0.0005740868, 
    0.0005607356, 0.0005912848, 0.0006201018, 0.0006339459, 0.0006378235, 
    0.0006625713, 0.0007052165, 0.0007335723, 0.0007311087, 0.0007197601, 
    0.0007194425, 0.0007079984, 0.0007224148, 0.000750469, 0.000773564, 
    0.0008223606, 0.0008387156, 0.0007313634, 0.0006537028, 0.0005986919, 
    0.0006075294, 0.000659711, 0.0005788554, 0.0004950911, 0.000522827, 
    0.0005582243, 0.0005188378, 0.0004583269, 0.0004444828, 0.0004772097, 
    0.0004963467, 0.0004787515, 0.0004698347, 0.0004767806, 0.0005350979, 
    0.0009038679, 0.0007150401, 0.0007346859, 0.000595147, 0.0004861106, 
    0.0003842576, 0.0001485888, -0.0001892978, -0.0004015057, -0.0003407085, 
    -7.304456e-005, 0.0002408577, 0.000464065, 0.0005554268, 0.0006565959, 
    0.0007316503,
  0.0006983345, 0.0006328644, 0.0006760501, 0.000765394, 0.00077172, 
    0.0007757253, 0.000738834, 0.0007596086, 0.0006722044, 0.000550563, 
    0.0004734905, 0.0004358519, 0.0003524532, 0.0002933092, 0.0002704372, 
    0.0002459754, 0.000229159, 0.0002224515, 0.0002279192, 0.0002448629, 
    0.000273648, 0.0003151328, 0.0002995718, 0.0002769857, 0.0002531119, 
    0.0002419699, 0.0002624262, 0.0002474218, 0.0002148856, 0.0002167134, 
    0.0002284438, 0.0002005805, 0.0001823971, 0.0001778832, 0.0001605738, 
    8.852378e-005, 8.057646e-005, 0.0001822858, 0.0004783857, 0.0009478321, 
    0.001006769, 0.0008454551, 0.0005198229, 0.0006267936, 0.000682679, 
    0.0005935258, 0.0005483695, 0.0005492915, 0.0005841006, 0.0006219614, 
    0.0006952982, 0.0007972778, 0.0008618098, 0.0008430702, 0.0007770443, 
    0.0007753749, 0.0007346375, 0.0007377211, 0.0007469086, 0.0007386911, 
    0.0007017367, 0.0007215245, 0.0005487669, 0.0004354387, 0.0004329751, 
    0.0004656066, 0.000499049, 0.0004821689, 0.0004993986, 0.0005072824, 
    0.0005058835, 0.0004717261, 0.0004950274, 0.0005088876, 0.0004716943, 
    0.0004583109, 0.0004177003, 0.000404937, 0.0003578733, 0.0003347466, 
    0.0003978638, 0.0006513507, 0.0007813523, 0.0004804202, 0.000336638, 
    0.0003751346, 0.0002765558, 4.309695e-005, -0.0001460803, -0.0001695883, 
    -1.192978e-005, 0.0002280148, 0.0004160311, 0.0004911651, 0.0004928177, 
    0.0005929694,
  0.0004768753, 0.000481612, 0.0004319889, 0.0005839413, 0.0006496499, 
    0.0007070927, 0.0005581288, 0.0005657582, 0.0004447052, 0.0004262357, 
    0.0004094194, 0.0003706842, 0.0002811978, 0.0002156008, 0.0001933485, 
    0.0002000084, 0.0001857033, 0.0001765321, 0.0001673609, 0.0001989116, 
    0.0002251217, 0.0002343089, 0.0002655417, 0.0002712478, 0.0002611389, 
    0.0002423516, 0.0002246608, 0.0001967499, 0.0001688392, 0.0001766752, 
    0.0001787096, 0.0001618454, 0.0001456171, 0.0001391797, 0.0001103152, 
    7.682538e-005, 8.675945e-005, 0.0001829375, 0.0004356135, 0.0006859849, 
    0.0006949652, 0.0005717189, 0.0003741491, 0.0004489174, 0.0008930116, 
    0.0007369588, 0.0008358071, 0.000963361, 0.0009844054, 0.00108319, 
    0.001180433, 0.001121989, 0.0009663175, 0.0008857157, 0.0007942268, 
    0.0007079984, 0.0006954414, 0.0007034685, 0.000694281, 0.0006324197, 
    0.0005993117, 0.0004498709, 0.000405414, 0.0004099121, 0.0004312107, 
    0.0004181454, 0.0003917445, 0.0003585725, 0.0003543763, 0.0003820329, 
    0.0003838289, 0.0003951936, 0.0004185903, 0.0004231045, 0.000402966, 
    0.0003844966, 0.0003502438, 0.0003299146, 0.0002701351, 0.0002320677, 
    0.0002914657, 0.0004894325, 0.0004454363, 4.996359e-005, 5.051959e-005, 
    0.0003578095, 0.0005473676, 0.0004814048, 0.0003372096, 0.0002686568, 
    0.0003093947, 0.0004013926, 0.0004849494, 0.0005177408, 0.0005146251, 
    0.0005585575,
  0.0003628479, 0.0003608926, 0.0004611402, 0.0004297327, 0.0004879227, 
    0.0007233371, 0.0005020212, 0.0004696279, 0.0004304479, 0.0003791243, 
    0.0003277212, 0.0002813409, 0.000237901, 0.0001945406, 0.0001595566, 
    0.0001584281, 0.000192681, 0.0002075583, 0.0001909008, 0.0001591434, 
    0.0001403877, 0.0001770406, 0.0002110393, 0.000217556, 0.0002000878, 
    0.0001884688, 0.0002006281, 0.0002171426, 0.0002118498, 0.000186323, 
    0.00016628, 0.0001539776, 0.0001431534, 0.0001250177, 9.80605e-005, 
    8.272222e-005, 8.971585e-005, 9.602599e-005, 9.949101e-005, 
    9.790156e-005, 0.0001194864, 0.0001616706, 0.0002130259, 0.0002726782, 
    0.0003639608, 0.0005088874, 0.0006879874, 0.001258794, 0.00148278, 
    0.001443393, 0.001280251, 0.001069235, 0.0007521542, 0.0006278268, 
    0.0005339375, 0.0004492988, 0.0003937791, 0.000364835, 0.000363818, 
    0.0003620377, 0.0003451098, 0.0003109684, 0.0002896219, 0.0002971401, 
    0.0003090133, 0.0003132413, 0.0003069947, 0.0003108731, 0.000334556, 
    0.0003478277, 0.0003379573, 0.0003457933, 0.0003281186, 0.000314767, 
    0.0003077576, 0.0003112384, 0.0002701032, 0.000225535, 0.0001924743, 
    0.0001580308, 0.0001620997, 0.0002013118, 0.0001397043, 0.0001199475, 
    0.0002354055, 0.0002316227, 0.0003638812, 0.0004565145, 0.0005542338, 
    0.0005733394, 0.0005498952, 0.0004547979, 0.0002545579, 0.0002167448, 
    0.0003372892, 0.0003684745,
  0.0002956134, 0.0003234129, 0.0003267669, 0.0005462239, 0.0004975864, 
    0.000450173, 0.0004635085, 0.0004038402, 0.0003971169, 0.0003729253, 
    0.0003497193, 0.0003241609, 0.0002897015, 0.0002374242, 0.0001826356, 
    0.0001482715, 0.0001527696, 0.0001793135, 0.000188151, 0.0001862913, 
    0.000181205, 0.0001883576, 0.0001981168, 0.0001991659, 0.0001966704, 
    0.0001999129, 0.0002049673, 0.0002036004, 0.0001770883, 0.0001459827, 
    0.0001335689, 0.0001319795, 0.0001295636, 0.0001177698, 9.92367e-005, 
    9.310138e-005, 9.306963e-005, 7.43299e-005, 5.479547e-005, 4.145992e-005, 
    5.269737e-005, 9.796515e-005, 0.0001444885, 0.0001901537, 0.0002370903, 
    0.0002828825, 0.000334667, 0.000395289, 0.0004592011, 0.0005058675, 
    0.0005324113, 0.0005704949, 0.0005028475, 0.0004430839, 0.0003753889, 
    0.0003157366, 0.000266384, 0.0002481051, 0.0002673217, 0.0002944696, 
    0.0003211407, 0.000324145, 0.0003055006, 0.0002817541, 0.0002620767, 
    0.0002541612, 0.000251761, 0.0002566724, 0.0002540339, 0.000243019, 
    0.0002198447, 0.000200501, 0.0001864979, 0.0001846541, 0.0002182871, 
    0.0002101491, 0.0001849562, 0.0001183737, 8.731577e-005, 8.776085e-005, 
    0.0001313596, 0.0001964797, 0.0002162209, 0.0002413343, 0.0002539387, 
    0.0002818812, 0.000336956, 0.0003854821, 0.0003860227, 0.0006098021, 
    0.0008467266, 0.0007933208, 0.0006533531, 0.0003925709, 0.0002676712, 
    0.0002672735,
  0.0002826282, 0.0002425262, 0.0002459593, 0.0002262343, 6.741565e-005, 
    0.0003561884, 0.0003450464, 0.0003639609, 0.0004036975, 0.0004365833, 
    0.0004325301, 0.0005080294, 0.0004214515, 0.0003258138, 0.0002396652, 
    0.000205031, 0.0001863231, 0.0001790592, 0.0001755942, 0.000170953, 
    0.0001636892, 0.0001589367, 0.0001612891, 0.0001627991, 0.0001616706, 
    0.0001615593, 0.0001434236, 0.0001315663, 0.000125876, 0.0001227448, 
    0.0001230627, 0.0001166572, 0.0001030197, 8.548789e-005, 8.041752e-005, 
    8.095797e-005, 8.618737e-005, 9.044702e-005, 8.175272e-005, 
    7.951159e-005, 8.782445e-005, 0.0001088211, 0.0001442819, 0.0001720497, 
    0.0001976559, 0.0002090046, 0.0002275377, 0.0002582619, 0.0003009388, 
    0.000371606, 0.0004279841, 0.0004629045, 0.0004922934, 0.0003988018, 
    0.0003596693, 0.000315689, 0.0002895425, 0.0002787501, 0.0002764295, 
    0.000259152, 0.0002420813, 0.0002302875, 0.0002147425, 0.0001981963, 
    0.0001872131, 0.0001838116, 0.0001848289, 0.0001893748, 0.0001941114, 
    0.0002151717, 0.0001834143, 0.0001700629, 0.0001558532, 0.0001599858, 
    0.0001373519, 0.0001459668, 0.0001179605, 0.000107629, 0.000102368, 
    0.0001180241, 0.0001237938, 0.0001588414, 0.0001546293, 0.0001522769, 
    0.0001345544, 0.0001162757, 0.000118644, 0.0001515139, 0.0002106417, 
    0.0002861886, 0.0004098961, 0.0005408673, 0.0007689387, 0.00100758, 
    0.0007096678, 0.0004497436,
  0.0005546797, 0.0003908859, 0.0002884455, 0.0002437818, 0.0002025673, 
    0.0002424149, 0.0004154118, 0.000640288, 0.0009025007, 0.0010727, 
    0.001025159, 0.0008102646, 0.000583926, 0.0003868331, 0.0003004143, 
    0.0002111026, 0.0002047925, 0.0001893271, 0.0001806169, 0.0001548836, 
    0.000152563, 0.0001509099, 0.0001514345, 0.0001500516, 0.000140356, 
    0.0001282284, 0.0001154015, 0.0001050859, 0.0001018116, 0.0001016845, 
    0.0001044025, 0.000106278, 0.0001056264, 0.0001023521, 0.0001003017, 
    0.000111714, 0.0001135737, 0.0001098225, 9.823535e-005, 9.615318e-005, 
    0.0001035601, 0.0001143365, 0.0001313755, 0.0001503854, 0.0001680125, 
    0.0001822381, 0.0001937141, 0.0002072562, 0.0002244223, 0.0002364228, 
    0.0002433051, 0.0002411434, 0.0002307961, 0.0002153148, 0.00020999, 
    0.0002121358, 0.0002224196, 0.000233816, 0.0002421766, 0.000245435, 
    0.0002437979, 0.0002349287, 0.0002247084, 0.0001582691, 0.0001396725, 
    0.0001284191, 0.0001224905, 0.0001218547, 0.0001292457, 0.0001624335, 
    0.0001454105, 0.0001439323, 0.000145331, 0.0001171499, 0.0001060555, 
    9.987249e-005, 0.0001013825, 0.0001203288, 0.0001261939, 0.0001328378, 
    0.0001529286, 0.0001434395, 0.0001504808, 0.0001498768, 0.0001365254, 
    0.0001160214, 9.057418e-005, 7.111921e-005, 7.065825e-005, 9.22749e-005, 
    0.000133712, 0.0002187161, 0.0003202507, 0.000451381, 0.0005983422, 
    0.0007639319,
  0.0005414874, 0.0005543461, 0.0005206019, 0.0005902997, 0.0007527261, 
    0.0009471009, 0.0008119972, 0.0006693273, 0.000533858, 0.0004220397, 
    0.0003626256, 0.0003057549, 0.0002614725, 0.0002248832, 0.0001986731, 
    0.0001829375, 0.0001712073, 0.0001666138, 0.0001640389, 0.0001613209, 
    0.0001613527, 0.0001614322, 0.000159191, 0.0001598109, 0.0001635938, 
    0.0001292457, 0.0001211235, 0.0001076131, 0.0001000791, 9.440475e-005, 
    9.092383e-005, 9.407094e-005, 9.48657e-005, 0.0001006195, 0.0001078198, 
    0.0001147657, 0.0001205513, 0.0001245408, 0.0001268455, 0.000126925, 
    0.000126035, 0.0001266231, 0.0001274973, 0.0001278469, 0.0001280854, 
    0.0001278787, 0.0001278469, 0.0001304536, 0.0001343637, 0.000140356, 
    0.0001471588, 0.0001540889, 0.0001609235, 0.0001667092, 0.0001722722, 
    0.0001758485, 0.0001768976, 0.0001753081, 0.0001718908, 0.0001675516, 
    0.00016326, 0.0001601606, 0.0001596043, 0.0001586665, 0.0001643885, 
    0.0001279582, 0.0001212984, 0.0001147498, 0.0001082171, 0.0001041163, 
    0.0001017163, 9.992017e-005, 9.866449e-005, 9.89665e-005, 0.0001007785, 
    0.0001188347, 0.0001181036, 0.0001219024, 9.856913e-005, 9.130526e-005, 
    8.57581e-005, 8.108508e-005, 7.911419e-005, 8.081491e-005, 8.345341e-005, 
    8.304016e-005, 7.917777e-005, 7.533128e-005, 7.227952e-005, 
    7.552202e-005, 8.617138e-005, 0.0001067072, 0.0001458078, 0.0001953829, 
    0.0002697378, 0.0004097531,
  0.0002100696, 0.0002451011, 0.000283725, 0.0003665993, 0.0002431779, 
    0.0002303351, 0.0002103875, 0.0002163161, 0.0001915842, 0.0001729558, 
    0.0001624654, 0.0001554718, 0.0001519431, 0.0001525153, 0.0001547247, 
    0.0001575062, 0.0001590162, 0.0001575539, 0.0001536915, 0.0001474132, 
    0.0001401176, 0.0001339187, 0.0001302152, 0.0001316935, 0.0001427561, 
    0.0001116026, 0.0001142571, 0.0001386394, 0.0001340776, 0.0001300245, 
    0.0001239846, 0.0001185168, 0.0001121113, 0.0001053243, 9.903006e-005, 
    9.410275e-005, 9.059005e-005, 8.833304e-005, 8.788798e-005, 
    8.836482e-005, 8.912776e-005, 9.059005e-005, 9.2259e-005, 9.465906e-005, 
    9.790155e-005, 0.0001018434, 0.0001068979, 0.0001128742, 0.0001194546, 
    0.0001260826, 0.0001316775, 0.0001351584, 0.0001352855, 0.0001323927, 
    0.0001272906, 0.0001199314, 0.0001123338, 0.0001066595, 0.0001024951, 
    0.0001011759, 0.0001030355, 0.0001071681, 0.0001134941, 0.0001197725, 
    0.0001249223, 0.0001255263, 0.000123158, 0.0001184691, 0.0001100132, 
    0.0001037826, 0.0001028925, 7.440938e-005, 7.192983e-005, 7.056291e-005, 
    7.256561e-005, 7.558559e-005, 7.860555e-005, 7.954333e-005, 
    7.916185e-005, 7.657105e-005, 7.097616e-005, 6.476138e-005, 
    5.876913e-005, 5.387361e-005, 5.134636e-005, 5.09013e-005, 5.307887e-005, 
    5.633726e-005, 6.002479e-005, 6.472959e-005, 7.129404e-005, 
    8.153015e-005, 0.0001065642, 0.0001232375, 0.0001480012, 0.0001778036,
  0.0001059601, 0.0001092344, 0.0001120319, 0.0001142095, 0.0001135419, 
    0.0001142571, 0.0001151154, 0.0001144638, 0.0001134783, 0.0001138915, 
    0.0001152267, 0.0001164824, 0.000117293, 0.0001182149, 0.0001182944, 
    0.0001164029, 0.0001133987, 0.0001094728, 0.0001053084, 0.0001008897, 
    9.672536e-005, 9.30696e-005, 9.030393e-005, 8.836482e-005, 8.796745e-005, 
    8.846019e-005, 9.073308e-005, 9.283116e-005, 9.551736e-005, 
    9.828301e-005, 0.0001000632, 0.0001008103, 0.000100842, 9.958637e-005, 
    9.790155e-005, 9.543787e-005, 9.318086e-005, 9.100331e-005, 
    8.923902e-005, 8.78085e-005, 8.698199e-005, 8.677536e-005, 8.688663e-005, 
    8.741114e-005, 8.820587e-005, 8.939796e-005, 9.090794e-005, 9.24815e-005, 
    9.457959e-005, 9.640747e-005, 9.786976e-005, 9.850555e-005, 
    9.871217e-005, 9.877574e-005, 9.914133e-005, 9.953869e-005, 0.0001001745, 
    0.0001010487, 0.0001025587, 0.0001048475, 0.0001072953, 0.0001101881, 
    0.000112906, 0.0001148293, 0.0001152584, 0.0001144001, 0.0001120318, 
    0.0001087893, 0.0001048157, 0.0001006672, 9.802872e-005, 9.470675e-005, 
    9.402328e-005, 9.507235e-005, 9.724989e-005, 9.987249e-005, 0.0001027653, 
    0.0001048475, 0.0001073271, 0.0001093774, 0.0001096317, 0.0001089006, 
    0.0001076449, 0.0001049111, 0.0001010646, 9.767903e-005, 9.42617e-005, 
    9.219541e-005, 9.038342e-005, 9.01768e-005, 9.113047e-005, 9.422992e-005, 
    9.411866e-005, 9.532666e-005, 9.871217e-005, 0.0001025269,
  0.000109743, 0.0001101086, 0.0001107444, 0.000111253, 0.0001113484, 
    0.000111698, 0.0001119365, 0.0001116981, 0.0001116662, 0.0001115391, 
    0.0001112689, 0.0001105537, 0.0001099814, 0.0001088688, 0.0001072635, 
    0.0001059124, 0.0001039256, 0.0001022408, 0.0001008738, 9.964994e-005, 
    9.885522e-005, 9.763133e-005, 9.690018e-005, 9.59624e-005, 9.53743e-005, 
    9.527894e-005, 9.507232e-005, 9.494516e-005, 9.502465e-005, 
    9.494516e-005, 9.512001e-005, 9.548558e-005, 9.583526e-005, 
    9.586704e-005, 9.605778e-005, 9.623262e-005, 9.650284e-005, 
    9.662998e-005, 9.674125e-005, 9.677304e-005, 9.699557e-005, 
    9.728167e-005, 9.732936e-005, 9.740883e-005, 9.75042e-005, 9.736114e-005, 
    9.713862e-005, 9.701147e-005, 9.713863e-005, 9.702736e-005, 
    9.669358e-005, 9.624853e-005, 9.597832e-005, 9.554917e-005, 
    9.473855e-005, 9.399148e-005, 9.329212e-005, 9.299014e-005, 
    9.237024e-005, 9.171856e-005, 9.108278e-005, 8.997016e-005, 
    8.935027e-005, 8.930259e-005, 8.906416e-005, 8.919132e-005, 
    8.915953e-005, 8.890522e-005, 8.846018e-005, 8.852375e-005, 
    8.853964e-005, 8.831712e-005, 8.84125e-005, 8.885755e-005, 8.957281e-005, 
    9.000196e-005, 9.070132e-005, 9.148015e-005, 9.22272e-005, 9.322856e-005, 
    9.410275e-005, 9.51359e-005, 9.624853e-005, 9.712273e-005, 9.817177e-005, 
    9.909365e-005, 0.0001003334, 0.0001014937, 0.0001023997, 0.0001032739, 
    0.0001050382, 0.0001061508, 0.0001066277, 0.0001069933, 0.0001077085, 
    0.0001086304,
  1.789812e-005, 1.662656e-005, 1.53391e-005, 1.427416e-005, 1.327279e-005, 
    1.233501e-005, 1.142903e-005, 1.071377e-005, 1.010978e-005, 
    9.489886e-006, 9.013047e-006, 8.583893e-006, 8.202425e-006, 
    7.900428e-006, 7.662013e-006, 7.391802e-006, 7.216961e-006, 6.89907e-006, 
    6.819597e-006, 6.66065e-006, 6.581176e-006, 6.422231e-006, 6.454022e-006, 
    6.342758e-006, 6.342761e-006, 6.422233e-006, 6.581176e-006, 
    6.724229e-006, 6.835491e-006, 7.042119e-006, 7.344115e-006, 
    7.614326e-006, 8.011692e-006, 8.472634e-006, 9.028947e-006, 
    9.664735e-006, 1.031642e-005, 1.107936e-005, 1.195355e-005, 
    1.270061e-005, 1.371786e-005, 1.47828e-005, 1.580006e-005, 1.681731e-005, 
    1.794581e-005, 1.891539e-005, 1.998033e-005, 2.099756e-005, 
    2.190355e-005, 2.26506e-005, 2.333406e-005, 2.381091e-005, 2.41447e-005, 
    2.460564e-005, 2.451028e-005, 2.478048e-005, 2.476459e-005, 
    2.447849e-005, 2.392217e-005, 2.346124e-005, 2.311155e-005, 
    2.257113e-005, 2.199892e-005, 2.123597e-005, 2.074325e-005, 
    2.018696e-005, 1.97737e-005, 1.956706e-005, 1.955116e-005, 1.980548e-005, 
    2.028233e-005, 2.085453e-005, 2.1538e-005, 2.183999e-005, 2.306388e-005, 
    2.404935e-005, 2.490765e-005, 2.606795e-005, 2.726004e-005, 
    2.819782e-005, 2.921507e-005, 2.999391e-005, 3.051842e-005, 
    3.096347e-005, 3.097936e-005, 3.083632e-005, 3.040716e-005, 
    2.977138e-005, 2.886539e-005, 2.783226e-005, 2.656066e-005, 
    2.516194e-005, 2.373144e-005, 2.223735e-005, 2.067969e-005, 1.921739e-005,
  2.571826e-005, 2.230093e-005, 1.980549e-005, 1.82637e-005, 1.718287e-005, 
    1.673781e-005, 1.646761e-005, 1.664245e-005, 1.67855e-005, 1.689676e-005, 
    1.681729e-005, 1.664245e-005, 1.61815e-005, 1.545035e-005, 1.457615e-005, 
    1.3543e-005, 1.255754e-005, 1.141313e-005, 1.052303e-005, 9.696512e-006, 
    8.949468e-006, 8.488527e-006, 8.011689e-006, 7.677902e-006, 
    7.487169e-006, 7.280539e-006, 7.137489e-006, 7.185172e-006, 
    7.264645e-006, 7.3918e-006, 7.773277e-006, 8.266001e-006, 9.076626e-006, 
    1.010978e-005, 1.160386e-005, 1.355891e-005, 1.602258e-005, 
    1.888361e-005, 2.204662e-005, 2.527321e-005, 2.810243e-005, 
    3.055019e-005, 3.161514e-005, 3.279134e-005, 3.260063e-005, 
    3.094759e-005, 3.213968e-005, 3.23463e-005, 3.277544e-005, 3.374502e-005, 
    3.684443e-005, 4.10724e-005, 4.661962e-005, 5.321577e-005, 5.904908e-005, 
    6.66944e-005, 7.160581e-005, 7.470525e-005, 7.535695e-005, 7.275026e-005, 
    6.767991e-005, 6.052732e-005, 5.245293e-005, 4.364725e-005, 
    3.523912e-005, 2.8023e-005, 2.198304e-005, 1.702394e-005, 1.424241e-005, 
    1.324105e-005, 1.382912e-005, 1.562518e-005, 1.820009e-005, 
    2.123597e-005, 2.528907e-005, 2.951703e-005, 3.372911e-005, 
    3.789349e-005, 4.162871e-005, 4.572951e-005, 4.989388e-005, 
    5.192838e-005, 5.572723e-005, 5.690343e-005, 6.051148e-005, 
    6.195788e-005, 6.311819e-005, 6.318177e-005, 6.18943e-005, 5.917635e-005, 
    5.534575e-005, 5.057735e-005, 4.523678e-005, 3.970547e-005, 
    3.447617e-005, 2.977138e-005,
  1.70875e-005, 1.220787e-005, 9.060743e-006, 7.296436e-006, 6.46992e-006, 
    6.342758e-006, 6.835489e-006, 7.646115e-006, 8.758734e-006, 
    9.871355e-006, 1.09045e-005, 1.155618e-005, 1.185818e-005, 1.220785e-005, 
    1.231912e-005, 1.239859e-005, 1.233502e-005, 1.214428e-005, 
    1.174692e-005, 1.136545e-005, 1.115882e-005, 1.114292e-005, 
    1.125418e-005, 1.128597e-005, 1.112702e-005, 1.068198e-005, 
    1.023693e-005, 9.760094e-006, 9.473994e-006, 9.29915e-006, 9.330938e-006, 
    9.426305e-006, 9.760093e-006, 1.077734e-005, 1.23827e-005, 1.454437e-005, 
    1.785044e-005, 2.231682e-005, 2.791172e-005, 3.415827e-005, 
    3.997568e-005, 4.428311e-005, 4.736664e-005, 4.892434e-005, 4.87177e-005, 
    5.021179e-005, 5.045022e-005, 5.016412e-005, 4.995747e-005, 
    5.032305e-005, 5.149917e-005, 5.43443e-005, 5.951006e-005, 6.720304e-005, 
    7.677163e-005, 8.899462e-005, 9.931019e-005, 0.0001061924, 0.0001101184, 
    0.0001101025, 0.0001090694, 0.0001052229, 9.978685e-005, 9.416018e-005, 
    8.816796e-005, 8.222336e-005, 7.694637e-005, 7.174886e-005, 
    6.626526e-005, 5.9224e-005, 5.316819e-005, 4.711223e-005, 4.140618e-005, 
    3.848162e-005, 3.862467e-005, 4.008696e-005, 4.065917e-005, 4.29003e-005, 
    4.580902e-005, 4.968727e-005, 5.270723e-005, 5.585435e-005, 
    5.935116e-005, 6.197378e-005, 6.551819e-005, 6.94601e-005, 7.460991e-005, 
    8.047497e-005, 8.373335e-005, 8.460757e-005, 8.23983e-005, 7.392648e-005, 
    6.19897e-005, 4.868591e-005, 3.55252e-005, 2.487585e-005,
  1.223967e-005, 1.297082e-005, 1.707162e-005, 2.115652e-005, 2.373145e-005, 
    2.527322e-005, 2.481228e-005, 2.257113e-005, 1.978958e-005, 
    1.762791e-005, 1.605435e-005, 1.533909e-005, 1.56093e-005, 1.73577e-005, 
    2.045714e-005, 2.443079e-005, 2.919916e-005, 3.377681e-005, 
    3.700341e-005, 3.843393e-005, 3.649479e-005, 3.1488e-005, 2.581363e-005, 
    2.082273e-005, 1.67855e-005, 1.324101e-005, 1.131776e-005, 1.026872e-005, 
    9.807778e-006, 9.601152e-006, 9.617046e-006, 9.903144e-006, 
    1.066608e-005, 1.136544e-005, 1.209659e-005, 1.276417e-005, 
    1.344764e-005, 1.495762e-005, 1.746898e-005, 2.102937e-005, 
    2.482815e-005, 2.883358e-005, 3.344299e-005, 3.789351e-005, 
    4.180358e-005, 4.917866e-005, 8.271617e-005, 9.522517e-005, 0.0001122164, 
    0.0001257745, 0.0001356293, 0.0001437513, 0.0001529542, 0.0001640646, 
    0.000175461, 0.0001887965, 0.0002092211, 0.0001680542, 0.0001613625, 
    0.0001533199, 0.0001435606, 0.0001398731, 0.0001367896, 0.0001329272, 
    0.0001280317, 0.000119528, 0.0001087832, 9.814979e-005, 8.656262e-005, 
    7.379922e-005, 6.326113e-005, 5.466217e-005, 4.841559e-005, 
    4.668316e-005, 5.008461e-005, 5.547286e-005, 6.515271e-005, 
    7.645373e-005, 8.899454e-005, 0.0001019962, 0.000143799, 0.0001510628, 
    0.0001667666, 0.0001789577, 0.0001909423, 0.000201401, 0.0002072025, 
    0.0002100634, 0.0002329675, 0.0001555292, 0.0001320847, 0.0001029976, 
    7.441913e-005, 4.792296e-005, 2.795937e-005, 1.654709e-005,
  6.419902e-005, 4.631765e-005, 3.752792e-005, 3.485763e-005, 3.633583e-005, 
    3.941938e-005, 4.493478e-005, 5.342249e-005, 6.24347e-005, 6.725077e-005, 
    6.510501e-005, 5.677626e-005, 4.595205e-005, 3.633583e-005, 
    3.148799e-005, 3.110653e-005, 3.436491e-005, 3.922865e-005, 4.3393e-005, 
    4.503015e-005, 5.097472e-005, 5.030715e-005, 4.035715e-005, 
    2.894486e-005, 2.091809e-005, 1.538678e-005, 1.413112e-005, 
    1.489405e-005, 1.678551e-005, 1.831138e-005, 1.792991e-005, 
    1.632457e-005, 1.583184e-005, 1.6865e-005, 1.827959e-005, 1.996442e-005, 
    2.044124e-005, 1.950347e-005, 1.851801e-005, 1.921738e-005, 
    2.168102e-005, 2.541624e-005, 3.013694e-005, 3.358607e-005, 
    3.856109e-005, 4.743024e-005, 8.835871e-005, 0.0001342783, 0.0001602976, 
    0.0001465648, 0.0001229454, 0.000119544, 0.0001440851, 0.0001969028, 
    0.0002585737, 0.0003115503, 0.000353989, 0.0003818999, 0.0004101761, 
    0.0004364817, 0.0004633436, 0.0004919061, 0.0005041448, 0.0005073556, 
    0.0004972942, 0.0004762976, 0.0004535365, 0.0004384685, 0.0004172175, 
    0.0003951557, 0.0003204671, 0.0003980804, 0.0004085233, 0.0004043906, 
    0.0003873676, 0.0003593453, 0.0003021884, 0.0002848792, 0.0002669978, 
    0.0002499588, 0.0002575088, 0.0002353517, 0.0002360193, 0.0002534874, 
    0.0002836553, 0.0003217388, 0.000353814, 0.0003726014, 0.0003794837, 
    0.0003773539, 0.000387272, 0.0002679992, 0.0002310126, 0.0001872547, 
    0.0001372027, 9.443043e-005,
  0.0009521018, 0.0007107744, 0.0003068773, 0.0002213645, 0.0001674184, 
    0.0001422572, 0.0001405565, 0.000162491, 0.0001983492, 0.0002332536, 
    0.0002477336, 0.0002314894, 0.0001891939, 0.0001383789, 9.520934e-005, 
    6.764814e-005, 5.31046e-005, 4.871769e-005, 5.369274e-005, 6.224395e-005, 
    7.119257e-005, 8.35268e-005, 8.311353e-005, 7.112895e-005, 5.704648e-005, 
    4.75892e-005, 4.291619e-005, 4.386986e-005, 5.107e-005, 5.944652e-005, 
    6.111542e-005, 6.000284e-005, 5.800014e-005, 5.827037e-005, 
    6.197381e-005, 6.671034e-005, 6.855412e-005, 6.335662e-005, 
    5.537752e-005, 4.981444e-005, 4.90197e-005, 5.108598e-005, 5.588619e-005, 
    6.040011e-005, 0.0001236289, 0.000188717, 0.0001985399, 0.0001693894, 
    6.740959e-005, -2.225162e-005, -8.726073e-005, -0.0001024082, 
    -7.150904e-005, -2.180715e-005, 3.202772e-005, 7.638964e-005, 
    0.0001288576, 0.000185617, 0.0002619904, 0.0003527643, 0.000433191, 
    0.0005095962, 0.0005702497, 0.000608206, 0.000612132, 0.0005912783, 
    0.0005694868, 0.0005609356, 0.0005901817, 0.0006762031, 0.0007714911, 
    0.0008144225, 0.0008131033, 0.0008070315, 0.0007932826, 0.0007420704, 
    0.0006761079, 0.0006280114, 0.0004719426, 0.0004593859, 0.0004775218, 
    0.0004683504, 0.0004666657, 0.0004767111, 0.0005122196, 0.0005755594, 
    0.0006465446, 0.0006922415, 0.000723983, 0.0007768165, 0.0008795114, 
    0.001028301, 0.001169794, 0.001259424, 0.001244705, 0.001140612,
  0.001374341, 0.001363707, 0.001330313, 0.00128274, 0.0012376, 0.001197164, 
    0.001149226, 0.001097425, 0.00103968, 0.0009969398, 0.0009850349, 
    0.0009853526, 0.0009960337, 0.001032496, 0.001073806, 0.001099841, 
    0.001079147, 0.001019829, 0.0009578398, 0.0009135891, 0.0008804646, 
    0.0008155989, 0.0007431197, 0.0006678591, 0.0005732072, 0.0004415838, 
    0.0003349949, 0.0002675226, 0.0002014327, 0.0001765257, 0.0001863008, 
    0.0002379103, 0.000328367, 0.00028809, 0.000330608, 0.0003917068, 
    0.0007350136, 0.0006117828, 0.0005348211, 0.0005379519, 0.0005494282, 
    0.0005208182, 0.0004620554, 0.0003794038, 0.0003012819, 0.0001778286, 
    7.006363e-005, 2.84519e-006, -4.323293e-005, -7.100124e-005, 
    -7.026992e-005, -4.723854e-005, -2.776785e-005, -2.234778e-005, 
    -2.640043e-005, -2.085348e-005, 1.896243e-005, 8.228631e-005, 
    0.0001414777, 0.0001908939, 0.000232792, 0.0002848469, 0.0003451188, 
    0.000404882, 0.0004426001, 0.0004545527, 0.0004568417, 0.0004591621, 
    0.0004709561, 0.0004953223, 0.0005279381, 0.0005728242, 0.0005971587, 
    0.0006074265, 0.0006041205, 0.0005716481, 0.000516224, 0.0004643439, 
    0.0005099298, 0.0007395272, 0.0007696473, 0.0007571385, 0.0007654515, 
    0.0007689481, 0.0008193657, 0.0008751876, 0.0009646262, 0.001023865, 
    0.00105904, 0.001086426, 0.001122014, 0.001174228, 0.001234357, 
    0.001298476, 0.001337545, 0.001361196,
  0.0006085555, 0.0006015936, 0.0006041049, 0.0006107173, 0.0006171227, 
    0.0006216688, 0.0006207628, 0.0006120042, 0.000597588, 0.0005856671, 
    0.0005820908, 0.0005867637, 0.0005982872, 0.0006151195, 0.0006408214, 
    0.0006564299, 0.000666793, 0.0006612781, 0.0006400587, 0.0005960623, 
    0.0005467255, 0.0004964669, 0.0004387696, 0.0003887655, 0.0003414312, 
    0.0002973399, 0.0002443632, 0.0001863637, 0.0001416525, 0.0001176996, 
    0.0001049999, 0.0001091165, 0.0001268866, 0.0001694206, 0.0002309959, 
    0.0002872946, 0.0003221512, 0.0003408594, 0.0003568013, 0.0003917054, 
    0.0004313623, 0.0004347956, 0.0004140059, 0.0003971416, 0.0003675781, 
    0.000286913, 0.0001617908, 5.552033e-005, 6.739516e-006, -1.73091e-005, 
    -3.531761e-005, -5.405815e-005, -8.098315e-005, -0.0001037749, 
    -9.919796e-005, -6.484985e-005, -1.525879e-005, 4.121428e-005, 
    7.271813e-005, 9.024981e-005, 0.0001256154, 0.000202179, 0.0002839407, 
    0.0003475659, 0.0004054704, 0.0004553157, 0.0005028723, 0.0005496508, 
    0.0005787215, 0.0005809776, 0.0005802624, 0.000597652, 0.0006304588, 
    0.0006688442, 0.0007004733, 0.0007094061, 0.0006837682, 0.0006268974, 
    0.0005573747, 0.0005437688, 0.0005979217, 0.0006080468, 0.0005239965, 
    0.0004337314, 0.0004450958, 0.0004856908, 0.0005274934, 0.0005590441, 
    0.0005921205, 0.0006227016, 0.0006299973, 0.0006205242, 0.000616455, 
    0.0006192047, 0.000625642, 0.0006241957,
  0.0004472572, 0.000452677, 0.0004479564, 0.0004393256, 0.0004336676, 
    0.0004353682, 0.0004402159, 0.0004475117, 0.0004531699, 0.0004668869, 
    0.0004827501, 0.0005034609, 0.0005199271, 0.0005364101, 0.0005547209, 
    0.000569439, 0.0005697412, 0.0005551819, 0.0005406383, 0.0005211667, 
    0.0004795869, 0.0004391985, 0.0004033246, 0.0003979201, 0.0003953939, 
    0.0003744122, 0.0003448008, 0.0003145691, 0.0002842741, 0.0002821758, 
    0.0002813023, 0.0002505458, 0.0002088863, 0.000185506, 0.0001871907, 
    0.0001954553, 0.0001974585, 0.000204436, 0.0002503553, 0.0003153961, 
    0.0003639702, 0.0004151352, 0.0004661405, 0.0004910314, 0.0004830691, 
    0.0004671584, 0.0004155319, 0.0003219447, 0.0002119862, 0.0001079086, 
    4.550675e-005, -6.516464e-006, -5.593244e-005, -8.053752e-005, 
    -9.245845e-005, -9.128219e-005, -5.214987e-005, 2.090167e-005, 
    7.683458e-005, 0.0001031877, 0.0001405249, 0.0002033086, 0.0002616737, 
    0.0003048112, 0.0003868593, 0.0004849122, 0.0005506203, 0.0005967459, 
    0.000647482, 0.0006827042, 0.0007064352, 0.0007209624, 0.0007382557, 
    0.0007645292, 0.0007891026, 0.0007876083, 0.0007478562, 0.0007317546, 
    0.0007161144, 0.0006979629, 0.0006886325, 0.000667477, 0.0005988432, 
    0.0004626112, 0.0004267218, 0.0004120674, 0.0004259432, 0.0004437761, 
    0.0004505471, 0.0004695414, 0.0004923819, 0.000502618, 0.0005113124, 
    0.0005123452, 0.0004919206, 0.0004631516,
  0.0004472411, 0.0004675542, 0.0004906491, 0.0004962119, 0.000488678, 
    0.0004934464, 0.0005002809, 0.0005100719, 0.0005281442, 0.0005440395, 
    0.0005563423, 0.0005761627, 0.0005966509, 0.0006060922, 0.0006275657, 
    0.0006684628, 0.0007282738, 0.0007700925, 0.0007446134, 0.0006668731, 
    0.0006047091, 0.000563669, 0.0005194186, 0.0005038427, 0.0005032388, 
    0.0004955614, 0.0004954343, 0.0004924936, 0.0004735156, 0.0004360201, 
    0.0004065358, 0.0003760029, 0.0003586616, 0.0003559124, 0.0003496967, 
    0.0003237091, 0.0003148876, 0.0003320859, 0.0003847131, 0.0004388969, 
    0.0004922552, 0.0005475529, 0.0005928362, 0.0005917079, 0.0005798666, 
    0.0005498258, 0.0004832591, 0.0004203324, 0.0003302582, 0.0002277535, 
    0.0001799273, 0.0001465483, 9.501819e-005, 7.128762e-005, 7.565878e-005, 
    6.338814e-005, 7.81063e-005, 0.0001479792, 0.000230615, 0.000266314, 
    0.000296291, 0.0003369339, 0.0003556418, 0.0004024352, 0.0005272869, 
    0.0006391848, 0.0006594188, 0.0006673657, 0.000715733, 0.000777706, 
    0.0008147722, 0.0008166479, 0.0007947609, 0.0007800898, 0.0007724292, 
    0.0007432308, 0.0007659919, 0.0008374215, 0.0008405689, 0.0007359195, 
    0.0006901906, 0.0006607533, 0.0006430629, 0.0005618581, 0.0004693042, 
    0.0004656324, 0.0005271281, 0.0005730316, 0.0005755266, 0.0005551185, 
    0.0005456759, 0.0005405103, 0.0005214848, 0.0004821774, 0.0004498637, 
    0.0004374501,
  0.0006223363, 0.0006094305, 0.0006450973, 0.0006883629, 0.0007003634, 
    0.000708438, 0.0007308652, 0.0007543731, 0.0007727942, 0.0007949355, 
    0.0007994971, 0.0008193976, 0.0008386457, 0.0008313661, 0.0008444311, 
    0.0008845017, 0.0009535793, 0.0009994037, 0.000966534, 0.0009023361, 
    0.0009044497, 0.0009344588, 0.0009090272, 0.0008577672, 0.0008097813, 
    0.0007745274, 0.0007547066, 0.00073638, 0.000699902, 0.0006499295, 
    0.0005964604, 0.000561222, 0.0005452638, 0.0005559768, 0.000550366, 
    0.0005266513, 0.0005212468, 0.000555357, 0.000601308, 0.0006651883, 
    0.0007428485, 0.0007793107, 0.0007605869, 0.0007487135, 0.0007869569, 
    0.0007462818, 0.0006302674, 0.0005581863, 0.0004966259, 0.0004363218, 
    0.0004244805, 0.0004314901, 0.0003877324, 0.0003585657, 0.0003712019, 
    0.0003698189, 0.0003786087, 0.0004358133, 0.0004847688, 0.0004899981, 
    0.0005414803, 0.0006117821, 0.0006248001, 0.0006451444, 0.0007175445, 
    0.0007616519, 0.0007923283, 0.0008295695, 0.0008760137, 0.0009023664, 
    0.0009062611, 0.0009010318, 0.0008859956, 0.0008612638, 0.0008382169, 
    0.0008346401, 0.0007973039, 0.0007899925, 0.0008389475, 0.0008504875, 
    0.0007303557, 0.0006256108, 0.0006145481, 0.0005474887, 0.0005324683, 
    0.0006332877, 0.00069782, 0.000719659, 0.0007300698, 0.000732136, 
    0.0007425789, 0.000737159, 0.0007008561, 0.0006671278, 0.0006584176, 
    0.0006453046,
  0.0008807662, 0.0008996492, 0.0009462992, 0.0009844145, 0.001025168, 
    0.00110631, 0.00121665, 0.001272107, 0.001252652, 0.001271582, 
    0.00132521, 0.001351723, 0.001333873, 0.001320998, 0.001331631, 
    0.001357111, 0.001413377, 0.001458884, 0.001461586, 0.001564614, 
    0.00171086, 0.001709366, 0.001535766, 0.001300638, 0.00112451, 
    0.001032066, 0.0009889286, 0.000935602, 0.0008846442, 0.0008430323, 
    0.0007971763, 0.0007615094, 0.0007583303, 0.0007546269, 0.0007620337, 
    0.0008023265, 0.0008428572, 0.0008726278, 0.0009022234, 0.0009598895, 
    0.001071437, 0.001128926, 0.001119453, 0.001133456, 0.001229715, 
    0.001158349, 0.001058594, 0.0009505595, 0.0008852961, 0.0008350057, 
    0.0008554142, 0.0008975817, 0.0008580685, 0.0007765442, 0.0007199449, 
    0.0006932253, 0.0006840862, 0.0007217093, 0.0007456141, 0.0007362524, 
    0.0007352033, 0.000732041, 0.0007304666, 0.0007965094, 0.0008921623, 
    0.0009523071, 0.001001866, 0.001033798, 0.001046816, 0.001041825, 
    0.001021401, 0.000991106, 0.0009677727, 0.0009591421, 0.0009584096, 
    0.0009417683, 0.0008492316, 0.0007398929, 0.00078524, 0.0009741932, 
    0.0008821329, 0.0006945776, 0.0005989717, 0.0005458351, 0.0006446368, 
    0.0008294103, 0.0009462195, 0.0009696013, 0.0009670579, 0.0009500827, 
    0.0009480962, 0.0009358404, 0.000896486, 0.0008825939, 0.0008966927, 
    0.0008888724,
  0.001434993, 0.001373385, 0.001341104, 0.001396481, 0.00152122, 
    0.001726229, 0.00197989, 0.002117967, 0.002190621, 0.002264388, 
    0.00234607, 0.002279726, 0.00208133, 0.001922226, 0.001876385, 
    0.001890086, 0.00192329, 0.001937309, 0.001957924, 0.002002047, 
    0.001959307, 0.001771131, 0.001488701, 0.001260597, 0.001148843, 
    0.001129707, 0.00114371, 0.001121871, 0.00108366, 0.001075632, 
    0.001078175, 0.001083341, 0.001104943, 0.001091067, 0.001078701, 
    0.001122268, 0.001152738, 0.001148477, 0.001162957, 0.001298442, 
    0.001538085, 0.001636027, 0.001618305, 0.001628334, 0.001702737, 
    0.001781606, 0.00158518, 0.00160845, 0.001600184, 0.001607974, 
    0.001590887, 0.001497443, 0.001350752, 0.001194412, 0.001088269, 
    0.001028823, 0.00101493, 0.0010317, 0.001042984, 0.001041507, 
    0.001018237, 0.001017999, 0.001033512, 0.001070037, 0.001112143, 
    0.001169283, 0.001209782, 0.001228968, 0.001204378, 0.001198259, 
    0.001211642, 0.001186354, 0.001126145, 0.001046784, 0.0009684553, 
    0.000920088, 0.0008565262, 0.000530879, 0.0005356474, 0.001076952, 
    0.001051123, 0.0009584893, 0.0009945389, 0.001074838, 0.001101605, 
    0.00113406, 0.001217238, 0.001268324, 0.001278369, 0.001280084, 
    0.001309648, 0.001325082, 0.001299238, 0.00132451, 0.001406558, 
    0.001444593,
  0.001534524, 0.001446611, 0.001427411, 0.001558382, 0.001786646, 
    0.002020012, 0.002155083, 0.002406822, 0.002467236, 0.002350697, 
    0.002141779, 0.001920098, 0.00172512, 0.001637127, 0.001617274, 
    0.001681235, 0.001818006, 0.001881124, 0.001865004, 0.001808945, 
    0.001716343, 0.00162336, 0.001504564, 0.001435708, 0.001432482, 
    0.00142525, 0.001393524, 0.001341501, 0.001308297, 0.001358206, 
    0.001335287, 0.001307916, 0.001286839, 0.001251458, 0.001303274, 
    0.001372877, 0.001354852, 0.001411881, 0.001495519, 0.001471646, 
    0.00200383, 0.002295384, 0.002287436, 0.002140746, 0.002130113, 
    0.002170278, 0.002162473, 0.001798962, 0.001889898, 0.001859079, 
    0.001706967, 0.001626588, 0.001531218, 0.00144588, 0.001443941, 
    0.001423278, 0.001391887, 0.001377709, 0.001348828, 0.001327689, 
    0.00131874, 0.001316578, 0.001366504, 0.001387007, 0.001426332, 
    0.001480057, 0.00148635, 0.001472745, 0.001421008, 0.001359147, 
    0.001298398, 0.001182209, 0.00102935, 0.0008816402, 0.0007997826, 
    0.0007432615, 0.0005630171, 0.000353639, 0.0007107262, 0.001125208, 
    0.00121692, 0.001329281, 0.001656058, 0.001822934, 0.0017444, 
    0.001669631, 0.001706634, 0.001716218, 0.001693315, 0.001656152, 
    0.001630514, 0.001632786, 0.001606482, 0.001593477, 0.001606511, 
    0.00159788,
  0.001519682, 0.00146262, 0.001453179, 0.00151315, 0.001664848, 0.001907271, 
    0.002193612, 0.002201591, 0.002117794, 0.002153193, 0.001770626, 
    0.001798728, 0.001747531, 0.001692473, 0.001689405, 0.001777316, 
    0.001876118, 0.001902931, 0.001904569, 0.001870667, 0.001840132, 
    0.001854104, 0.001835141, 0.001789572, 0.001721924, 0.00165423, 
    0.001635171, 0.001630038, 0.001628735, 0.001563312, 0.00143436, 
    0.001471569, 0.001445089, 0.0014198, 0.001526787, 0.001533463, 
    0.001544716, 0.001753281, 0.001897271, 0.001973024, 0.002269553, 
    0.002628995, 0.002752768, 0.002563685, 0.00241852, 0.002365289, 
    0.002245396, 0.002086912, 0.001897464, 0.001736373, 0.001727647, 
    0.001766398, 0.001806563, 0.00181858, 0.001872685, 0.001847365, 
    0.001772104, 0.001702533, 0.001602874, 0.001619945, 0.001661255, 
    0.001696637, 0.001767559, 0.001781769, 0.001784932, 0.001730429, 
    0.001666931, 0.001589729, 0.00141535, 0.001266736, 0.00107438, 
    0.0008713109, 0.0008126767, 0.0007748641, 0.0006597703, 0.0005806154, 
    0.0005329922, 0.0008622962, 0.001276095, 0.001494009, 0.001687322, 
    0.002113345, 0.002341622, 0.002383091, 0.002257587, 0.002098039, 
    0.002060065, 0.00194607, 0.001875182, 0.001882747, 0.001857061, 
    0.001835125, 0.001797314, 0.001754922, 0.001665769, 0.001588585,
  0.001374548, 0.001343205, 0.001297062, 0.001519269, 0.001839575, 
    0.002026827, 0.002239973, 0.002330192, 0.00246355, 0.002280636, 
    0.002141478, 0.002158707, 0.002188733, 0.002069873, 0.00203074, 
    0.002143544, 0.002263453, 0.002324631, 0.002344532, 0.002330529, 
    0.002311724, 0.002258955, 0.002163333, 0.002113202, 0.002032251, 
    0.001907066, 0.001885211, 0.001827481, 0.001765539, 0.001767511, 
    0.001797329, 0.002002654, 0.002240307, 0.002088101, 0.001973326, 
    0.002005751, 0.00210142, 0.002276531, 0.002395566, 0.002644745, 
    0.002697437, 0.002695118, 0.00233795, 0.002307639, 0.002331529, 
    0.002300916, 0.002215245, 0.002095717, 0.002097243, 0.002203546, 
    0.002292889, 0.002367944, 0.002409365, 0.002294304, 0.002201098, 
    0.002145085, 0.00205676, 0.001967782, 0.001851862, 0.001905952, 
    0.001988684, 0.00205552, 0.00210589, 0.002067441, 0.002013335, 
    0.001878423, 0.00178156, 0.001620136, 0.001398088, 0.001158367, 
    0.0008739969, 0.0007952871, 0.0007177861, 0.0006425567, 0.0005268119, 
    0.0006164107, 0.0008606138, 0.001024229, 0.001647138, 0.00206388, 
    0.002292047, 0.002626723, 0.002643539, 0.002690063, 0.002631284, 
    0.002370279, 0.002325696, 0.002306066, 0.002231266, 0.002173902, 
    0.002140841, 0.002036144, 0.001888659, 0.001745575, 0.001598328, 
    0.001463987,
  0.001405512, 0.001389919, 0.001545955, 0.001905173, 0.002219314, 
    0.002002667, 0.002053149, 0.002262577, 0.00230721, 0.00236176, 
    0.002342101, 0.002400942, 0.002430458, 0.002362859, 0.002385556, 
    0.002584222, 0.00275782, 0.00287781, 0.002861264, 0.002720676, 
    0.002596094, 0.002483068, 0.002365877, 0.002262276, 0.002141733, 
    0.002043789, 0.002058555, 0.002039816, 0.002129032, 0.002378642, 
    0.00260997, 0.002859943, 0.002812957, 0.002414607, 0.001863321, 
    0.002186584, 0.002120827, 0.002366732, 0.002835989, 0.002877713, 
    0.002785509, 0.002564273, 0.002392786, 0.002565115, 0.002603421, 
    0.002649517, 0.002673644, 0.002700632, 0.002782109, 0.00285346, 
    0.002830778, 0.002800291, 0.002822973, 0.002652789, 0.002479571, 
    0.002458352, 0.002275643, 0.002209029, 0.002191864, 0.002267648, 
    0.002302935, 0.002265058, 0.002194867, 0.002072098, 0.001997996, 
    0.001768799, 0.00157161, 0.001300893, 0.001166871, 0.001060233, 
    0.0008678772, 0.0008916389, 0.0006671762, 0.0006297128, 0.0006054109, 
    0.0008467538, 0.001341822, 0.000670386, 0.001800472, 0.002634147, 
    0.002777498, 0.002790024, 0.002673024, 0.002814502, 0.002912367, 
    0.00265168, 0.002501887, 0.002443348, 0.002385762, 0.002245492, 
    0.002108258, 0.001977828, 0.001807152, 0.001617163, 0.001507554, 
    0.001411869,
  0.001661525, 0.001727981, 0.002144609, 0.00261016, 0.00196438, 0.002091677, 
    0.002156656, 0.002546026, 0.002699855, 0.002426659, 0.002529876, 
    0.002687296, 0.002544787, 0.002703527, 0.002829077, 0.002936684, 
    0.002950607, 0.00295477, 0.002837835, 0.002678733, 0.002541689, 
    0.002523618, 0.002488155, 0.002395283, 0.002318686, 0.002306813, 
    0.002357487, 0.002521694, 0.002764722, 0.003159732, 0.003445581, 
    0.003159271, 0.0027582, 0.001840846, 0.001645518, 0.002084255, 
    0.002070555, 0.002531624, 0.003014932, 0.003001915, 0.00307673, 
    0.002865429, 0.003065065, 0.003195417, 0.003168555, 0.003170589, 
    0.003247853, 0.003221706, 0.003200214, 0.003160877, 0.003159367, 
    0.003079494, 0.003029253, 0.002919214, 0.00285295, 0.00281536, 
    0.002623798, 0.002593631, 0.002544755, 0.002513109, 0.002375621, 
    0.002227724, 0.002121421, 0.001949472, 0.001805929, 0.001512704, 
    0.001327677, 0.00120888, 0.001139992, 0.001085125, 0.0009621158, 
    0.0008912263, 0.0007752283, 0.0008830251, 0.0008498216, 0.001310685, 
    0.002027482, 0.0008571791, 0.001679501, 0.002884899, 0.003076874, 
    0.00280684, 0.002771872, 0.002601387, 0.002691, 0.002693163, 0.002544215, 
    0.002405092, 0.002314109, 0.002203882, 0.00202311, 0.001855582, 
    0.001718586, 0.001583673, 0.001601395, 0.001594116,
  0.002195727, 0.002271734, 0.00261827, 0.002785275, 0.002319274, 
    0.002156863, 0.002577244, 0.002792996, 0.002512315, 0.002420858, 
    0.002807796, 0.002954582, 0.0026742, 0.002636942, 0.002966123, 
    0.003022293, 0.002969254, 0.002961449, 0.002879621, 0.002861088, 
    0.002822321, 0.002851456, 0.002763256, 0.002689015, 0.002710711, 
    0.002812292, 0.002952101, 0.003167901, 0.003390824, 0.003773628, 
    0.004130429, 0.003754236, 0.002898425, 0.001265256, 0.001739836, 
    0.002026748, 0.002513869, 0.003078383, 0.00336369, 0.003126734, 
    0.003113128, 0.003314704, 0.003434468, 0.003443591, 0.003450682, 
    0.00342932, 0.00341427, 0.003319267, 0.003300019, 0.003315039, 
    0.003345668, 0.003215218, 0.003114128, 0.003046766, 0.00302108, 
    0.002955293, 0.002859259, 0.002795728, 0.002696946, 0.002585398, 
    0.002381645, 0.002208538, 0.00210125, 0.001906093, 0.001741255, 
    0.001550583, 0.001448872, 0.001369525, 0.001312243, 0.0012558, 
    0.001199502, 0.001189425, 0.00120559, 0.001259646, 0.00129258, 
    0.001876913, 0.002300312, 0.001580921, 0.002330843, 0.003099237, 
    0.003181525, 0.003025473, 0.003181365, 0.002493606, 0.002276263, 
    0.00264392, 0.002528351, 0.002522122, 0.002361586, 0.002228105, 
    0.00209971, 0.002019394, 0.002024513, 0.001990527, 0.002089867, 
    0.002064008,
  0.002673693, 0.002681609, 0.002848119, 0.002840299, 0.002364559, 
    0.001978033, 0.002554054, 0.002453217, 0.002634575, 0.00246665, 
    0.002662724, 0.0031607, 0.002912128, 0.002777612, 0.002965752, 
    0.002996285, 0.002998384, 0.003104862, 0.003119374, 0.003150687, 
    0.003107978, 0.003117545, 0.00311836, 0.003220098, 0.003238317, 
    0.003288573, 0.00342172, 0.003556315, 0.003678434, 0.003771719, 
    0.004054133, 0.004140105, 0.003833152, 0.003546845, 0.003266958, 
    0.002834879, 0.002917306, 0.003489928, 0.003332984, 0.003282374, 
    0.003403857, 0.00348247, 0.0035419, 0.003501272, 0.003583018, 
    0.003584433, 0.003497284, 0.003352134, 0.003274934, 0.003179949, 
    0.003129005, 0.003077062, 0.002963368, 0.002883879, 0.002891541, 
    0.002902016, 0.002894528, 0.002842713, 0.002798922, 0.00267493, 
    0.002529908, 0.00245546, 0.002374699, 0.002204308, 0.002067363, 
    0.001992801, 0.001932355, 0.001872811, 0.001810028, 0.001745082, 
    0.001771516, 0.001761151, 0.001759261, 0.001777793, 0.001977763, 
    0.002419254, 0.001985568, 0.002355656, 0.002480254, 0.003182796, 
    0.00320689, 0.002916309, 0.002736078, 0.002572061, 0.002412989, 
    0.002522616, 0.002540544, 0.002535267, 0.002453728, 0.002454124, 
    0.002436737, 0.00247431, 0.00259619, 0.00258602, 0.002704322, 0.002623564,
  0.003031733, 0.003011629, 0.003053648, 0.003144456, 0.002721534, 
    0.001736166, 0.002192372, 0.00220949, 0.002287342, 0.002353925, 
    0.002485721, 0.003174512, 0.003393602, 0.003118133, 0.003064077, 
    0.003015153, 0.003118865, 0.003257576, 0.003283929, 0.003357299, 
    0.003389612, 0.003402201, 0.003392966, 0.003532346, 0.003554121, 
    0.003631052, 0.003652383, 0.003531408, 0.003465859, 0.003358619, 
    0.003419129, 0.003619814, 0.003787771, 0.003597958, 0.003624089, 
    0.003142565, 0.003270755, 0.003494661, 0.00327651, 0.003191249, 
    0.003344519, 0.003483439, 0.003440903, 0.003292527, 0.003253348, 
    0.003264396, 0.003268225, 0.003191343, 0.003140369, 0.003069084, 
    0.003006332, 0.00295496, 0.002837149, 0.002773762, 0.002832444, 
    0.002867095, 0.002900474, 0.002960555, 0.002988562, 0.00291883, 
    0.002863232, 0.002784461, 0.002730595, 0.002709171, 0.002597954, 
    0.002516557, 0.002439821, 0.002361318, 0.002366785, 0.002425611, 
    0.002442524, 0.002357026, 0.00232242, 0.002458053, 0.002813548, 
    0.003179919, 0.002835577, 0.002390544, 0.002558457, 0.002952103, 
    0.002805106, 0.002210793, 0.002551719, 0.00265179, 0.002019996, 
    0.002410416, 0.002685245, 0.002826231, 0.002846098, 0.002940416, 
    0.003018161, 0.003101144, 0.003155218, 0.003101399, 0.003180934, 
    0.003094833,
  0.003208224, 0.003153292, 0.003059832, 0.003107835, 0.003298061, 
    0.003054397, 0.003179077, 0.002978835, 0.002764784, 0.002743913, 
    0.00286872, 0.003161207, 0.003211182, 0.003090905, 0.003185544, 
    0.003136411, 0.003318485, 0.003358603, 0.003355503, 0.003270229, 
    0.00334549, 0.003429508, 0.003431194, 0.003526593, 0.003481038, 
    0.003462458, 0.003408685, 0.003286839, 0.003197003, 0.003261423, 
    0.003334252, 0.003290016, 0.003336383, 0.003339354, 0.003351418, 
    0.003236182, 0.003120374, 0.003231781, 0.002935492, 0.002918467, 
    0.003219923, 0.003297059, 0.003252937, 0.003238296, 0.003156424, 
    0.003026884, 0.003068956, 0.003061643, 0.003057066, 0.003061486, 
    0.003017981, 0.002959998, 0.002912205, 0.00280579, 0.0028855, 
    0.002840266, 0.002824927, 0.002892558, 0.002879189, 0.002875168, 
    0.00288666, 0.002859354, 0.002873324, 0.002849041, 0.002870454, 
    0.002882533, 0.002867462, 0.002881497, 0.002878875, 0.002939465, 
    0.00295029, 0.002956774, 0.003033036, 0.003163962, 0.003148401, 
    0.002993636, 0.002273609, 0.002004197, 0.00240989, 0.002992839, 
    0.002527226, 0.002373205, 0.002342992, 0.002667492, 0.002586829, 
    0.00228682, 0.002569709, 0.003029745, 0.003079224, 0.003157727, 
    0.003286934, 0.00335981, 0.003389295, 0.003414251, 0.003358128, 
    0.003280384,
  0.003151322, 0.003094068, 0.003075313, 0.00289523, 0.003134873, 
    0.003263731, 0.003711035, 0.003224712, 0.003001836, 0.002899093, 
    0.002715353, 0.00307234, 0.003219588, 0.003260311, 0.003324637, 
    0.003351832, 0.003444511, 0.003498316, 0.003585799, 0.003459325, 
    0.003525097, 0.003565598, 0.003590409, 0.003597593, 0.003577773, 
    0.003453683, 0.003325684, 0.003293451, 0.003259091, 0.00331332, 
    0.003260899, 0.003425788, 0.003461441, 0.003208844, 0.003125302, 
    0.003199751, 0.003098583, 0.002816062, 0.002527365, 0.002749857, 
    0.003113827, 0.00316062, 0.003203455, 0.003212675, 0.003099363, 
    0.00293587, 0.002982616, 0.002972476, 0.002986128, 0.002944501, 
    0.00289863, 0.002961285, 0.00301571, 0.002990786, 0.003075887, 
    0.003075471, 0.003083643, 0.003087236, 0.003043985, 0.002998289, 
    0.003010195, 0.003051313, 0.003042681, 0.002985494, 0.003043907, 
    0.003069703, 0.003114669, 0.003175229, 0.00316493, 0.003192969, 
    0.003177822, 0.003182428, 0.003200499, 0.003208812, 0.003092766, 
    0.003038729, 0.002130336, 0.002817031, 0.00307535, 0.002910361, 
    0.002617441, 0.002637198, 0.002817394, 0.002794554, 0.002981331, 
    0.0027768, 0.002781283, 0.003068766, 0.003122712, 0.003172683, 
    0.003274456, 0.003344791, 0.003360877, 0.003393332, 0.003302766, 
    0.003239488,
  0.003124079, 0.003088681, 0.003137479, 0.002381852, 0.002821384, 
    0.002910489, 0.003166139, 0.002813898, 0.002786464, 0.002783888, 
    0.002758492, 0.003206221, 0.003227249, 0.003409561, 0.003516421, 
    0.003593571, 0.003583893, 0.003512397, 0.003481485, 0.00343976, 
    0.003538594, 0.003510524, 0.003534762, 0.003403712, 0.003432527, 
    0.003222037, 0.003325669, 0.00347794, 0.003187278, 0.00324529, 
    0.003047405, 0.003130376, 0.002882117, 0.003067, 0.003216377, 
    0.003223786, 0.003114544, 0.002810655, 0.002723409, 0.002990054, 
    0.003031889, 0.002954895, 0.002883561, 0.002779707, 0.002598176, 
    0.002441883, 0.002418963, 0.002443472, 0.002542257, 0.002533961, 
    0.002563223, 0.002651976, 0.002751382, 0.002848515, 0.003018443, 
    0.003106132, 0.003179852, 0.00323922, 0.003259612, 0.003262267, 
    0.003291877, 0.003283914, 0.003256671, 0.003315449, 0.003317134, 
    0.003339672, 0.003346713, 0.003334396, 0.003323603, 0.003261836, 
    0.003175259, 0.003113477, 0.003043557, 0.002966326, 0.00288992, 
    0.003137542, 0.00271079, 0.003445134, 0.003234625, 0.002631031, 
    0.002391787, 0.002174332, 0.002324488, 0.002814516, 0.002940767, 
    0.003052585, 0.003044605, 0.003144359, 0.003237853, 0.003213199, 
    0.003215868, 0.003224881, 0.003209146, 0.003180567, 0.003162464, 
    0.003124475,
  0.003191631, 0.003193315, 0.003195699, 0.00268857, 0.00254056, 0.002866589, 
    0.002591914, 0.002315652, 0.002813423, 0.003245135, 0.003281565, 
    0.003420023, 0.003422689, 0.003401231, 0.003563913, 0.003626155, 
    0.003548004, 0.003406461, 0.003435405, 0.003409624, 0.003408099, 
    0.003379123, 0.003391633, 0.00335053, 0.003402948, 0.003178691, 
    0.003397195, 0.003236663, 0.00298945, 0.003093466, 0.003316117, 
    0.002797291, 0.002458051, 0.002995744, 0.003022067, 0.003007555, 
    0.002933249, 0.002918083, 0.002959205, 0.003030809, 0.002912967, 
    0.002841171, 0.002873644, 0.00287536, 0.002826119, 0.00278597, 
    0.00275944, 0.002711773, 0.002732914, 0.002713203, 0.002707435, 
    0.002675295, 0.002687564, 0.002713583, 0.002759043, 0.00286077, 
    0.002953755, 0.003049331, 0.003112067, 0.003186531, 0.00320125, 
    0.003201075, 0.003242847, 0.00328031, 0.00328503, 0.00336789, 
    0.003352629, 0.003391922, 0.003380679, 0.003281401, 0.003177373, 
    0.003087489, 0.002943419, 0.002832651, 0.002659721, 0.002902621, 
    0.002786099, 0.003213836, 0.003212899, 0.002105778, 0.002326634, 
    0.001770547, 0.00217217, 0.00287573, 0.002819749, 0.002860995, 
    0.002891401, 0.003045628, 0.003147634, 0.003234593, 0.003263632, 
    0.003255844, 0.003295073, 0.003257623, 0.003275173, 0.003200913,
  0.003051504, 0.003360573, 0.003036007, 0.002963608, 0.003115704, 
    0.003386391, 0.003294105, 0.002879191, 0.003124161, 0.003408132, 
    0.003171414, 0.003343809, 0.003538676, 0.003430782, 0.003617112, 
    0.003705421, 0.003646707, 0.003550928, 0.003520664, 0.003475316, 
    0.003435502, 0.003393428, 0.003268655, 0.003286839, 0.003204869, 
    0.003365468, 0.003527388, 0.002734631, 0.002894593, 0.003136411, 
    0.003189724, 0.002948081, 0.003046608, 0.003129084, 0.002988324, 
    0.003054539, 0.003102113, 0.003223991, 0.003241984, 0.003242841, 
    0.003260121, 0.00330116, 0.003306165, 0.003339227, 0.003396034, 
    0.003412565, 0.003366152, 0.003370842, 0.003376961, 0.003350336, 
    0.003307167, 0.003252523, 0.003200103, 0.003136715, 0.0030248, 
    0.002962368, 0.002860673, 0.002796475, 0.002789833, 0.00284891, 
    0.002839534, 0.002860213, 0.002929719, 0.003002118, 0.003124699, 
    0.003233019, 0.003319582, 0.003418159, 0.003316863, 0.003313906, 
    0.003124889, 0.003096946, 0.003132105, 0.002978103, 0.002833797, 
    0.002722615, 0.002674122, 0.00307487, 0.003052127, 0.001490925, 
    0.002048764, 0.002507865, 0.002734583, 0.002650533, 0.002680272, 
    0.002664901, 0.002717847, 0.002792185, 0.002856113, 0.003020003, 
    0.003030924, 0.003105832, 0.003181346, 0.003121281, 0.002794681, 
    0.002816696,
  0.003357062, 0.003062826, 0.002674423, 0.002262516, 0.002467539, 
    0.002942739, 0.002740007, 0.002349524, 0.002605058, 0.002901062, 
    0.002456764, 0.002873518, 0.003132888, 0.002923602, 0.003471203, 
    0.00358841, 0.00346089, 0.003712878, 0.003699971, 0.003819242, 
    0.00365483, 0.003355948, 0.003265843, 0.003295677, 0.003079144, 
    0.003186416, 0.003377231, 0.003419479, 0.002882544, 0.002808459, 
    0.002993902, 0.002931755, 0.002961811, 0.002819158, 0.002962081, 
    0.003167534, 0.003206158, 0.003294166, 0.003294008, 0.003368346, 
    0.003368711, 0.003377199, 0.003370952, 0.003386592, 0.003404856, 
    0.003441684, 0.003412057, 0.003447039, 0.003447406, 0.003467228, 
    0.003445707, 0.003459839, 0.003431134, 0.003397785, 0.003277021, 
    0.003148766, 0.002961401, 0.002759159, 0.002591677, 0.002499506, 
    0.00245136, 0.002437294, 0.002483197, 0.002593361, 0.002714524, 
    0.002920851, 0.00320673, 0.003344154, 0.003378168, 0.003406746, 
    0.003261089, 0.003310522, 0.003150193, 0.003101923, 0.002781712, 
    0.002658578, 0.002806971, 0.002546553, 0.002373494, 0.00257591, 
    0.002804631, 0.002662966, 0.002667682, 0.002556929, 0.002486138, 
    0.002508119, 0.002589436, 0.00264346, 0.002732027, 0.002838915, 
    0.002850328, 0.003108868, 0.00312602, 0.003170731, 0.003554966, 
    0.003499368,
  0.003573374, 0.002925573, 0.002196887, 0.001650828, 0.001136336, 
    0.001541171, 0.001508222, 0.001653578, 0.001938123, 0.002200462, 
    0.001963666, 0.001433724, 0.001168504, 0.001256198, 0.002969552, 
    0.003220798, 0.003242906, 0.003476495, 0.003497412, 0.003736863, 
    0.003445724, 0.003867596, 0.003634008, 0.003386782, 0.003296375, 
    0.003241284, 0.003175052, 0.003225107, 0.002928767, 0.002385413, 
    0.002822367, 0.002877442, 0.002776591, 0.002988914, 0.002939383, 
    0.003069751, 0.003104066, 0.003207255, 0.003193393, 0.003209177, 
    0.003125383, 0.003125429, 0.003093772, 0.003120188, 0.003106438, 
    0.003138656, 0.003103737, 0.003136367, 0.003125319, 0.003149306, 
    0.003166439, 0.003180888, 0.003173813, 0.003163578, 0.003053509, 
    0.002922093, 0.002765642, 0.002589341, 0.002471816, 0.002382822, 
    0.002338301, 0.002335377, 0.00234749, 0.002361586, 0.002365418, 
    0.002427803, 0.002535393, 0.002936013, 0.003384478, 0.003359539, 
    0.003434896, 0.003274487, 0.002906658, 0.002429058, 0.002903845, 
    0.002931407, 0.002803916, 0.002719073, 0.002669051, 0.002638392, 
    0.002623117, 0.002520502, 0.002507007, 0.002383679, 0.002349729, 
    0.002365289, 0.002422128, 0.002497151, 0.002553831, 0.00258233, 
    0.002698948, 0.002710932, 0.00346567, 0.003713691, 0.004090486, 
    0.004017787,
  0.001270643, 0.001121919, 0.001107819, 0.0007234416, 3.004121e-005, 
    0.0005298941, 0.0007291953, 0.0007817908, 0.0009884671, 0.001590683, 
    0.002367323, 0.002202545, 0.0005118852, 0.0004672688, 0.001277796, 
    0.002624721, 0.00307104, 0.003034754, 0.003284028, 0.003501657, 
    0.003034164, 0.003933179, 0.003923718, 0.003607322, 0.003280386, 
    0.003177376, 0.003285584, 0.003545621, 0.002812419, 0.002162889, 
    0.002477013, 0.002595566, 0.002585048, 0.002601897, 0.002781631, 
    0.002799274, 0.002841221, 0.002881227, 0.002913004, 0.002914958, 
    0.002779266, 0.002754785, 0.002700172, 0.002708483, 0.002675742, 
    0.002725635, 0.002705785, 0.002728626, 0.002720868, 0.002746633, 
    0.002794381, 0.002791342, 0.002768202, 0.002749191, 0.002685804, 
    0.002559601, 0.002392962, 0.002231711, 0.002086259, 0.001967242, 
    0.001922022, 0.001912532, 0.00190948, 0.001924198, 0.001905094, 
    0.001813986, 0.001881966, 0.002288677, 0.002647944, 0.002988645, 
    0.002824882, 0.002606601, 0.001891218, 0.002700284, 0.002846736, 
    0.002728989, 0.002621781, 0.002478635, 0.002429761, 0.002303443, 
    0.002294098, 0.002253263, 0.00222405, 0.002168228, 0.002181612, 
    0.002119717, 0.002148709, 0.002145387, 0.00215378, 0.00217794, 
    0.00230276, 0.002340239, 0.002396044, 0.002010535, 0.001667405, 
    0.001450206,
  0.0007085651, 0.0007315008, 0.0003748108, 0.000445589, -0.0002854026, 
    0.0003050179, 0.000274658, 0.0001958848, 0.0003879545, 0.001101414, 
    0.002218185, 0.00108765, 0.0005616988, 0.0002275468, -0.0003381087, 
    0.0008629644, 0.002904166, 0.002967011, 0.002989472, 0.003000803, 
    0.002704034, 0.003035181, 0.004088566, 0.004112165, 0.003444418, 
    0.003380733, 0.00310507, 0.003577488, 0.002714716, 0.001960075, 
    0.002044173, 0.002371298, 0.002386462, 0.002331467, 0.002343722, 
    0.002421575, 0.002461104, 0.002515383, 0.002550017, 0.002548905, 
    0.002452696, 0.002407061, 0.002399623, 0.002395539, 0.002320534, 
    0.00233015, 0.002305287, 0.002300488, 0.002303379, 0.002291157, 
    0.002311454, 0.002347154, 0.002386254, 0.002344769, 0.002296418, 
    0.002195281, 0.002021077, 0.001868712, 0.001725278, 0.001601602, 
    0.001500991, 0.001444454, 0.00143328, 0.001482109, 0.001451639, 
    0.00138755, 0.001544732, 0.001805054, 0.001799284, 0.001774966, 
    0.001953986, 0.001957689, 0.001837605, 0.002659896, 0.002531849, 
    0.002463534, 0.00240401, 0.002262959, 0.002192721, 0.002154003, 
    0.002087388, 0.00196945, 0.002012556, 0.001964206, 0.001897846, 
    0.00188656, 0.001899038, 0.001822696, 0.001819914, 0.001814781, 
    0.001905603, 0.001914679, 0.001736864, 0.001033879, 0.0004455097, 
    0.0005335333,
  0.001194906, 0.0008851378, 0.0001978399, 7.192325e-005, 0.0002010188, 
    0.0002080281, -0.0002038949, 4.255027e-005, 0.0002178194, 0.0008725165, 
    0.001704981, 0.0004858975, 0.0005587265, 0.00036583, 4.959293e-006, 
    0.0005699326, 0.002659736, 0.002661612, 0.002182581, 0.002293939, 
    0.002351318, 0.002226656, 0.002625579, 0.003176786, 0.003433595, 
    0.003703675, 0.003058529, 0.002811735, 0.002316143, 0.001347894, 
    0.001517013, 0.002005977, 0.001875625, 0.001962841, 0.001920193, 
    0.00204449, 0.002150347, 0.002175412, 0.00215041, 0.00219369, 
    0.002206837, 0.002199635, 0.002114218, 0.002051943, 0.00195551, 
    0.001886481, 0.001834759, 0.00181637, 0.001888818, 0.001970213, 
    0.002015799, 0.002048447, 0.002073878, 0.002014512, 0.001954844, 
    0.001879758, 0.001757544, 0.001632582, 0.001519651, 0.001382274, 
    0.001268977, 0.001232468, 0.001214379, 0.001250682, 0.001251811, 
    0.001203412, 0.001323893, 0.001898021, 0.001442336, 0.001719318, 
    0.001845965, 0.002215451, 0.002380325, 0.002333929, 0.002239341, 
    0.00219342, 0.002060225, 0.002025892, 0.002024986, 0.002042916, 
    0.002095987, 0.002057364, 0.00202327, 0.00194429, 0.001964683, 
    0.001914757, 0.001882555, 0.00183047, 0.001772359, 0.001702978, 
    0.001679947, 0.001699847, 0.001394813, 0.001254575, 0.001257611, 
    0.00106314,
  0.0007834753, 0.001124319, 0.0009065471, 0.0004564128, 0.0009608911, 
    0.0009731296, 0.0003709313, 7.605576e-005, 0.0003247256, 0.0004545054, 
    0.0006552222, 0.0002479551, 0.0006190622, 0.0007030647, 0.001371908, 
    0.00126737, 0.001074202, 0.001142152, 0.001416095, 0.001711765, 
    0.00216826, 0.002190907, 0.001665512, 0.001455292, 0.002007977, 
    0.002560663, 0.002405293, 0.002139837, 0.001855104, 0.001281931, 
    0.001308316, 0.001293582, 0.001541155, 0.001714072, 0.001734816, 
    0.001843216, 0.001872574, 0.001882412, 0.001956131, 0.00202537, 
    0.00204441, 0.002018596, 0.001954654, 0.001820996, 0.00166906, 
    0.001558989, 0.001514612, 0.001493121, 0.001533082, 0.001640308, 
    0.001690581, 0.001708159, 0.001713453, 0.001671586, 0.001650081, 
    0.001610138, 0.001504916, 0.001422169, 0.00132235, 0.001183703, 
    0.00106991, 0.001041904, 0.001046417, 0.001075108, 0.001030587, 
    0.001094325, 0.0009216471, 0.001129341, 0.00119063, 0.001558512, 
    0.002153192, 0.002179943, 0.002272321, 0.002097768, 0.002028658, 
    0.001937948, 0.001887102, 0.001868632, 0.001847652, 0.001863705, 
    0.001851958, 0.00183902, 0.001852181, 0.001879822, 0.001945069, 
    0.001915568, 0.001916092, 0.001832598, 0.001738884, 0.001689723, 
    0.001547752, 0.001513292, 0.001670425, 0.001344474, 0.001111047, 
    0.0006447318,
  0.0008952143, 0.0007647509, 0.0002077899, 0.0008889521, 0.001311509, 
    0.001465383, 0.001252524, 0.0008011982, 0.001663843, 0.001139562, 
    0.000875426, 0.0006991234, 0.001042398, 0.001261298, 0.0006149458, 
    0.000473341, 0.0004432206, 0.0004158821, 0.0004645512, 0.001440031, 
    0.001790999, 0.0009505746, 0.001035389, 0.000878572, 0.0008383589, 
    0.001331981, 0.001361466, 0.001789634, 0.001742665, 0.001684492, 
    0.001794227, 0.001615603, 0.001552851, 0.00112063, 0.001429382, 
    0.001723304, 0.001666388, 0.001714278, 0.001822268, 0.001827354, 
    0.001803082, 0.001762503, 0.001725009, 0.001660126, 0.001538231, 
    0.001431848, 0.001372037, 0.001335877, 0.001332377, 0.001364055, 
    0.001417874, 0.001498253, 0.001544697, 0.001506963, 0.001463491, 
    0.001387341, 0.001260772, 0.001134856, 0.001078875, 0.001034799, 
    0.0009687254, 0.0008695908, 0.0008325409, 0.0008573839, 0.0008555884, 
    0.000965707, 0.0008422057, 0.001010704, 0.001147747, 0.001643101, 
    0.001455449, 0.001726201, 0.00183333, 0.001749262, 0.001769496, 
    0.001829834, 0.001858681, 0.001735723, 0.00171757, 0.001701612, 
    0.001616401, 0.001549055, 0.001505727, 0.001529425, 0.001618435, 
    0.001712054, 0.001728425, 0.00160661, 0.001591335, 0.001604416, 
    0.001489416, 0.001419496, 0.00141433, 0.001520298, 0.001518138, 
    0.0008900329,
  0.001351197, 0.001288764, 0.001044734, 0.001379155, 0.001452859, 
    0.001468244, 0.001365883, 0.00138049, 0.001596577, 0.001504499, 
    0.001314767, 0.0009012865, 0.0007148273, 0.0007279562, 0.0005518598, 
    0.0003204187, 0.0006361012, 0.0009100121, 0.001308998, 0.001496108, 
    0.001264763, 0.001260265, 0.001233769, 0.0009071187, 0.001020034, 
    0.0008569246, 0.0008532838, 0.0008129287, 0.001183049, 0.001408132, 
    0.001722241, 0.001549117, 0.001374786, 0.000933568, 0.001424885, 
    0.001534222, 0.001383814, 0.001459901, 0.001543649, 0.001591205, 
    0.001575993, 0.001494661, 0.001454256, 0.001424645, 0.001398562, 
    0.001395272, 0.001395209, 0.001356298, 0.001301288, 0.001285472, 
    0.001303132, 0.001326306, 0.001348351, 0.001333237, 0.001287205, 
    0.001213836, 0.001117833, 0.00101269, 0.0008888887, 0.000835482, 
    0.0008247849, 0.0007761475, 0.0007474413, 0.0007309755, 0.0004764241, 
    0.0003809775, 0.0005234722, 0.0005942825, 0.0008058716, 0.0006973115, 
    0.001203123, 0.001520967, 0.001612742, 0.001681026, 0.001690594, 
    0.001762198, 0.001703994, 0.001667502, 0.001623601, 0.001587965, 
    0.001572865, 0.001505839, 0.001342553, 0.001291007, 0.001252049, 
    0.001238934, 0.001265668, 0.001252603, 0.001241524, 0.001267639, 
    0.001326847, 0.001306628, 0.001240714, 0.00135792, 0.001357984, 
    0.001457945,
  0.001368428, 0.001191266, 0.001205604, 0.001254638, 0.001260169, 
    0.001342837, 0.001302767, 0.001186594, 0.001220178, 0.001307821, 
    0.001251984, 0.001405637, 0.001462969, 0.001259471, 0.0009136675, 
    0.0003773845, -0.00042208, -0.0001492337, 0.001435931, 0.001213201, 
    0.000776625, 0.0008885388, 0.001023086, 0.0006775693, 0.0006376421, 
    0.0007286868, 0.0006465917, 0.0007197065, 0.0007800106, 0.0008910028, 
    0.0007937592, 0.0008666199, 0.0009502256, 0.0008327961, 0.0008723256, 
    0.001156267, 0.001156314, 0.001092403, 0.001204379, 0.001305945, 
    0.001311144, 0.001260344, 0.00127864, 0.001249536, 0.001213805, 
    0.001216269, 0.00121611, 0.001204666, 0.001171843, 0.001151863, 
    0.001148272, 0.001137558, 0.001142201, 0.001170381, 0.001148717, 
    0.001074854, 0.001008988, 0.0009097736, 0.0008055684, 0.000749032, 
    0.0007151444, 0.0007267636, 0.000683785, 0.0004487359, 0.0003862069, 
    0.0006116717, 0.0006338283, 0.0004776311, 0.000580057, 0.0007609529, 
    0.001017157, 0.001632484, 0.001743983, 0.001805146, 0.00167648, 0.00172, 
    0.001814477, 0.001715214, 0.001589234, 0.00154395, 0.001598771, 
    0.001541852, 0.001333983, 0.001003217, 0.0005201008, 0.0003064303, 
    0.000535694, 0.0007487927, 0.0007842211, 0.0008158358, 0.001000388, 
    0.001092005, 0.001050122, 0.001106993, 0.001147111, 0.00117197,
  0.001088985, 0.001121457, 0.001073011, 0.000977437, 0.001193809, 
    0.001259629, 0.001329613, 0.001244879, 0.001249663, 0.001314783, 
    0.001258596, 0.001672793, 0.001623043, 0.001017969, 0.0005246168, 
    0.0004440155, 0.0003614114, -0.0001437338, 0.0004055984, 0.0009014453, 
    0.0007000444, 0.0006868527, 0.0007317704, 0.0008016429, 0.0007824583, 
    0.0006732943, 0.0006084125, 0.0006101767, 0.0008112746, 0.0007944899, 
    0.000691684, 0.0006684775, 0.0007172583, 0.0006906504, 0.0006552697, 
    0.0007130143, 0.0008940543, 0.0009272425, 0.0009837304, 0.001183367, 
    0.001105261, 0.0009867991, 0.0008982825, 0.0008151373, 0.0007692343, 
    0.0007736688, 0.0007813303, 0.000840331, 0.0009100125, 0.0009415313, 
    0.000942294, 0.0009078663, 0.0008899537, 0.000916895, 0.0009029713, 
    0.0008735978, 0.0008216389, 0.000741371, 0.0006844681, 0.0006479896, 
    0.0006127357, 0.0006145481, 0.0006034849, 0.0003931369, 0.0005726661, 
    0.0008925283, 0.0008373894, 0.0005539414, 0.0006842613, 0.001261187, 
    0.001088302, 0.001681424, 0.002024492, 0.001940903, 0.001375437, 
    0.001941157, 0.001939711, 0.001778794, 0.001638206, 0.001599853, 
    0.001302529, 0.001085139, 0.0008790977, 0.0006008311, 0.0003773696, 
    0.0002725916, 0.000258971, 0.0003129486, 0.0003780685, 0.0004872484, 
    0.000655476, 0.0008372627, 0.0009583635, 0.001010546, 0.001018588, 
    0.001015917,
  0.000928482, 0.001021211, 0.001017873, 0.00109706, 0.001250649, 0.00139219, 
    0.001403475, 0.001484347, 0.001339214, 0.001189614, 0.001137702, 
    0.001435455, 0.001440844, 0.001166932, 0.0009471579, 0.0008808468, 
    0.0007862574, 0.000613308, 0.0006595938, 0.0008404106, 0.0009117927, 
    0.0007620649, 0.0005716165, 0.0006051385, 0.0006663164, 0.0005485213, 
    0.0006443814, 0.000659402, 0.0007159547, 0.0007056552, 0.0007176874, 
    0.000669813, 0.0006254034, 0.0006442389, 0.0006140394, 0.0005555314, 
    0.0005162081, 0.0007062596, 0.0007297988, 0.0006969774, 0.0006971681, 
    0.0006389937, 0.0006368316, 0.0006333827, 0.0006461458, 0.0006568593, 
    0.0006661573, 0.0006968337, 0.000744279, 0.0007600943, 0.0007483168, 
    0.0007316116, 0.0007065139, 0.0007009516, 0.0006714505, 0.0006231153, 
    0.0005833949, 0.0005654502, 0.0005753678, 0.0005956497, 0.0005911356, 
    0.0006160904, 0.0006835307, 0.0005353931, 0.0007699812, 0.0009240475, 
    0.0007232351, 0.0005542273, 0.0006603552, 0.0009384002, 0.00111483, 
    0.001349338, 0.001403427, 0.001124716, 0.00137488, 0.001528884, 
    0.001581796, 0.001481279, 0.001361609, 0.001230177, 0.0009879747, 
    0.0007610801, 0.0006572406, 0.0005270955, 0.0004285183, 0.0004351619, 
    0.0003671013, 0.0002110009, 0.0001180009, 0.0002085692, 0.0004305206, 
    0.0006574155, 0.0008311905, 0.0009148284, 0.0009337272, 0.0009141448,
  0.0008145333, 0.0009480002, 0.001032639, 0.001143058, 0.001184305, 
    0.001223628, 0.001254574, 0.001315895, 0.001312876, 0.001241557, 
    0.001156807, 0.001162942, 0.001133665, 0.00101881, 0.000833781, 
    0.0006723716, 0.0005728565, 0.0005776407, 0.0005461378, 0.0004747228, 
    0.0004489101, 0.000504192, 0.0005372998, 0.0005352974, 0.0004511995, 
    0.0004763766, 0.0005625251, 0.0006369117, 0.0005906743, 0.0005357109, 
    0.0006436349, 0.0006053611, 0.0005884808, 0.0005636378, 0.0004838309, 
    0.0003955367, 0.0002943361, 0.0003883846, 0.0005398754, 0.0006450657, 
    0.00076464, 0.0007076899, 0.0006871542, 0.0006743756, 0.0006808916, 
    0.0006607689, 0.0006612933, 0.0006668884, 0.0006619773, 0.0006653629, 
    0.0006863112, 0.000700505, 0.0006942106, 0.0006697495, 0.0006398684, 
    0.0005914695, 0.0005441676, 0.0005447553, 0.0005562468, 0.0005507474, 
    0.000549031, 0.0006462899, 0.000632382, 0.0007462979, 0.0005434195, 
    0.0005490144, 0.0005890527, 0.0005771634, 0.0006783807, 0.0008007046, 
    0.0009593484, 0.001094564, 0.001097107, 0.001122793, 0.001201741, 
    0.001220099, 0.001079448, 0.0009065315, 0.0008515203, 0.0008013886, 
    0.0007795019, 0.0007545156, 0.0005686446, 0.0006252928, 0.0005598865, 
    0.0004635011, 0.0002813349, -3.925525e-006, -0.0001665745, 
    -9.614555e-005, 0.0001807059, 0.0004795236, 0.0006650132, 0.0007400992, 
    0.0007547061, 0.0007471885,
  0.0006687492, 0.0007018414, 0.0008766018, 0.001010147, 0.001070213, 
    0.00110898, 0.001064443, 0.001056273, 0.00105478, 0.0009617642, 
    0.0009638306, 0.0009411494, 0.0008510591, 0.0007357914, 0.0006347022, 
    0.0005337875, 0.0004191878, 0.0003616812, 0.0003596945, 0.0003770355, 
    0.000354243, 0.0004113996, 0.0004163587, 0.0003492839, 0.0003159689, 
    0.0002663459, 0.0002659329, 0.0003197361, 0.0003162872, 0.0003721882, 
    0.0003848244, 0.0003503968, 0.0003352492, 0.0003050495, 0.0002975791, 
    0.0002593365, 0.0002578584, 0.0003293204, 0.0005133159, 0.0006312693, 
    0.000743469, 0.0007028105, 0.0005355519, 0.0005811851, 0.0006376584, 
    0.0006167251, 0.000624832, 0.0006400582, 0.0006441909, 0.0006693837, 
    0.0007288458, 0.0008046944, 0.0008246419, 0.0007600305, 0.0007055923, 
    0.0006701155, 0.000607904, 0.0006172666, 0.0006236718, 0.0006285356, 
    0.0006206995, 0.0006237188, 0.0006708147, 0.000437228, 0.0003465656, 
    0.0003694694, 0.0005052248, 0.0005942185, 0.0007356959, 0.000863584, 
    0.0009434861, 0.001021354, 0.001087093, 0.001135238, 0.001089049, 
    0.0009040682, 0.0007980831, 0.0006757108, 0.0005919624, 0.0005166538, 
    0.0004433163, 0.0004091745, 0.0004688583, 0.0004545848, 0.0003795945, 
    0.0003711698, 0.0002289615, -2.382603e-005, -0.0002243356, -0.0001978711, 
    2.722768e-005, 0.000310644, 0.0005471869, 0.0006273594, 0.0006049797, 
    0.0006537922,
  0.0005215812, 0.0006122594, 0.0006618812, 0.000868177, 0.0008829911, 
    0.0008854235, 0.0007607935, 0.000991964, 0.000966629, 0.0008910501, 
    0.0008661749, 0.0008660795, 0.0008544924, 0.0007610642, 0.0007056398, 
    0.0006776338, 0.0006110512, 0.0004928592, 0.0003971737, 0.0003696762, 
    0.0004115426, 0.0003851098, 0.000444921, 0.0004641376, 0.0004470197, 
    0.0003446903, 0.0002928264, 0.0002986599, 0.0003335485, 0.0003244408, 
    0.0002909671, 0.0002635967, 0.0002354155, 0.0002017826, 0.0001904498, 
    0.000191753, 0.0002344936, 0.0003367433, 0.0005145239, 0.00055434, 
    0.0004738651, 0.000381788, 0.0003231856, 0.000351621, 0.0004887264, 
    0.0005837444, 0.0007218681, 0.000862662, 0.0009827774, 0.001072137, 
    0.001132695, 0.001059628, 0.0009091855, 0.0008638704, 0.0007013318, 
    0.0006741839, 0.0006191093, 0.000602548, 0.0006059809, 0.0006018798, 
    0.0006680968, 0.0004328571, 0.000313648, 0.0002952896, 0.0003923895, 
    0.000472371, 0.0005579793, 0.0006308239, 0.0006847065, 0.0007496201, 
    0.0007433741, 0.0008099406, 0.0007010471, 0.0007261605, 0.0007434855, 
    0.0007354588, 0.0006770464, 0.0006117832, 0.0005433729, 0.0004759323, 
    0.0004205077, 0.0003662752, 0.0002361939, 1.843786e-005, 2.299971e-005, 
    0.0002583507, 0.0004000021, 0.0003263312, 0.000216166, 0.0001612832, 
    0.0002167234, 0.0003482662, 0.0004605618, 0.0004876619, 0.0004869783, 
    0.0005184505,
  0.0004017996, 0.0004367027, 0.0006186329, 0.0005508587, 0.0005621277, 
    0.0004715126, 0.0006898406, 0.0007468385, 0.0007613027, 0.0007484439, 
    0.0007603015, 0.0007749721, 0.0007528949, 0.0006978837, 0.0006299184, 
    0.0006042805, 0.0005667377, 0.0004580346, 0.0003791022, 0.0003072113, 
    0.0002706059, 0.0002788393, 0.0003001221, 0.0003235029, 0.000317622, 
    0.0003105965, 0.0003163348, 0.0003418296, 0.000350222, 0.0003130605, 
    0.0002591619, 0.0002346206, 0.000220999, 0.0001827409, 0.000164144, 
    0.0001868734, 0.0002340168, 0.0002207288, 0.000210588, 0.0001711694, 
    0.0001757154, 0.0001963783, 0.0002059788, 0.0002281676, 0.0002917777, 
    0.0004191248, 0.0005772285, 0.0009313112, 0.001002455, 0.0009717152, 
    0.0009119036, 0.0007881008, 0.0008847876, 0.0007995607, 0.0006922884, 
    0.0005455657, 0.000428661, 0.0003729505, 0.0003552439, 0.0003519538, 
    0.000361999, 0.000345167, 0.0003484094, 0.0004025623, 0.000513236, 
    0.0006262304, 0.0006617073, 0.0006436037, 0.0006372619, 0.0006473553, 
    0.0006504866, 0.0006082704, 0.0005886883, 0.0005846829, 0.0005970648, 
    0.0006085566, 0.0005302281, 0.0004434597, 0.0003884484, 0.0003524155, 
    0.0003257601, 0.0002907127, 0.0001817711, 9.805406e-005, 0.0001744751, 
    0.0001360897, 0.0002192657, 0.0003205938, 0.0003687218, 0.0003604568, 
    0.0003619357, 0.0003044452, 0.0001625703, 0.0001864284, 0.0003282558, 
    0.0003790064,
  0.0002337615, 0.0002711294, 0.0002917447, 0.0005452158, 0.0005108519, 
    0.0004703046, 0.0004076008, 0.0005378253, 0.0005856204, 0.0006063788, 
    0.0006469418, 0.0006711013, 0.0006769504, 0.0006546823, 0.0006106388, 
    0.0005471556, 0.0004744381, 0.0004171223, 0.0003805329, 0.0003527651, 
    0.0003432761, 0.000339954, 0.0003233441, 0.0003057806, 0.0002901403, 
    0.000284339, 0.0002948612, 0.000293685, 0.00026366, 0.0002168664, 
    0.0001904338, 0.0001889715, 0.0001763669, 0.0001655269, 0.0001632541, 
    0.0001928021, 0.0002235102, 0.0002062487, 0.0001673549, 0.0001417169, 
    0.0001393011, 0.0001778133, 0.0001911966, 0.0001964101, 0.0002129565, 
    0.0002486239, 0.0002954017, 0.0003444683, 0.0003930739, 0.0004386274, 
    0.0005266358, 0.0005986857, 0.0006673505, 0.0006278362, 0.0005343121, 
    0.0004511042, 0.0003609983, 0.0003070679, 0.0002907122, 0.0002995655, 
    0.0003241862, 0.0003930258, 0.0004446674, 0.0004743901, 0.0004934319, 
    0.0005250307, 0.0005211044, 0.0005552302, 0.0005625576, 0.000542133, 
    0.0005004258, 0.0004561433, 0.000427676, 0.0004143883, 0.0004365136, 
    0.000417154, 0.0003859688, 0.0002908556, 0.0002350657, 0.0002328405, 
    0.0002688895, 0.0002806354, 0.000230949, 0.0001933742, 0.0001546233, 
    0.0001200525, 9.865849e-005, 0.0001288892, 0.0001562119, 0.0003524781, 
    0.0004904908, 0.0005027298, 0.000373268, 0.0001516659, 8.344604e-005, 
    0.0001400942,
  0.0002122084, 0.0001642541, 0.0001589614, 0.0001174291, -1.122127e-005, 
    0.0002611643, 0.0003197677, 0.0004083485, 0.0005204848, 0.0005966674, 
    0.000619762, 0.000634274, 0.0005801369, 0.0005256186, 0.0004640431, 
    0.0004381188, 0.0004128782, 0.0003949493, 0.0003776559, 0.0003648289, 
    0.0003433077, 0.0003161121, 0.0003039209, 0.0002899814, 0.0002752473, 
    0.000269843, 0.0002312191, 0.0002082355, 0.000183297, 0.0001685944, 
    0.0001672435, 0.0001577386, 0.0001454521, 0.0001264738, 0.0001268713, 
    0.000137457, 0.0001493623, 0.000153479, 0.0001327999, 0.0001216579, 
    0.0001231996, 0.0001568008, 0.0001954723, 0.0002088397, 0.0002288191, 
    0.0002364008, 0.0002511827, 0.0002767411, 0.0003107873, 0.0003682304, 
    0.0004470199, 0.0005260636, 0.000586781, 0.0005454232, 0.0005253325, 
    0.0005141904, 0.0005088656, 0.0005187043, 0.0005108365, 0.0005166857, 
    0.0005194355, 0.0005395423, 0.0005483, 0.0005542604, 0.0005530525, 
    0.0005461702, 0.0005361407, 0.0005109637, 0.000496722, 0.0005026826, 
    0.0004622944, 0.0004397559, 0.0004039772, 0.0003947743, 0.000353957, 
    0.0003458826, 0.0002937484, 0.0002722112, 0.0002501814, 0.0002360353, 
    0.0001984447, 0.0001841395, 0.0001275389, 0.0001084336, 9.239593e-005, 
    7.300457e-005, 5.691923e-005, 6.599509e-005, 0.0001065105, 0.0001832971, 
    0.0002847522, 0.0003953942, 0.0005367446, 0.0006045981, 0.0004332229, 
    0.0003025692,
  0.0004564764, 0.0003394922, 0.0002507369, 0.000210301, 0.0002006216, 
    0.0002594313, 0.0004211904, 0.0006133877, 0.0008360709, 0.0009107279, 
    0.0008658736, 0.0007655155, 0.0006073802, 0.0004805573, 0.0004232575, 
    0.0003513343, 0.0003450402, 0.00033962, 0.0003459621, 0.0003329762, 
    0.0003316252, 0.0003208964, 0.0003094999, 0.0002949881, 0.0002721635, 
    0.0002489574, 0.0002206811, 0.000186762, 0.0001734106, 0.0001505066, 
    0.0001463421, 0.0001280952, 0.0001180339, 9.710074e-005, 7.654907e-005, 
    8.030009e-005, 8.390821e-005, 7.917167e-005, 8.920114e-005, 0.000103999, 
    0.000111088, 0.0001282064, 0.0001561649, 0.000181024, 0.0002000021, 
    0.0002074249, 0.0002095865, 0.0002183922, 0.0002389915, 0.0002667753, 
    0.0003029354, 0.0003384438, 0.0003668793, 0.0003912457, 0.0004195221, 
    0.0004457163, 0.0004683025, 0.0004839428, 0.0004918742, 0.000493432, 
    0.0004888702, 0.0004862794, 0.0004882503, 0.0004273422, 0.0003981757, 
    0.0003732054, 0.0003557691, 0.0003382691, 0.000344166, 0.0003728716, 
    0.0003512867, 0.0003397632, 0.0003212301, 0.0002649951, 0.0002338895, 
    0.0002111284, 0.0002030222, 0.0002161352, 0.0002122728, 0.0002020844, 
    0.0001842191, 0.0001555928, 0.0001247573, 0.0001121689, 0.0001014559, 
    7.929886e-005, 5.394695e-005, 3.916497e-005, 5.388341e-005, 0.000107019, 
    0.0001918642, 0.0003147135, 0.0004381032, 0.0005556276, 0.000629394, 
    0.0005852066,
  0.0005597757, 0.0005356953, 0.0005189423, 0.0005655927, 0.0007022389, 
    0.0007924885, 0.0007800431, 0.0006299824, 0.00055674, 0.0004913814, 
    0.0004483867, 0.0004009256, 0.0003571677, 0.000308133, 0.000270892, 
    0.0002453971, 0.0002293436, 0.0002231447, 0.0002274999, 0.0002365597, 
    0.0002441732, 0.0002491959, 0.0002449202, 0.0002372431, 0.0002246228, 
    0.0002092847, 0.0001885423, 0.0001573094, 0.0001426706, 0.0001291601, 
    0.0001105635, 9.505043e-005, 8.389237e-005, 7.567497e-005, 7.348147e-005, 
    7.786835e-005, 8.624478e-005, 9.559083e-005, 0.0001088628, 0.0001214354, 
    0.0001393327, 0.0001562604, 0.0001719801, 0.0001839965, 0.0001914033, 
    0.0001968552, 0.0002030064, 0.0002132425, 0.000229439, 0.0002525974, 
    0.0002809374, 0.0003093568, 0.0003356465, 0.0003574856, 0.0003717748, 
    0.000380644, 0.000383362, 0.0003845858, 0.0003867793, 0.0003936935, 
    0.0003998606, 0.0004086662, 0.0004143087, 0.0004132914, 0.0004174717, 
    0.000328637, 0.0003090866, 0.0002948769, 0.0002874065, 0.0002910145, 
    0.0002866594, 0.0002756763, 0.0002604651, 0.0002429812, 0.0002238918, 
    0.0002106039, 0.0001834401, 0.0001762239, 0.0001430997, 0.0001300821, 
    0.0001146484, 9.732321e-005, 8.258902e-005, 7.122432e-005, 6.233924e-005, 
    5.599734e-005, 5.432841e-005, 6.31022e-005, 8.400355e-005, 0.0001234222, 
    0.000176065, 0.0002442209, 0.000320165, 0.00037551, 0.0004330168, 
    0.0005211841,
  0.0003484575, 0.0003656872, 0.0003897834, 0.0004230826, 0.0003442931, 
    0.0003370293, 0.0003254104, 0.0003444362, 0.0003242501, 0.0003089277, 
    0.000295163, 0.0002831149, 0.0002739914, 0.0002658693, 0.0002592572, 
    0.0002532013, 0.0002465097, 0.0002399294, 0.0002333013, 0.0002252746, 
    0.0002184241, 0.0002124, 0.0002072025, 0.0002006062, 0.0002011148, 
    0.0001622845, 0.0001522232, 0.0001551636, 0.0001401274, 0.0001269031, 
    0.0001165239, 0.0001064468, 9.819746e-005, 9.449403e-005, 9.350857e-005, 
    9.670333e-005, 0.0001034744, 0.0001109926, 0.000122548, 0.0001341033, 
    0.0001451183, 0.0001564988, 0.0001671005, 0.0001756359, 0.0001836627, 
    0.0001906563, 0.0001991122, 0.0002092053, 0.0002195367, 0.0002305517, 
    0.0002428223, 0.0002526928, 0.0002597182, 0.0002629925, 0.0002629925, 
    0.0002609421, 0.0002571592, 0.0002540439, 0.0002535352, 0.000256444, 
    0.0002615143, 0.0002673159, 0.0002736419, 0.0002801586, 0.0002841799, 
    0.0002797293, 0.0002765346, 0.0002702562, 0.000260799, 0.0002526928, 
    0.0002533126, 0.0002024659, 0.0001849341, 0.0001592485, 0.0001452136, 
    0.000130972, 0.0001173663, 0.0001043645, 9.431917e-005, 8.587915e-005, 
    7.842467e-005, 7.30523e-005, 7.13357e-005, 7.233702e-005, 7.685111e-005, 
    8.417849e-005, 9.52729e-005, 0.0001080839, 0.0001245507, 0.0001459924, 
    0.0001714714, 0.0001986352, 0.0002551882, 0.0002765981, 0.0003021089, 
    0.0003251401,
  0.0002245116, 0.0002178836, 0.0002120821, 0.000205915, 0.0001972842, 
    0.0001886217, 0.0001808969, 0.0001746663, 0.0001680541, 0.0001629997, 
    0.0001596618, 0.0001578021, 0.0001569438, 0.000156769, 0.0001569278, 
    0.0001564828, 0.0001557675, 0.0001538443, 0.0001513489, 0.0001485515, 
    0.0001456428, 0.0001417804, 0.0001380451, 0.0001342305, 0.0001308926, 
    0.000127221, 0.0001252501, 0.0001206565, 0.0001173981, 0.0001155702, 
    0.0001166193, 0.0001171278, 0.0001188763, 0.0001209743, 0.0001248685, 
    0.0001281269, 0.0001322913, 0.0001377273, 0.0001433222, 0.0001502681, 
    0.000156896, 0.0001636672, 0.0001696912, 0.0001756834, 0.0001808809, 
    0.0001858083, 0.0001900203, 0.0001937874, 0.0001968709, 0.0002008605, 
    0.0002047069, 0.0002094753, 0.0002139894, 0.0002185194, 0.0002229222, 
    0.0002270389, 0.0002309331, 0.000235304, 0.0002408513, 0.0002467322, 
    0.0002513575, 0.0002559034, 0.0002603061, 0.0002629606, 0.0002636123, 
    0.0002624201, 0.0002594797, 0.0002542662, 0.0002466845, 0.000239818, 
    0.0002334444, 0.0002246229, 0.000221285, 0.000218122, 0.0002118119, 
    0.0002088078, 0.0002058514, 0.0002003678, 0.000198699, 0.0002003996, 
    0.0001976975, 0.0001978883, 0.0002012738, 0.0002015599, 0.0002029428, 
    0.0002055176, 0.0002093164, 0.0002131788, 0.0002187419, 0.0002238123, 
    0.0002279131, 0.0002364961, 0.0002342391, 0.0002297887, 0.0002283741, 
    0.0002268322,
  0.0002116689, 0.0002072502, 0.0002061217, 0.0002043256, 0.0002027202, 
    0.0002009241, 0.0001987942, 0.0001965848, 0.0001946933, 0.0001927701, 
    0.000191435, 0.000189766, 0.0001878269, 0.0001865395, 0.0001849023, 
    0.0001830267, 0.0001816439, 0.0001804995, 0.0001791484, 0.0001770663, 
    0.0001758265, 0.0001740622, 0.0001727748, 0.000171837, 0.0001703906, 
    0.0001683879, 0.0001669574, 0.0001660514, 0.0001644778, 0.0001628725, 
    0.0001614738, 0.0001599479, 0.0001583901, 0.0001569596, 0.0001561172, 
    0.0001559583, 0.0001563079, 0.0001559265, 0.0001551477, 0.0001544166, 
    0.0001537808, 0.0001533993, 0.0001536854, 0.0001542576, 0.0001543053, 
    0.0001540351, 0.0001542099, 0.000154957, 0.0001557199, 0.0001566577, 
    0.0001576908, 0.0001592961, 0.0001607584, 0.0001621413, 0.0001628883, 
    0.0001643983, 0.000165956, 0.0001679905, 0.000169723, 0.0001716304, 
    0.0001730291, 0.0001742371, 0.0001757947, 0.0001772888, 0.0001784332, 
    0.0001794346, 0.0001806585, 0.0001813578, 0.0001818824, 0.0001822956, 
    0.0001828996, 0.0001828678, 0.0001827725, 0.0001834718, 0.0001842348, 
    0.0001851884, 0.0001862216, 0.000186762, 0.000187811, 0.0001888919, 
    0.0001900522, 0.0001917847, 0.0001939781, 0.00019641, 0.0001985716, 
    0.0002009081, 0.0002031016, 0.0002054222, 0.0002071229, 0.0002092052, 
    0.0002112874, 0.0002130357, 0.0002130198, 0.0002123681, 0.0002117483, 
    0.000211955,
  6.462073e-006, 5.937552e-006, 5.540191e-006, 5.190508e-006, 4.936195e-006, 
    4.76135e-006, 4.475254e-006, 4.3481e-006, 4.205047e-006, 4.061996e-006, 
    3.966628e-006, 3.871259e-006, 3.744106e-006, 3.616949e-006, 
    3.569266e-006, 3.521583e-006, 3.473901e-006, 3.489793e-006, 
    3.410321e-006, 3.585163e-006, 3.744108e-006, 3.966632e-006, 
    4.205051e-006, 4.618305e-006, 5.079248e-006, 5.603768e-006, 
    6.144184e-006, 6.827649e-006, 7.479328e-006, 8.258161e-006, 
    9.084681e-006, 9.799931e-006, 1.061056e-005, 1.145297e-005, 
    1.229538e-005, 1.320138e-005, 1.412326e-005, 1.501336e-005, 
    1.599882e-005, 1.695249e-005, 1.795384e-005, 1.893931e-005, 1.98453e-005, 
    2.087844e-005, 2.186391e-005, 2.288118e-005, 2.370768e-005, 
    2.447062e-005, 2.531303e-005, 2.601241e-005, 2.667998e-005, 
    2.725219e-005, 2.758596e-005, 2.80787e-005, 2.803102e-005, 2.820585e-005, 
    2.831712e-005, 2.814228e-005, 2.757007e-005, 2.710913e-005, 
    2.682303e-005, 2.629851e-005, 2.575808e-005, 2.515409e-005, 
    2.448651e-005, 2.386662e-005, 2.323084e-005, 2.27699e-005, 2.230896e-005, 
    2.18957e-005, 2.15937e-005, 2.137118e-005, 2.121223e-005, 2.087844e-005, 
    2.079897e-005, 2.086255e-005, 2.075129e-005, 2.086255e-005, 
    2.092613e-005, 2.081487e-005, 2.052876e-005, 2.021087e-005, 
    1.960688e-005, 1.898699e-005, 1.811279e-005, 1.72068e-005, 1.614186e-005, 
    1.507692e-005, 1.385304e-005, 1.269274e-005, 1.156424e-005, 1.04834e-005, 
    9.545616e-006, 8.591942e-006, 7.765429e-006, 7.097857e-006,
  1.488619e-005, 1.437757e-005, 1.393252e-005, 1.371e-005, 1.345569e-005, 
    1.324906e-005, 1.318548e-005, 1.291527e-005, 1.280401e-005, 
    1.248612e-005, 1.202517e-005, 1.140529e-005, 1.075361e-005, 
    9.815829e-006, 8.97342e-006, 7.797224e-006, 6.716393e-006, 5.699137e-006, 
    4.777253e-006, 4.014311e-006, 3.473896e-006, 3.028848e-006, 
    2.869901e-006, 2.981164e-006, 3.219584e-006, 3.569265e-006, 4.17326e-006, 
    4.888516e-006, 5.842189e-006, 6.795864e-006, 7.987956e-006, 
    9.211837e-006, 1.062646e-005, 1.22318e-005, 1.421863e-005, 1.630082e-005, 
    1.846247e-005, 2.083076e-005, 2.329443e-005, 2.588527e-005, 
    2.817406e-005, 3.041521e-005, 3.194108e-005, 3.413454e-005, 3.56286e-005, 
    3.529483e-005, 3.793332e-005, 3.923668e-005, 4.066718e-005, 
    4.163677e-005, 4.340106e-005, 4.678663e-005, 4.905957e-005, 
    5.309675e-005, 5.211133e-005, 6.051951e-005, 6.279245e-005, 
    6.373021e-005, 6.406399e-005, 6.268118e-005, 6.051955e-005, 
    5.734061e-005, 5.285833e-005, 4.775617e-005, 4.262224e-005, 
    3.791745e-005, 3.332391e-005, 2.949333e-005, 2.691841e-005, 2.48998e-005, 
    2.359644e-005, 2.327855e-005, 2.39779e-005, 2.559915e-005, 2.771313e-005, 
    3.031982e-005, 3.289476e-005, 3.599421e-005, 3.844197e-005, 
    4.085795e-005, 4.33216e-005, 4.373488e-005, 4.465676e-005, 4.311498e-005, 
    4.279708e-005, 4.07467e-005, 3.858503e-005, 3.591474e-005, 3.284708e-005, 
    2.946154e-005, 2.617136e-005, 2.326265e-005, 2.075132e-005, 
    1.863734e-005, 1.698428e-005, 1.579218e-005,
  1.243843e-005, 8.480685e-006, 5.794504e-006, 3.775895e-006, 2.234121e-006, 
    9.466603e-007, -1.500648e-007, -8.812131e-007, -1.135526e-006, 
    -9.76579e-007, -2.931156e-007, 8.830848e-007, 2.440749e-006, 
    3.998417e-006, 5.571981e-006, 6.923019e-006, 8.035639e-006, 
    8.703213e-006, 8.591951e-006, 7.876697e-006, 6.795863e-006, 
    5.317666e-006, 4.125573e-006, 3.23548e-006, 2.997058e-006, 3.251372e-006, 
    3.505686e-006, 4.07789e-006, 4.6342e-006, 5.206406e-006, 5.921662e-006, 
    6.621025e-006, 7.638278e-006, 8.830364e-006, 1.024498e-005, 
    1.208875e-005, 1.472725e-005, 1.8383e-005, 2.299242e-005, 2.871449e-005, 
    3.478621e-005, 3.98089e-005, 4.475213e-005, 4.847145e-005, 5.002912e-005, 
    5.249277e-005, 5.317623e-005, 5.368485e-005, 5.447958e-005, 
    5.541735e-005, 5.641869e-005, 5.772208e-005, 5.691146e-005, 5.72135e-005, 
    5.784931e-005, 5.905732e-005, 5.955005e-005, 5.940703e-005, 
    6.088521e-005, 6.174349e-005, 6.277664e-005, 6.419123e-005, 
    6.614625e-005, 6.76403e-005, 7.037417e-005, 7.423654e-005, 7.689091e-005, 
    7.884596e-005, 7.944995e-005, 7.852809e-005, 7.422063e-005, 
    6.857807e-005, 6.357129e-005, 5.929563e-005, 5.600548e-005, 
    5.292193e-005, 5.026754e-005, 4.990195e-005, 5.018806e-005, 
    5.060132e-005, 5.077616e-005, 5.091922e-005, 5.150729e-005, 5.28901e-005, 
    5.544914e-005, 5.956585e-005, 6.366665e-005, 6.735422e-005, 
    6.949995e-005, 6.940457e-005, 6.44773e-005, 5.625979e-005, 4.589652e-005, 
    3.516769e-005, 2.55038e-005, 1.787437e-005,
  1.444115e-005, 1.407557e-005, 1.467956e-005, 1.533124e-005, 1.531535e-005, 
    1.448883e-005, 1.307422e-005, 1.134171e-005, 9.291307e-006, 
    7.240909e-006, 5.746822e-006, 4.618305e-006, 4.01431e-006, 4.236839e-006, 
    5.142829e-006, 6.811753e-006, 9.354892e-006, 1.208875e-005, 
    1.420273e-005, 1.51723e-005, 1.405967e-005, 1.200928e-005, 9.704567e-006, 
    8.115112e-006, 7.463441e-006, 7.193225e-006, 6.779968e-006, 
    6.589235e-006, 6.493868e-006, 6.795865e-006, 7.09786e-006, 7.701852e-006, 
    8.369425e-006, 9.084679e-006, 9.927091e-006, 1.075361e-005, 
    1.191391e-005, 1.385304e-005, 1.645976e-005, 1.981351e-005, 
    2.424811e-005, 2.941384e-005, 3.486568e-005, 3.939566e-005, 
    4.252687e-005, 4.634156e-005, 6.633696e-005, 7.17729e-005, 8.191366e-005, 
    9.03855e-005, 9.389821e-005, 9.491551e-005, 9.60757e-005, 9.728369e-005, 
    9.739486e-005, 0.0001015751, 0.0001209982, 8.995616e-005, 9.197486e-005, 
    9.427959e-005, 9.604392e-005, 9.998583e-005, 9.979514e-005, 0.0001015911, 
    0.0001023859, 0.0001036892, 0.0001053423, 0.0001091888, 0.0001158168, 
    0.0001232236, 0.0001300901, 0.0001333007, 0.0001339524, 0.000133857, 
    0.0001328716, 0.0001313616, 0.0001310596, 0.0001316954, 0.0001322517, 
    0.000132506, 0.0001621654, 0.0001533121, 0.0001494497, 0.0001481146, 
    0.0001482576, 0.0001508167, 0.0001565864, 0.0001640568, 0.0001826535, 
    0.0001262595, 0.0001067886, 8.105533e-005, 5.665715e-005, 3.729753e-005, 
    2.421632e-005, 1.720683e-005,
  4.300369e-005, 3.635976e-005, 3.237024e-005, 2.688661e-005, 2.173676e-005, 
    1.843069e-005, 1.857375e-005, 2.119634e-005, 2.615545e-005, 
    3.025627e-005, 2.898469e-005, 2.313549e-005, 1.518818e-005, 9.45025e-006, 
    7.39986e-006, 8.957519e-006, 1.281991e-005, 1.792206e-005, 2.267453e-005, 
    2.297656e-005, 2.48521e-005, 2.548789e-005, 2.242023e-005, 1.820818e-005, 
    1.452062e-005, 1.248612e-005, 1.189802e-005, 1.216823e-005, 
    1.281991e-005, 1.369411e-005, 1.413915e-005, 1.440936e-005, 
    1.485441e-005, 1.601471e-005, 1.762006e-005, 1.8987e-005, 1.95592e-005, 
    1.955919e-005, 2.075129e-005, 2.466137e-005, 3.066951e-005, 
    3.737703e-005, 4.300371e-005, 4.534022e-005, 4.6882e-005, 5.225436e-005, 
    6.972248e-005, 8.407535e-005, 9.331011e-005, 9.392988e-005, 
    9.106874e-005, 8.423405e-005, 7.805094e-005, 7.965643e-005, 
    8.590298e-005, 9.826897e-005, 0.0001212048, 0.0001579531, 0.0002016313, 
    0.0002457704, 0.0002855545, 0.0003188856, 0.000340089, 0.0003556657, 
    0.0003684767, 0.0003799845, 0.0003955294, 0.0004095484, 0.0004250456, 
    0.0004351545, 0.0003937492, 0.0004298456, 0.0004325, 0.0004313238, 
    0.000423313, 0.0004050342, 0.0003556975, 0.0003420442, 0.0003293285, 
    0.0003207136, 0.0003431568, 0.0003110497, 0.0002845693, 0.0002682774, 
    0.0002667356, 0.0002737769, 0.0002840925, 0.0002872397, 0.0002814541, 
    0.0002696444, 0.0002632071, 0.0001707167, 0.0001328558, 0.0001000017, 
    7.132781e-005, 5.397094e-005,
  0.0004194982, 0.0003596233, 0.0002093722, 0.000161927, 0.0001205216, 
    9.396169e-005, 8.477463e-005, 9.24835e-005, 0.0001167546, 0.0001482418, 
    0.0001711776, 0.0001717657, 0.0001391023, 9.168875e-005, 5.223847e-005, 
    2.809459e-005, 1.795385e-005, 1.480673e-005, 1.952742e-005, 2.63462e-005, 
    3.376897e-005, 4.289242e-005, 4.759723e-005, 4.651639e-005, 
    4.165267e-005, 3.866448e-005, 3.999964e-005, 4.448192e-005, 
    4.915487e-005, 5.055363e-005, 4.497463e-005, 3.631206e-005, 
    2.807871e-005, 2.528126e-005, 2.885755e-005, 3.589883e-005, 
    4.106456e-005, 4.131888e-005, 3.721807e-005, 3.488157e-005, 
    3.581935e-005, 3.972941e-005, 4.287655e-005, 4.049236e-005, 
    3.764729e-005, 3.639163e-005, 3.799697e-005, 4.562619e-005, 
    4.799443e-005, 3.313308e-005, 5.190261e-006, -3.297464e-006, 
    8.766772e-006, 3.885524e-005, 8.712697e-005, 0.0001365909, 0.0001860865, 
    0.0002331663, 0.0002966492, 0.0003618806, 0.0004239011, 0.0004780063, 
    0.0005214462, 0.000576648, 0.00064207, 0.000713548, 0.0007790335, 
    0.0008534202, 0.0009246279, 0.0009873002, 0.001028849, 0.0009368508, 
    0.0009004839, 0.0008771667, 0.0008512425, 0.000795548, 0.0007094153, 
    0.0006136345, 0.0005181718, 0.0005049317, 0.0005425541, 0.0004972388, 
    0.0004429269, 0.0004020778, 0.0003928589, 0.0004179723, 0.0004598228, 
    0.0004956015, 0.0005193798, 0.0005437144, 0.0005790163, 0.0006238389, 
    0.0006510505, 0.0006286391, 0.0005631216, 0.0004843005,
  0.001426817, 0.001439119, 0.001423813, 0.001366004, 0.001329081, 
    0.00130206, 0.001268015, 0.001211128, 0.001148932, 0.001136948, 
    0.001184631, 0.001238498, 0.001239944, 0.001139825, 0.0009802432, 
    0.0007470696, 0.0005570341, 0.0004555472, 0.000434471, 0.0004607128, 
    0.00047292, 0.0004540689, 0.0004229156, 0.000378538, 0.0003236062, 
    0.0002772418, 0.0002484568, 0.0002533045, 0.0002659885, 0.0002695966, 
    0.0002571193, 0.00018437, 0.0001474943, 0.0001213956, 0.0001513887, 
    0.0001990724, 0.0004389692, 0.0005255311, 0.0005373249, 0.0004526228, 
    0.0003528207, 0.0003285338, 0.0003514696, 0.0003149757, 0.0002210388, 
    0.0001048653, 1.74134e-005, -2.685282e-005, -3.418047e-005, 
    -2.078107e-005, -1.261104e-005, -1.275423e-005, -9.384472e-006, 
    1.628511e-005, 4.286109e-005, 7.889397e-005, 0.0001160395, 0.0001590659, 
    0.0002238683, 0.0002727441, 0.0003014179, 0.0003202369, 0.0003540127, 
    0.0004022054, 0.000449762, 0.0004862561, 0.0005203974, 0.0005720232, 
    0.0006384465, 0.0006943636, 0.0007317634, 0.0007478329, 0.0007571152, 
    0.0007606281, 0.000756257, 0.0007402191, 0.0007197787, 0.0007492953, 
    0.0008626713, 0.0009797185, 0.0008279729, 0.0007618357, 0.0007089861, 
    0.0006770537, 0.0007337657, 0.0008062606, 0.0008807271, 0.0009293963, 
    0.0009528409, 0.0009830564, 0.00101394, 0.001068093, 0.001133991, 
    0.001207234, 0.001290569, 0.001367514,
  0.0009512356, 0.000910609, 0.0008722555, 0.0008287046, 0.0007924011, 
    0.0007681779, 0.0007379148, 0.0007102424, 0.0006800585, 0.0006516548, 
    0.000639877, 0.0006483488, 0.0006722384, 0.0006992433, 0.0007251191, 
    0.0007356256, 0.0007308573, 0.000717649, 0.0007091775, 0.0007134688, 
    0.0006997834, 0.0006575678, 0.0006023333, 0.0005247525, 0.0004403049, 
    0.0003749144, 0.000328534, 0.0002856345, 0.0002514296, 0.0002271743, 
    0.0002060025, 0.0001769317, 0.0001495455, 0.0001545835, 0.000180651, 
    0.0002250446, 0.0002908001, 0.0003471305, 0.0003666172, 0.0003790313, 
    0.0003917788, 0.0003934002, 0.0003702259, 0.0003403758, 0.0002880348, 
    0.0002027759, 9.022653e-005, -4.679896e-007, -1.207134e-005, 
    -1.97906e-007, 1.350325e-005, 1.531537e-005, 5.603768e-006, 
    8.401228e-006, 2.771383e-005, 4.872633e-005, 8.072215e-005, 0.0001224135, 
    0.000158526, 0.0001847197, 0.0002007573, 0.0002300194, 0.000279038, 
    0.0003238132, 0.0003592581, 0.0003934153, 0.0004520346, 0.0005249111, 
    0.0005899039, 0.0006326765, 0.0006572176, 0.0006825693, 0.0007229256, 
    0.0007528232, 0.0007590861, 0.0007525852, 0.0007363092, 0.0007106555, 
    0.0006741777, 0.0006282581, 0.0006050679, 0.0006233146, 0.0006106626, 
    0.000569623, 0.0006018253, 0.0006703627, 0.0007607075, 0.0008513222, 
    0.0009124053, 0.0009391876, 0.0009337994, 0.0009321144, 0.0009429865, 
    0.0009619964, 0.0009710402, 0.0009702933,
  0.0005629312, 0.0005476091, 0.0005409177, 0.0005284087, 0.0004979065, 
    0.0004720462, 0.0004575506, 0.0004538789, 0.0004600461, 0.0004617311, 
    0.0004623982, 0.0004664832, 0.0004763855, 0.0004959041, 0.0005239579, 
    0.0005453362, 0.0005586082, 0.0005653317, 0.0005645845, 0.0005475776, 
    0.0005016103, 0.0004560407, 0.0004339949, 0.0004227574, 0.0004121717, 
    0.0003989155, 0.0003951485, 0.0003881389, 0.0003769968, 0.0003636773, 
    0.0003543629, 0.0003307271, 0.0002890197, 0.0002687385, 0.0002671652, 
    0.0002701525, 0.0002744603, 0.0002979841, 0.0003207452, 0.000329487, 
    0.0003390084, 0.0003619287, 0.0003897594, 0.0003940035, 0.0003745169, 
    0.0003580023, 0.0003179, 0.000222215, 0.0001206649, 5.95185e-005, 
    5.055405e-005, 6.6448e-005, 6.791018e-005, 6.291969e-005, 6.508129e-005, 
    6.442983e-005, 5.486095e-005, 7.698592e-005, 0.0001324108, 0.0001735617, 
    0.0001855143, 0.0002212771, 0.0002663541, 0.0002860478, 0.0003176779, 
    0.0003920165, 0.0004962212, 0.0005876147, 0.0006552949, 0.0006923131, 
    0.0007136436, 0.0007537617, 0.0008089794, 0.0008546598, 0.0008728271, 
    0.000853674, 0.0008034953, 0.0007516788, 0.000722337, 0.000702756, 
    0.0006872267, 0.0006850013, 0.0006647515, 0.000539789, 0.0004789445, 
    0.0004670555, 0.0004833476, 0.0005098437, 0.0005325729, 0.0005486263, 
    0.0005595139, 0.0005710216, 0.0005875521, 0.0005962939, 0.0005920979, 
    0.0005773955,
  0.0005440488, 0.0005673503, 0.000595849, 0.0006013648, 0.0005806065, 
    0.0005508673, 0.0005388351, 0.0005281537, 0.0005060444, 0.0004889574, 
    0.0004939325, 0.0005202699, 0.0005494524, 0.0005654106, 0.0005811616, 
    0.0006245226, 0.0006800261, 0.0007194127, 0.0007099714, 0.0006543719, 
    0.0005995841, 0.000552393, 0.0005091755, 0.0004981286, 0.0005025472, 
    0.0005177585, 0.000566571, 0.0005932576, 0.0005711168, 0.0005326676, 
    0.0005098903, 0.0004901178, 0.000463272, 0.0004425934, 0.0004361398, 
    0.0004198635, 0.0003899983, 0.0003705113, 0.0003758045, 0.0004086741, 
    0.0004655765, 0.0005107652, 0.000543349, 0.0005498338, 0.0005806061, 
    0.0005573677, 0.0004650997, 0.0003891401, 0.0003009886, 0.0002304642, 
    0.0002001692, 0.0002124878, 0.0002104687, 0.0001834002, 0.0001560934, 
    0.0001490521, 0.0001715273, 0.0002122172, 0.0002434975, 0.0002553235, 
    0.0002672602, 0.0002969829, 0.0003332072, 0.0003514695, 0.0004088967, 
    0.0005058218, 0.0005938779, 0.0006481898, 0.0006789612, 0.0007177442, 
    0.0007706732, 0.0008126507, 0.0008445191, 0.0008768332, 0.0008975593, 
    0.0008672327, 0.0008536587, 0.0009188424, 0.0008829846, 0.0007700371, 
    0.0007339567, 0.0007084459, 0.0006570271, 0.0005610874, 0.0005125771, 
    0.0005006241, 0.0005269777, 0.0005385964, 0.0005359263, 0.0005331766, 
    0.0005431108, 0.0005639323, 0.000573803, 0.0005613263, 0.000542793, 
    0.0005354339,
  0.0006600628, 0.0006908509, 0.000736373, 0.000743255, 0.000722656, 
    0.000717029, 0.00071536, 0.0007143747, 0.0007124511, 0.0007083979, 
    0.0006979397, 0.0006967792, 0.0007086205, 0.0007101786, 0.0007195403, 
    0.0007784138, 0.0008670739, 0.0009128023, 0.0008752113, 0.0008174507, 
    0.0008349344, 0.000893347, 0.0009163152, 0.0009136926, 0.0009137876, 
    0.0009279819, 0.0009533656, 0.0009661284, 0.0009613289, 0.000943304, 
    0.0008708406, 0.0007721512, 0.0007259618, 0.0006834753, 0.000636078, 
    0.000592161, 0.0005585123, 0.0005493411, 0.0005607693, 0.0006068796, 
    0.000700451, 0.0007582116, 0.0007362613, 0.0007598801, 0.0008821576, 
    0.0008468074, 0.0006792475, 0.0005463213, 0.0004947432, 0.000450572, 
    0.0004319116, 0.0004625404, 0.0004686755, 0.0004366166, 0.0004178449, 
    0.0004273024, 0.0004685964, 0.0004911032, 0.0004748111, 0.0004681041, 
    0.0004849993, 0.0005002581, 0.0005036443, 0.0005254997, 0.0005695592, 
    0.0006180694, 0.0006695199, 0.0007237205, 0.0007758234, 0.0008494151, 
    0.0009192713, 0.0009618057, 0.0009733131, 0.0009808312, 0.0009654928, 
    0.000939203, 0.0009008655, 0.0008374932, 0.0008570123, 0.0009253277, 
    0.0008245879, 0.0006940453, 0.0006486187, 0.0006020796, 0.0005775858, 
    0.0006410847, 0.0006997832, 0.0006929962, 0.0006705849, 0.0006515118, 
    0.0006386363, 0.0006391769, 0.0006544841, 0.0006585531, 0.0006615729, 
    0.0006609689,
  0.0009110696, 0.0009611859, 0.0009798296, 0.0009755702, 0.001016022, 
    0.001082032, 0.001153081, 0.001210826, 0.001190703, 0.001163873, 
    0.00118282, 0.001202052, 0.001186014, 0.00115707, 0.001137377, 
    0.001143862, 0.001201225, 0.001289901, 0.001292461, 0.001384887, 
    0.001538889, 0.001589212, 0.001468413, 0.00129087, 0.00115804, 
    0.001081952, 0.001019042, 0.0009734086, 0.0009549391, 0.0009104502, 
    0.0008535949, 0.00083174, 0.0008539767, 0.0008777068, 0.0008902475, 
    0.0008776113, 0.0008577751, 0.0008593164, 0.0008898983, 0.000948438, 
    0.001078122, 0.001132513, 0.001082064, 0.001097911, 0.00119873, 
    0.00112768, 0.0009918143, 0.0008840016, 0.0008264631, 0.0007782546, 
    0.0008160518, 0.0008809338, 0.000906969, 0.0008580773, 0.0008160206, 
    0.0007978845, 0.0007697036, 0.0007371036, 0.0007249448, 0.0007232595, 
    0.000713564, 0.0007027872, 0.000713103, 0.0007535866, 0.0007673511, 
    0.0007684953, 0.0007885867, 0.0008604769, 0.0009493916, 0.001009298, 
    0.001024826, 0.001041516, 0.001057141, 0.001035047, 0.001023635, 
    0.001003593, 0.0009151548, 0.0007862975, 0.0008065631, 0.0009824997, 
    0.0009146933, 0.0007526958, 0.0007033432, 0.0006620171, 0.0006703301, 
    0.0007887608, 0.0009055701, 0.0009194459, 0.0008864966, 0.0008554547, 
    0.0008371123, 0.0008397987, 0.0008430574, 0.0008190563, 0.0008270987, 
    0.0008730185,
  0.001246747, 0.00126927, 0.001284735, 0.00131244, 0.001411748, 0.001584825, 
    0.001782935, 0.001946887, 0.002057768, 0.00215854, 0.002188643, 
    0.002102653, 0.001894022, 0.00171597, 0.001629027, 0.001613164, 
    0.001610144, 0.001634304, 0.001679396, 0.001732707, 0.00172867, 
    0.001565116, 0.001283352, 0.001017993, 0.0008370969, 0.000809567, 
    0.0009125955, 0.001000794, 0.001006358, 0.001030454, 0.001060909, 
    0.001073847, 0.00110287, 0.001104491, 0.001111453, 0.001140143, 
    0.001145117, 0.001176159, 0.001212494, 0.001321245, 0.001507322, 
    0.001533787, 0.001473992, 0.001458271, 0.001465408, 0.001480842, 
    0.001205199, 0.001339715, 0.001354941, 0.001409762, 0.001479031, 
    0.00145673, 0.00136931, 0.001278329, 0.00122033, 0.001131003, 
    0.001054456, 0.001014004, 0.0009989035, 0.0009577046, 0.0009153462, 
    0.0009343075, 0.0009572431, 0.0009185239, 0.0008846205, 0.0009156624, 
    0.0009612171, 0.001004244, 0.001065104, 0.001111468, 0.00114545, 
    0.001193389, 0.001191879, 0.001128714, 0.001054947, 0.00102346, 
    0.0009182058, 0.0006348859, 0.0006654034, 0.0009944211, 0.001006898, 
    0.0009664157, 0.001011905, 0.001038734, 0.001033378, 0.001032648, 
    0.001074799, 0.001082603, 0.00105784, 0.001060893, 0.001072591, 
    0.001102822, 0.001109164, 0.001081825, 0.001140397, 0.001217088,
  0.001427279, 0.001427692, 0.001393851, 0.001431745, 0.001605583, 
    0.001810368, 0.001931041, 0.002121887, 0.002142979, 0.002175611, 
    0.002013693, 0.001766992, 0.001574271, 0.001470416, 0.001411177, 
    0.001399686, 0.001381788, 0.001366116, 0.001337457, 0.001286405, 
    0.001218027, 0.001136232, 0.00108467, 0.001108845, 0.001179243, 
    0.001222953, 0.00126048, 0.001306876, 0.001314823, 0.001376351, 
    0.00136583, 0.001312917, 0.001274499, 0.001222254, 0.00124797, 
    0.001316858, 0.001360743, 0.001418218, 0.001345898, 0.001212415, 
    0.001731007, 0.002014121, 0.001982015, 0.001832113, 0.001790183, 
    0.001783078, 0.001740751, 0.00130322, 0.001546137, 0.00151945, 
    0.001416327, 0.001374635, 0.001341908, 0.001339191, 0.001327826, 
    0.001262389, 0.001216326, 0.001198286, 0.001181358, 0.00116896, 
    0.001129207, 0.001086673, 0.001104522, 0.001110181, 0.001136551, 
    0.001185521, 0.001210777, 0.001274245, 0.001312441, 0.001288916, 
    0.001269081, 0.001209412, 0.001157644, 0.00109168, 0.001047651, 
    0.0009974884, 0.0007528076, 0.0004136967, 0.0005906038, 0.0009491844, 
    0.001104173, 0.001271305, 0.001579803, 0.00166514, 0.001555276, 
    0.001367021, 0.001278568, 0.001276073, 0.001283529, 0.001291301, 
    0.001261783, 0.001222841, 0.001221459, 0.001234811, 0.001303237, 
    0.001387811,
  0.001538508, 0.001495291, 0.001407568, 0.00144082, 0.001626771, 
    0.001803264, 0.002086219, 0.002067003, 0.002005857, 0.00203496, 
    0.00153897, 0.001430585, 0.001409636, 0.001409207, 0.001395632, 
    0.001367515, 0.001362348, 0.001365321, 0.001348807, 0.001309515, 
    0.001305573, 0.00142464, 0.001538938, 0.001565211, 0.001597891, 
    0.00161806, 0.001556278, 0.001523106, 0.001471337, 0.001405646, 
    0.001315412, 0.001259305, 0.001247177, 0.001272307, 0.001395967, 
    0.001479079, 0.001381184, 0.001324137, 0.001301282, 0.001339571, 
    0.001660021, 0.002281866, 0.002453686, 0.002248805, 0.002052682, 
    0.00199349, 0.001870514, 0.001707181, 0.001545598, 0.00133528, 
    0.001330019, 0.00140803, 0.001452645, 0.001524759, 0.001537587, 
    0.001482782, 0.001473356, 0.001449783, 0.001396807, 0.001410303, 
    0.001444889, 0.001415341, 0.001459464, 0.001521405, 0.001544787, 
    0.001517924, 0.001430727, 0.0013421, 0.001255602, 0.001134151, 
    0.001029009, 0.0009319233, 0.0008900734, 0.0008639423, 0.0007949602, 
    0.0007758383, 0.0005884264, 0.0005330965, 0.0007960568, 0.001121514, 
    0.001227737, 0.001583379, 0.002032878, 0.002090718, 0.001945585, 
    0.001740481, 0.001619348, 0.001549381, 0.001462231, 0.001437768, 
    0.001429344, 0.001406647, 0.001436338, 0.001456158, 0.001469111, 
    0.001522406,
  0.00132522, 0.001318481, 0.001281001, 0.001483387, 0.001594617, 
    0.001117032, 0.001170135, 0.001638087, 0.001967184, 0.002043192, 
    0.001849628, 0.001851949, 0.00189558, 0.001793871, 0.001796669, 
    0.001871644, 0.001892689, 0.001869164, 0.001823388, 0.001832511, 
    0.001871485, 0.001926923, 0.001949192, 0.001912825, 0.001833671, 
    0.001751797, 0.001642697, 0.001526523, 0.001473356, 0.001426611, 
    0.001345437, 0.001112485, 0.001155481, 0.001052421, 0.0009700544, 
    0.001045713, 0.00110082, 0.001213178, 0.001648387, 0.00206271, 
    0.002185209, 0.002374468, 0.00215479, 0.002089892, 0.001993761, 
    0.001882467, 0.001829443, 0.001711632, 0.001683261, 0.001734807, 
    0.001822163, 0.001846785, 0.001818778, 0.00183232, 0.00184866, 
    0.001852458, 0.001862266, 0.001840888, 0.001804728, 0.001818476, 
    0.001840569, 0.001858101, 0.001870102, 0.001826932, 0.001708422, 
    0.001470067, 0.001202545, 0.0009755539, 0.0008947309, 0.0008940641, 
    0.0008764686, 0.0008792663, 0.0008123498, 0.000737343, 0.0006158929, 
    0.0007007373, 0.0007820064, 0.0006664358, 0.001003704, 0.001495592, 
    0.001565592, 0.001978152, 0.002253748, 0.002432482, 0.002341534, 
    0.00212621, 0.001994588, 0.001906183, 0.001778072, 0.001647132, 
    0.001581774, 0.001532597, 0.001533233, 0.001515827, 0.001440709, 
    0.001386271,
  0.001273006, 0.001350333, 0.001555612, 0.001917435, 0.00200112, 
    0.0009458135, 0.001008646, 0.001607219, 0.001928164, 0.002164054, 
    0.002059024, 0.002212344, 0.002301241, 0.002202155, 0.002204888, 
    0.002354249, 0.002468118, 0.002420212, 0.002388931, 0.002348211, 
    0.002300161, 0.002195114, 0.00207743, 0.002004125, 0.001921091, 
    0.001792552, 0.001712745, 0.001691447, 0.001815964, 0.00197901, 
    0.001977946, 0.001699393, 0.001715763, 0.001406536, 0.0008166395, 
    0.0009526019, 0.001519944, 0.001990979, 0.002344171, 0.002471438, 
    0.002516549, 0.00238275, 0.002224804, 0.002225662, 0.002193746, 
    0.002138496, 0.002147175, 0.002088063, 0.002067479, 0.002099968, 
    0.002101685, 0.002114639, 0.002124971, 0.002158348, 0.002156712, 
    0.002220131, 0.002261044, 0.002308283, 0.002276334, 0.002194462, 
    0.002119614, 0.002081579, 0.002020845, 0.00185516, 0.001580104, 
    0.001209268, 0.001019296, 0.0008963514, 0.0008949684, 0.0008994825, 
    0.0008801073, 0.0009371368, 0.0007877452, 0.0007159496, 0.0006871959, 
    0.0009295717, 0.001350429, 0.0005960553, 0.001234667, 0.002079369, 
    0.002132758, 0.002207335, 0.002355727, 0.002463445, 0.002608674, 
    0.002333189, 0.002150957, 0.002015694, 0.00191006, 0.001792027, 
    0.001716495, 0.001623147, 0.00154833, 0.001475201, 0.001402452, 
    0.001282241,
  0.001671704, 0.001861216, 0.002235454, 0.002516993, 0.001611797, 
    0.001069761, 0.001386763, 0.001751876, 0.00200991, 0.00216164, 
    0.002286843, 0.002429432, 0.002513021, 0.002561437, 0.002614366, 
    0.00256007, 0.002609185, 0.00259866, 0.002617145, 0.002587215, 
    0.002483028, 0.002371972, 0.00227643, 0.002273028, 0.002274554, 
    0.002258691, 0.002289193, 0.002425441, 0.002570431, 0.002753428, 
    0.002789792, 0.002345731, 0.002093895, 0.001713714, 0.001881163, 
    0.002037788, 0.00213449, 0.002547939, 0.002644992, 0.002705377, 
    0.002721382, 0.002607752, 0.002806976, 0.002846409, 0.002656883, 
    0.002486412, 0.002434311, 0.002368951, 0.00230604, 0.002268497, 
    0.00232766, 0.002412998, 0.002510209, 0.002610567, 0.002631135, 
    0.002655008, 0.002702342, 0.002703996, 0.002569783, 0.002486192, 
    0.002349945, 0.002169143, 0.002007082, 0.001779551, 0.00153733, 
    0.001243584, 0.001222221, 0.001224685, 0.001138537, 0.001073989, 
    0.001032171, 0.001012827, 0.0009197174, 0.0009204159, 0.0009170631, 
    0.001319815, 0.002110762, 0.001015339, 0.001249068, 0.00256285, 
    0.002516073, 0.0021501, 0.002225408, 0.002169125, 0.002199215, 
    0.002264638, 0.002189107, 0.002035419, 0.001950575, 0.001852585, 
    0.001787719, 0.001710663, 0.001639503, 0.00158972, 0.001566292, 
    0.001506433,
  0.002264858, 0.002454655, 0.002770433, 0.002689451, 0.001783618, 
    0.00161663, 0.001955344, 0.001950177, 0.001915353, 0.002137669, 
    0.002588267, 0.002758449, 0.002452765, 0.002512194, 0.002800364, 
    0.002667643, 0.002681712, 0.002686718, 0.002712784, 0.002823649, 
    0.002880823, 0.002805561, 0.002749834, 0.00279903, 0.002857553, 
    0.002889421, 0.002989257, 0.003106048, 0.00320779, 0.003362205, 
    0.003374223, 0.003091091, 0.002564057, 0.002073217, 0.002300335, 
    0.002076237, 0.002292259, 0.002840417, 0.003022918, 0.002859062, 
    0.002986299, 0.003076279, 0.003219329, 0.003138395, 0.002956798, 
    0.002790399, 0.002723133, 0.00266186, 0.002603717, 0.002624029, 
    0.002768399, 0.002881536, 0.002992306, 0.003142796, 0.003162744, 
    0.00312075, 0.003086004, 0.00302214, 0.002918778, 0.002838319, 
    0.002593957, 0.002312129, 0.002132013, 0.001942804, 0.001853509, 
    0.001678765, 0.001546567, 0.001399367, 0.001348313, 0.001310675, 
    0.001264836, 0.001237958, 0.00122227, 0.00122238, 0.001261926, 
    0.001813055, 0.00242347, 0.001673421, 0.001762129, 0.002766158, 
    0.002496808, 0.002361864, 0.002638875, 0.001996431, 0.001855335, 
    0.002177439, 0.002254862, 0.002236376, 0.002149846, 0.001996162, 
    0.001912906, 0.001871849, 0.001867891, 0.001877619, 0.00196124, 
    0.002026313,
  0.00270986, 0.002881681, 0.003063675, 0.002822347, 0.001942708, 
    0.001699028, 0.001982285, 0.002005936, 0.002219797, 0.002156634, 
    0.002491498, 0.003061749, 0.002666086, 0.002542965, 0.0028027, 
    0.002823886, 0.002862496, 0.002875783, 0.00294273, 0.003011204, 
    0.003071303, 0.00306933, 0.003120925, 0.003238212, 0.003286166, 
    0.003349505, 0.003506448, 0.003579816, 0.003597237, 0.003610002, 
    0.003641583, 0.003657367, 0.003484562, 0.003510755, 0.003455872, 
    0.002790396, 0.002900516, 0.003321119, 0.003022967, 0.003107496, 
    0.003208457, 0.003345165, 0.0034148, 0.003345437, 0.003246477, 
    0.003122373, 0.003088165, 0.003004638, 0.002907474, 0.002946878, 
    0.003067805, 0.003144717, 0.003255645, 0.003309639, 0.003238957, 
    0.003200395, 0.003143542, 0.00304633, 0.002983753, 0.002867961, 
    0.002731396, 0.002633311, 0.002510985, 0.002319075, 0.002228891, 
    0.002126053, 0.002000135, 0.001909026, 0.001880177, 0.001834082, 
    0.001847371, 0.001821049, 0.001798686, 0.001781314, 0.001899697, 
    0.002340694, 0.002001502, 0.002126813, 0.00224553, 0.002963267, 
    0.002575994, 0.002428493, 0.002322619, 0.002182843, 0.002002853, 
    0.002078971, 0.00239877, 0.002412235, 0.002354728, 0.002285063, 
    0.002335543, 0.002360308, 0.00244431, 0.002418528, 0.002541426, 
    0.002573976,
  0.003074847, 0.003170261, 0.003215991, 0.003104616, 0.002234755, 
    0.001615152, 0.002081483, 0.00192408, 0.002004283, 0.001980742, 
    0.002271486, 0.003237989, 0.003185648, 0.002933497, 0.002960071, 
    0.002967685, 0.003052784, 0.003017608, 0.003168114, 0.003250083, 
    0.003331067, 0.003363682, 0.003426051, 0.003481602, 0.003545228, 
    0.003703397, 0.003762349, 0.003789021, 0.003833571, 0.003825482, 
    0.003838293, 0.003920849, 0.00398376, 0.003837278, 0.003584236, 
    0.003183391, 0.003411971, 0.003463453, 0.00310554, 0.003275516, 
    0.003419043, 0.003558487, 0.003562411, 0.003497846, 0.003381848, 
    0.003268074, 0.003166858, 0.003060063, 0.002978824, 0.002960054, 
    0.002997709, 0.003034584, 0.003130443, 0.003134511, 0.003025698, 
    0.003027575, 0.003053911, 0.002995294, 0.003012268, 0.002950598, 
    0.002924642, 0.002867835, 0.002767446, 0.002694648, 0.002626937, 
    0.002569908, 0.002532223, 0.002490563, 0.00248233, 0.002518618, 
    0.002511227, 0.002393734, 0.002369128, 0.002456724, 0.002655549, 
    0.003105587, 0.002563995, 0.00222641, 0.002493486, 0.00246459, 
    0.002084916, 0.001650693, 0.002119074, 0.002419147, 0.001867304, 
    0.002120886, 0.002528582, 0.00264005, 0.002671998, 0.002723005, 
    0.002787188, 0.002841832, 0.002945673, 0.002917919, 0.003022872, 
    0.003049115,
  0.003239324, 0.003207088, 0.003138201, 0.003227146, 0.002870236, 
    0.002478594, 0.002642721, 0.002631197, 0.002511336, 0.002387136, 
    0.002346016, 0.003052751, 0.003021648, 0.002930811, 0.003018307, 
    0.002982847, 0.003107127, 0.003133925, 0.003219899, 0.003276419, 
    0.003415864, 0.003422124, 0.003451323, 0.003496353, 0.003487818, 
    0.003502838, 0.003425051, 0.003475515, 0.003424654, 0.003592959, 
    0.003830791, 0.003720371, 0.003726428, 0.003760394, 0.003723821, 
    0.003586523, 0.00345269, 0.003321068, 0.003052691, 0.003301803, 
    0.003548773, 0.003622111, 0.00357678, 0.003513439, 0.003370071, 
    0.003173534, 0.003040085, 0.003042404, 0.003011107, 0.002840512, 
    0.002843166, 0.002837013, 0.002864067, 0.002942156, 0.002958639, 
    0.00290614, 0.002940122, 0.002892375, 0.00290061, 0.002910368, 
    0.002934845, 0.002928821, 0.002936339, 0.002891343, 0.002902422, 
    0.002914963, 0.002917664, 0.002950042, 0.002958594, 0.00300391, 
    0.002973568, 0.002962807, 0.002996361, 0.003114423, 0.003102073, 
    0.002915648, 0.001992999, 0.001764322, 0.002023802, 0.002095534, 
    0.001714922, 0.001808795, 0.001932455, 0.002413284, 0.002346938, 
    0.002076984, 0.002485381, 0.002909446, 0.003030801, 0.003076434, 
    0.003131321, 0.003253296, 0.003290012, 0.003309118, 0.003314251, 
    0.003280396,
  0.003179289, 0.003109528, 0.002981449, 0.002987441, 0.003173728, 
    0.003077646, 0.003446956, 0.003222665, 0.003110227, 0.002519872, 
    0.002412646, 0.002850255, 0.003026778, 0.002930108, 0.003021343, 
    0.003077785, 0.003137691, 0.003263259, 0.003376968, 0.003451642, 
    0.003516382, 0.003495956, 0.003407422, 0.0033633, 0.003335485, 
    0.003283748, 0.00321966, 0.003158817, 0.003226114, 0.003322275, 
    0.003359802, 0.003358547, 0.003321115, 0.003251115, 0.003321147, 
    0.003328443, 0.003148612, 0.002838194, 0.002633058, 0.003097925, 
    0.003477296, 0.003434157, 0.003321448, 0.003257886, 0.003166111, 
    0.003017465, 0.002942666, 0.003008215, 0.003069187, 0.002983339, 
    0.003019199, 0.002986073, 0.002997883, 0.003049763, 0.00307928, 
    0.003033949, 0.003019676, 0.002965443, 0.002954364, 0.002897238, 
    0.002915392, 0.002948357, 0.003005115, 0.003010171, 0.003084905, 
    0.003133146, 0.003119273, 0.003106555, 0.003125472, 0.003171835, 
    0.003144003, 0.00312404, 0.003083922, 0.003108654, 0.00308292, 
    0.002974042, 0.002280816, 0.002760801, 0.00276937, 0.00229587, 
    0.002007796, 0.002086921, 0.00252248, 0.002748612, 0.00276662, 
    0.002597375, 0.002720732, 0.002921861, 0.003051765, 0.003082348, 
    0.003143031, 0.003307654, 0.003286799, 0.003347343, 0.003271349, 
    0.003242388,
  0.003071506, 0.00311099, 0.003083922, 0.002429526, 0.002754746, 
    0.003167098, 0.003247892, 0.003016928, 0.002861603, 0.002612599, 
    0.002641261, 0.003023062, 0.002845421, 0.002938883, 0.002976999, 
    0.003230944, 0.003374601, 0.003483018, 0.003446206, 0.003501169, 
    0.003512392, 0.003530527, 0.003535565, 0.003407836, 0.003306651, 
    0.00316616, 0.003131222, 0.002873844, 0.003124103, 0.003305761, 
    0.002594832, 0.003021507, 0.002947675, 0.003067628, 0.003194308, 
    0.003228879, 0.002948929, 0.002825461, 0.002968941, 0.003175568, 
    0.003283111, 0.003089722, 0.002984786, 0.002965696, 0.002982497, 
    0.002904756, 0.002860285, 0.002838159, 0.00290045, 0.002921764, 
    0.002968365, 0.00303112, 0.003105426, 0.003129171, 0.003184009, 
    0.00318579, 0.003182499, 0.003194483, 0.003224604, 0.003187506, 
    0.003193974, 0.00314448, 0.003157545, 0.003198361, 0.003170023, 
    0.003193086, 0.003198775, 0.00318433, 0.003227463, 0.003172327, 
    0.0031032, 0.003016576, 0.002978157, 0.0028644, 0.002865322, 0.003204532, 
    0.002809979, 0.003175555, 0.003082747, 0.002808994, 0.00272488, 
    0.002451938, 0.002456009, 0.003116205, 0.003069697, 0.002976665, 
    0.002939628, 0.003077865, 0.003225509, 0.003205243, 0.003164252, 
    0.00319113, 0.003173631, 0.003190778, 0.003151838, 0.003142556,
  0.003162201, 0.003217658, 0.003151393, 0.002422806, 0.002451733, 
    0.002990654, 0.002726914, 0.002669027, 0.00304549, 0.003152716, 
    0.002991577, 0.00310762, 0.003046934, 0.003073128, 0.003335245, 
    0.003500739, 0.003521625, 0.003537266, 0.003535787, 0.003542272, 
    0.003561029, 0.003564032, 0.003634732, 0.003634444, 0.003576636, 
    0.003190033, 0.003205387, 0.003089488, 0.003124198, 0.003178302, 
    0.003090279, 0.00299841, 0.002816433, 0.002963105, 0.003027303, 
    0.003001427, 0.003004782, 0.002932874, 0.003021931, 0.003012776, 
    0.002927503, 0.002881391, 0.003003065, 0.002930522, 0.002814395, 
    0.002811376, 0.002847107, 0.002838952, 0.002883045, 0.002888178, 
    0.002881614, 0.00292607, 0.002948005, 0.002952758, 0.002979398, 
    0.002997486, 0.003050113, 0.003057489, 0.003078613, 0.003139777, 
    0.003173107, 0.003173949, 0.003187444, 0.00316966, 0.003162824, 
    0.003222937, 0.003216626, 0.003186841, 0.003229562, 0.003122974, 
    0.003075736, 0.00296231, 0.002863605, 0.00270207, 0.002679691, 
    0.002996344, 0.002844648, 0.003091427, 0.003086435, 0.002745433, 
    0.00291676, 0.002221355, 0.002100859, 0.002847617, 0.002862256, 
    0.002973692, 0.002969401, 0.00310096, 0.003258936, 0.003206134, 
    0.003214383, 0.003147595, 0.00322176, 0.003240386, 0.003234522, 
    0.003208041,
  0.003120067, 0.003323849, 0.002887497, 0.003029643, 0.00335367, 
    0.003440805, 0.003276851, 0.0031022, 0.00319412, 0.003326807, 
    0.003297659, 0.00320555, 0.003217993, 0.003158387, 0.003360853, 
    0.003580833, 0.003721561, 0.003668237, 0.003644871, 0.003576303, 
    0.003571089, 0.003599364, 0.003593849, 0.003543273, 0.003559614, 
    0.003196757, 0.00307321, 0.003128285, 0.002972897, 0.002964679, 
    0.003094841, 0.00314022, 0.003021376, 0.00302886, 0.003018944, 
    0.002985025, 0.003019197, 0.003008883, 0.003026254, 0.003016654, 
    0.003086224, 0.003052307, 0.003132781, 0.003170514, 0.003166668, 
    0.00317595, 0.003172882, 0.003205705, 0.003233537, 0.003211649, 
    0.003179049, 0.003122656, 0.003081935, 0.003022345, 0.002951026, 
    0.002919888, 0.002904885, 0.002869248, 0.002881091, 0.002946496, 
    0.00296708, 0.002984961, 0.003040895, 0.003084382, 0.003201205, 
    0.003230419, 0.003290487, 0.003322022, 0.003330573, 0.003330048, 
    0.003254564, 0.003218994, 0.003174378, 0.002889881, 0.002891485, 
    0.002967481, 0.002776458, 0.002963729, 0.002919717, 0.001906786, 
    0.002296124, 0.002669647, 0.002830166, 0.002784166, 0.002810042, 
    0.002856694, 0.002824252, 0.002884857, 0.002971787, 0.002993848, 
    0.003041403, 0.002996992, 0.003131095, 0.003153348, 0.002725357, 
    0.002860524,
  0.003149835, 0.00312992, 0.003248114, 0.003289996, 0.003344309, 
    0.003569389, 0.003472671, 0.003254391, 0.003445188, 0.00334809, 
    0.002924562, 0.003127745, 0.003318414, 0.003414068, 0.003540063, 
    0.003673784, 0.003839215, 0.003820809, 0.003794709, 0.003769074, 
    0.003601829, 0.003455536, 0.003515935, 0.003562061, 0.003451133, 
    0.003279136, 0.003389351, 0.003203893, 0.003182229, 0.003046965, 
    0.003065785, 0.00296228, 0.003122037, 0.002967447, 0.002953062, 
    0.002997629, 0.002994878, 0.003085859, 0.003171578, 0.003276404, 
    0.003283381, 0.003242994, 0.003230579, 0.003312502, 0.003352666, 
    0.003371311, 0.003321784, 0.003309147, 0.00332935, 0.003297528, 
    0.003279582, 0.003257822, 0.00326631, 0.003202969, 0.00312542, 0.0030524, 
    0.002983404, 0.002891516, 0.002834359, 0.002779683, 0.002812553, 
    0.002784958, 0.002860697, 0.00293839, 0.003042674, 0.003129825, 
    0.003308002, 0.003389604, 0.003446762, 0.003401924, 0.003348328, 
    0.003440833, 0.003128981, 0.003005147, 0.002871428, 0.00274354, 
    0.002813747, 0.002693696, 0.002577489, 0.002566077, 0.002863513, 
    0.002789857, 0.002740964, 0.00264366, 0.002594052, 0.002653005, 
    0.002690818, 0.002709812, 0.00278059, 0.002846552, 0.002878565, 
    0.002934193, 0.002867864, 0.002741762, 0.003081951, 0.003148928,
  0.003657876, 0.003517432, 0.003167082, 0.002907446, 0.002377266, 
    0.00245329, 0.002177883, 0.002318279, 0.002624156, 0.002514374, 
    0.00202199, 0.001310803, 0.001718594, 0.002761452, 0.003707306, 
    0.003672529, 0.003684465, 0.003777957, 0.003715046, 0.003732625, 
    0.003596747, 0.003883721, 0.003787538, 0.003657347, 0.003539886, 
    0.003238065, 0.003175855, 0.003216451, 0.003225034, 0.003079168, 
    0.003032168, 0.00293548, 0.00291547, 0.003185598, 0.002823504, 
    0.00297606, 0.003010424, 0.003164997, 0.003196597, 0.003230531, 
    0.003147213, 0.003198218, 0.003214875, 0.003250115, 0.003232598, 
    0.003274847, 0.003261942, 0.003233761, 0.003192833, 0.003116349, 
    0.003056869, 0.002995024, 0.002995182, 0.002950439, 0.002928872, 
    0.00288392, 0.002864022, 0.002769036, 0.002759818, 0.002745211, 
    0.002766684, 0.002712166, 0.002720604, 0.00267165, 0.002694823, 
    0.002778411, 0.002872601, 0.003178285, 0.003569311, 0.003426863, 
    0.003423827, 0.003328951, 0.002793623, 0.002382148, 0.002725294, 
    0.002587218, 0.002559815, 0.002464829, 0.002531316, 0.002617354, 
    0.002555158, 0.002454691, 0.002466578, 0.00239135, 0.002407005, 
    0.002417576, 0.00244423, 0.002455436, 0.002502151, 0.002548482, 
    0.002682585, 0.002865674, 0.00300944, 0.003639709, 0.003984986, 
    0.003887076,
  0.002923276, 0.002739551, 0.00227144, 0.001855621, 0.001104539, 
    0.001002162, 0.0009570853, 0.0006844928, 0.0007680813, 0.001118972, 
    0.002234151, 0.002393733, 0.0001719571, 0.0008831746, 0.002207399, 
    0.003476677, 0.003524629, 0.003473658, 0.003570931, 0.003730195, 
    0.003451072, 0.004169141, 0.003979277, 0.003645187, 0.00354162, 
    0.003294555, 0.002793116, 0.003344083, 0.00333396, 0.002964457, 
    0.002874302, 0.002802713, 0.002672505, 0.002612518, 0.002673667, 
    0.002859266, 0.002935704, 0.003026778, 0.003049923, 0.003090946, 
    0.002954364, 0.002969671, 0.002967987, 0.002981879, 0.002972661, 
    0.002954938, 0.002935132, 0.002913134, 0.00283101, 0.002743049, 
    0.00266294, 0.002596945, 0.002563249, 0.002497795, 0.002503025, 
    0.002436966, 0.002395529, 0.002309538, 0.002273186, 0.002232354, 
    0.002266941, 0.002282009, 0.002270247, 0.002190568, 0.002075254, 
    0.001905102, 0.002014965, 0.002461394, 0.002933273, 0.003082175, 
    0.00312002, 0.002929174, 0.002262443, 0.002727121, 0.002722591, 
    0.002451716, 0.002394065, 0.002291054, 0.00225305, 0.002201965, 
    0.002254434, 0.002234804, 0.002266751, 0.002219622, 0.002292864, 
    0.002242638, 0.002221831, 0.002157411, 0.002106277, 0.002045561, 
    0.002234006, 0.002452398, 0.002251429, 0.001781345, 0.002371256, 
    0.002766872,
  0.001758217, 0.001847069, 0.001258001, 0.001490157, 0.0004237583, 
    0.0009869509, 0.0007218928, 0.0003292011, 0.0004953477, 0.001080522, 
    0.002372831, 0.001266695, 0.0005272478, 0.00023172, 0.000523719, 
    0.002007287, 0.00342262, 0.003410429, 0.003457144, 0.00354485, 
    0.003159264, 0.003757425, 0.004233912, 0.003699167, 0.003216052, 
    0.002937896, 0.002502418, 0.002907619, 0.003054725, 0.002919316, 
    0.002757493, 0.002763994, 0.002718458, 0.002655324, 0.002528612, 
    0.002708538, 0.002731776, 0.002762772, 0.002756158, 0.002756827, 
    0.002670122, 0.002669344, 0.002708748, 0.002681568, 0.002622614, 
    0.002615303, 0.002571911, 0.002576586, 0.002534861, 0.002429386, 
    0.002301417, 0.002169588, 0.002112445, 0.00207832, 0.002115576, 
    0.002012755, 0.001928895, 0.00187258, 0.001778945, 0.001690603, 
    0.001659721, 0.001627614, 0.001670832, 0.001691844, 0.00161544, 
    0.001363302, 0.00151314, 0.002038743, 0.001959206, 0.002465861, 
    0.002884891, 0.002726915, 0.002218463, 0.00278803, 0.002663622, 
    0.002468405, 0.002303069, 0.00210415, 0.002006622, 0.001995718, 
    0.001994843, 0.001936365, 0.002049519, 0.002048216, 0.002052651, 
    0.00202059, 0.001989024, 0.001880115, 0.001808254, 0.001700141, 
    0.00179546, 0.002086617, 0.00132053, 0.0006994815, 0.000587313, 
    0.001104268,
  0.00192643, 0.001793535, 0.001101264, 0.0008398308, 0.0008935062, 
    0.0007931162, 0.0001022746, 0.0001857372, 0.0001466523, 0.0007169815, 
    0.001764434, 0.0006493023, 0.0009467532, 0.000527184, 0.0001393091, 
    0.0009647938, 0.002971025, 0.003240356, 0.002592192, 0.003041897, 
    0.002995263, 0.003330369, 0.004412918, 0.004058165, 0.003216563, 
    0.003330113, 0.002690499, 0.00274853, 0.002680488, 0.002606673, 
    0.002594275, 0.003150791, 0.002573309, 0.002629114, 0.002403747, 
    0.002353597, 0.002414061, 0.002509318, 0.002469519, 0.0025272, 
    0.002596961, 0.00258272, 0.002539741, 0.002498781, 0.002427066, 
    0.00234505, 0.002256691, 0.002196909, 0.00216129, 0.002111015, 
    0.00207743, 0.001953403, 0.001814931, 0.001744343, 0.001734457, 
    0.001690254, 0.001614007, 0.001609828, 0.001546679, 0.001456413, 
    0.001361602, 0.001296706, 0.001387383, 0.001364987, 0.001354831, 
    0.001264693, 0.001480144, 0.002037327, 0.00232262, 0.002618624, 
    0.002903186, 0.002728201, 0.002776904, 0.002661174, 0.002548832, 
    0.002311479, 0.002062013, 0.002040541, 0.002001535, 0.001884533, 
    0.001867255, 0.001919629, 0.001992759, 0.002010767, 0.002075776, 
    0.002006078, 0.001942469, 0.001862139, 0.00178284, 0.001669751, 
    0.001611608, 0.001705498, 0.001347073, 0.001566895, 0.001461165, 
    0.001316874,
  0.001066423, 0.001799687, 0.001802422, 0.001240453, 0.001522676, 
    0.001175078, 0.0003555538, 0.0003768215, 0.0007686545, 0.0006798678, 
    0.0008860994, 0.0003488148, 0.0008009993, 0.001006597, 0.001718706, 
    0.001538079, 0.001591994, 0.001936523, 0.00212025, 0.002660602, 
    0.003124404, 0.002988205, 0.002344649, 0.002282517, 0.002434882, 
    0.00264358, 0.00240295, 0.002184084, 0.002120535, 0.002235056, 
    0.002239046, 0.002279768, 0.002530027, 0.00249608, 0.002467024, 
    0.002318152, 0.002257436, 0.002272854, 0.002268943, 0.002292785, 
    0.00237542, 0.002426744, 0.00243954, 0.002394001, 0.00228018, 
    0.002177659, 0.002082882, 0.001976276, 0.001870212, 0.001774527, 
    0.001757742, 0.001687138, 0.001589753, 0.001511742, 0.001473691, 
    0.001492097, 0.001409096, 0.00138066, 0.001360983, 0.00132363, 
    0.001270954, 0.001178115, 0.001213782, 0.001151189, 0.001202751, 
    0.001325061, 0.001354879, 0.0017562, 0.0018986, 0.002677338, 0.002840783, 
    0.00280793, 0.002811301, 0.002593891, 0.002604891, 0.002196211, 
    0.001946522, 0.001861565, 0.001907897, 0.001898664, 0.001824038, 
    0.001839806, 0.001892845, 0.001971445, 0.002067718, 0.002000787, 
    0.001972542, 0.001890828, 0.001746553, 0.001641459, 0.001522169, 
    0.001493925, 0.001654427, 0.001510882, 0.001457016, 0.0004888787,
  0.001205532, 0.001044886, 0.0004157473, 0.001344594, 0.001536775, 
    0.001474676, 0.001273498, 0.0008420558, 0.001738859, 0.001305272, 
    0.001100072, 0.0007575275, 0.001394073, 0.001668431, 0.0008231406, 
    0.0006007599, 0.0008996893, 0.0009580064, 0.0008768006, 0.002054891, 
    0.002243258, 0.001590992, 0.001330051, 0.0007900805, 0.0009166012, 
    0.001095638, 0.00124217, 0.001726715, 0.001853746, 0.002171971, 
    0.002336209, 0.002294566, 0.002168616, 0.001488741, 0.00195601, 
    0.00208881, 0.002041001, 0.00205734, 0.00209846, 0.002045165, 
    0.001997322, 0.002011182, 0.002030399, 0.002044625, 0.002028555, 
    0.002011913, 0.00196763, 0.001897472, 0.001799562, 0.00166673, 
    0.00158284, 0.001497103, 0.001448863, 0.001403722, 0.001368818, 
    0.001377862, 0.001283336, 0.001192897, 0.001141906, 0.001112979, 
    0.001156005, 0.001086483, 0.001062959, 0.001084846, 0.001157404, 
    0.001573699, 0.001598716, 0.001637865, 0.002016617, 0.002612123, 
    0.002708763, 0.002568842, 0.002562834, 0.002468199, 0.002461681, 
    0.00241689, 0.002278527, 0.002022911, 0.001935364, 0.001848532, 
    0.001717846, 0.001695371, 0.001661279, 0.001663201, 0.0017274, 
    0.001772652, 0.001802693, 0.001737556, 0.001710774, 0.001656399, 
    0.00155321, 0.001464264, 0.001469732, 0.001797081, 0.00206387, 0.001392357,
  0.001840251, 0.001856415, 0.001536506, 0.001610113, 0.001533104, 
    0.001476218, 0.001357405, 0.001361538, 0.001653982, 0.00167091, 
    0.001745917, 0.001331608, 0.001033522, 0.0008516726, 0.0005091755, 
    0.0006387322, 0.001171519, 0.0006707273, 0.0005509788, 0.001182628, 
    0.001340112, 0.001353082, 0.001271844, 0.0008513858, 0.001022491, 
    0.0007147719, 0.0008916627, 0.001320275, 0.001950828, 0.002287013, 
    0.002285918, 0.002138433, 0.002031478, 0.00140981, 0.001989962, 
    0.001959492, 0.002036119, 0.002163069, 0.002066161, 0.001975846, 
    0.00185473, 0.001748762, 0.001734663, 0.001757328, 0.001740958, 
    0.001732645, 0.001733868, 0.001720709, 0.001692194, 0.001642141, 
    0.001598764, 0.001488218, 0.001367483, 0.00130462, 0.001266488, 
    0.001290855, 0.001271256, 0.00114178, 0.0009934353, 0.0008960972, 
    0.0008989424, 0.0009178426, 0.0009628236, 0.001040198, 0.001417534, 
    0.001456269, 0.001547869, 0.001342226, 0.00179794, 0.002464845, 
    0.002579508, 0.002353312, 0.002369255, 0.002382019, 0.002345985, 
    0.002413917, 0.002332316, 0.002215824, 0.001967599, 0.001775211, 
    0.001695421, 0.001617679, 0.001461182, 0.00137303, 0.001302904, 
    0.001279857, 0.001368803, 0.001376828, 0.001415659, 0.001416693, 
    0.001410096, 0.001388145, 0.001340272, 0.001448291, 0.00154598, 
    0.001962131,
  0.001864649, 0.001421397, 0.00137535, 0.001368326, 0.001288137, 
    0.001234779, 0.001318178, 0.001311613, 0.001137313, 0.001269922, 
    0.001317955, 0.00130953, 0.001424099, 0.001491793, 0.001198461, 
    0.001056918, -4.298985e-006, -8.065673e-005, 0.00132018, 0.001530418, 
    0.001547202, 0.001337887, 0.0007693698, 0.001035174, 0.001552448, 
    0.00168798, 0.001176541, 0.001334819, 0.001818602, 0.001994269, 
    0.001962924, 0.002040251, 0.002018571, 0.001894944, 0.001878524, 
    0.001585618, 0.001613482, 0.001749906, 0.001644286, 0.001743548, 
    0.001688044, 0.001566769, 0.001566402, 0.00159239, 0.001557566, 
    0.001500488, 0.001464614, 0.001465583, 0.001435654, 0.001393962, 
    0.001362682, 0.001283686, 0.001210857, 0.001190178, 0.001169166, 
    0.001171471, 0.001145403, 0.00106992, 0.000963998, 0.000864164, 
    0.000817148, 0.0008631637, 0.0008932361, 0.0009977901, 0.0009898916, 
    0.0009947545, 0.000905348, 0.001159438, 0.001746312, 0.002145396, 
    0.002248408, 0.002177581, 0.002219432, 0.002306646, 0.00218049, 
    0.002216062, 0.002356553, 0.002181857, 0.001983539, 0.001726079, 
    0.001675201, 0.001539875, 0.001330829, 0.001052436, 0.0006315168, 
    0.0003388971, 0.0005448591, 0.0008497173, 0.001011238, 0.001068284, 
    0.001121785, 0.001220776, 0.001230837, 0.001242965, 0.001369628, 
    0.001606362,
  0.00118541, 0.001101328, 0.00112943, 0.001266171, 0.00123497, 0.001182294, 
    0.001186046, 0.001161329, 0.001215325, 0.001296785, 0.001357056, 
    0.001477743, 0.001423018, 0.001181483, 0.0009973142, 0.0007842947, 
    0.0006739385, 5.122134e-005, 0.0006405604, 0.00102036, 0.001366306, 
    0.001411081, 0.001505336, 0.001615882, 0.00150238, 0.001285991, 
    0.001237831, 0.001397428, 0.001434796, 0.00155267, 0.001549046, 
    0.001621128, 0.001598097, 0.001605679, 0.001546964, 0.001454442, 
    0.001208807, 0.001251038, 0.001381406, 0.001402149, 0.001336647, 
    0.001171248, 0.001071144, 0.001014797, 0.0009801956, 0.0009541917, 
    0.0009696414, 0.001009123, 0.001021315, 0.0010319, 0.001037908, 
    0.0010041, 0.0009695296, 0.0009520454, 0.0009226566, 0.000907477, 
    0.0008903751, 0.0008392585, 0.0008130162, 0.0007931795, 0.0007772218, 
    0.0008356026, 0.0008581574, 0.0007664771, 0.0008994192, 0.001005643, 
    0.001171931, 0.001472641, 0.001845766, 0.001977914, 0.001367482, 
    0.00180374, 0.002204061, 0.002108169, 0.001763622, 0.002113541, 
    0.002209798, 0.002137923, 0.001962543, 0.001838486, 0.001392262, 
    0.001177081, 0.00100987, 0.0007619313, 0.0005079671, 0.0004500644, 
    0.0004475843, 0.0005094297, 0.0005979938, 0.000767923, 0.0008939514, 
    0.0009904951, 0.00108103, 0.001128619, 0.001220219, 0.001315635,
  0.00101421, 0.0009014062, 0.001101709, 0.001242377, 0.001149567, 
    0.001145372, 0.001167862, 0.001250959, 0.001177113, 0.001190163, 
    0.001151142, 0.001264787, 0.001325281, 0.001144942, 0.001141144, 
    0.001278202, 0.001278536, 0.001137011, 0.001216182, 0.001459432, 
    0.001508944, 0.001456397, 0.001311438, 0.001224924, 0.001145308, 
    0.001045999, 0.0009582611, 0.001167465, 0.001290489, 0.001247399, 
    0.00125719, 0.00115858, 0.001215816, 0.001294828, 0.001345135, 
    0.001168626, 0.001022634, 0.001001399, 0.0009587379, 0.0007326689, 
    0.0007885862, 0.0007672557, 0.0007577669, 0.0007712133, 0.0007684319, 
    0.0007598167, 0.0007776036, 0.0008230619, 0.0008338061, 0.0008351412, 
    0.0008678208, 0.0008792649, 0.00085981, 0.0008485089, 0.0008161473, 
    0.0008006189, 0.0007799873, 0.0007686066, 0.0008076434, 0.0008733515, 
    0.000896113, 0.0008986243, 0.0008949689, 0.0008279732, 0.0008833022, 
    0.001022825, 0.00135046, 0.001690825, 0.001820811, 0.001817362, 
    0.001561777, 0.00208331, 0.002071342, 0.00150532, 0.001910854, 
    0.00211564, 0.002164357, 0.002067209, 0.001866286, 0.001679859, 
    0.001160042, 0.0008157184, 0.0006430401, 0.0005709734, 0.0005095252, 
    0.0005126405, 0.0004398595, 0.0003371807, 0.0002839179, 0.0004058303, 
    0.0006663576, 0.0008463785, 0.0009579421, 0.001034269, 0.001077438, 
    0.001138696,
  0.0008319155, 0.0007740902, 0.0008676932, 0.0009055063, 0.0008543734, 
    0.0008691717, 0.001015672, 0.001078074, 0.001077136, 0.00104681, 
    0.001163937, 0.001275517, 0.001339143, 0.001472784, 0.001351444, 
    0.00134728, 0.001384919, 0.001512123, 0.001503746, 0.00147129, 
    0.001546884, 0.001611797, 0.001350205, 0.001004053, 0.0008449801, 
    0.0008407841, 0.0008405615, 0.000836906, 0.0008672485, 0.0009326867, 
    0.000896574, 0.0008194377, 0.0008625914, 0.0009153299, 0.0008597779, 
    0.0007837065, 0.0007789861, 0.0006740026, 0.0004922643, 0.0006328516, 
    0.0008469515, 0.0008279572, 0.0008108071, 0.0008066581, 0.0008077393, 
    0.0007872353, 0.00079318, 0.0008024299, 0.0007862812, 0.0007768879, 
    0.0007978845, 0.0008138907, 0.00081904, 0.0008266699, 0.0008177529, 
    0.0007987428, 0.000786107, 0.0007966929, 0.0008120467, 0.000829387, 
    0.0008300073, 0.0008806475, 0.0009171576, 0.001066217, 0.001180864, 
    0.00106253, 0.001191069, 0.001279856, 0.001331847, 0.001314538, 
    0.001529528, 0.001588624, 0.0016265, 0.001665442, 0.001742547, 
    0.001703049, 0.001506893, 0.001365655, 0.001295465, 0.001150617, 
    0.0009221162, 0.000876944, 0.0005979792, 0.0006465362, 0.0005681915, 
    0.0004248866, 0.000211725, -4.905835e-005, -0.0001609721, -2.896693e-005, 
    0.0003029755, 0.0006050197, 0.000789572, 0.0008621146, 0.0008446937, 
    0.0008130637,
  0.0007851049, 0.0007302528, 0.0007688766, 0.0006331052, 0.0007286952, 
    0.0007065861, 0.0009272504, 0.001154145, 0.00130651, 0.001246651, 
    0.001278345, 0.001391228, 0.001410699, 0.001250817, 0.00115556, 
    0.001175937, 0.001118113, 0.001081619, 0.001107352, 0.001074212, 
    0.001090631, 0.001143496, 0.001111771, 0.0009132312, 0.0008014133, 
    0.0007396149, 0.0007294584, 0.0007029148, 0.0007496772, 0.0007765705, 
    0.0008200263, 0.0007901443, 0.0007420792, 0.000695667, 0.0006482855, 
    0.0006250157, 0.0005939261, 0.0006065306, 0.0004602843, 0.000547196, 
    0.0007913208, 0.0008355393, 0.0007827058, 0.00070735, 0.0007503759, 
    0.0007532998, 0.0007585296, 0.0007455917, 0.0007378189, 0.0007732003, 
    0.0008313581, 0.0008842717, 0.0009125955, 0.0009144871, 0.0009117532, 
    0.0008881502, 0.0008655, 0.0008699824, 0.0008854317, 0.0009108791, 
    0.0009044576, 0.001010475, 0.001200828, 0.001155592, 0.001071351, 
    0.0009886674, 0.001058365, 0.001118017, 0.00116292, 0.001212081, 
    0.00124031, 0.001283289, 0.001315619, 0.001218121, 0.001116046, 
    0.0008350941, 0.0009761741, 0.0009390446, 0.0008410546, 0.000693108, 
    0.0005888394, 0.000263589, 0.0003519948, 0.0003971506, 0.0003302186, 
    0.0003294074, 0.0001784894, -7.232744e-005, -0.0002426533, -0.0001478107, 
    0.0001640883, 0.0004654969, 0.0006516222, 0.0007252144, 0.0008107433, 
    0.0008579185,
  0.000583387, 0.0006436277, 0.0006662775, 0.0008416586, 0.0008249213, 
    0.0008887695, 0.0008160044, 0.00114774, 0.001303555, 0.001369359, 
    0.001271002, 0.001194502, 0.001183185, 0.001168625, 0.00107302, 
    0.0009811651, 0.0009054905, 0.0008873711, 0.0008681705, 0.0008473322, 
    0.0008545639, 0.0008436292, 0.000835666, 0.0008055773, 0.0007839766, 
    0.0007343544, 0.0006318346, 0.0006069911, 0.0006099159, 0.0006073408, 
    0.0005513283, 0.0006104244, 0.0006319298, 0.0005780628, 0.0005072844, 
    0.0004719666, 0.0004937104, 0.0005244506, 0.0004276524, 0.0003556823, 
    0.0003805729, 0.0003971667, 0.0005162647, 0.0005732786, 0.0005443506, 
    0.0006521798, 0.0007274086, 0.0008038932, 0.0009129292, 0.001003656, 
    0.001078042, 0.001023619, 0.0009117057, 0.0009203679, 0.0008148602, 
    0.0008435654, 0.0008327095, 0.0008300235, 0.0008323281, 0.0008538649, 
    0.001051912, 0.001203562, 0.000819549, 0.0008102187, 0.0008736541, 
    0.001007692, 0.001046444, 0.0009919098, 0.0009846459, 0.001009521, 
    0.0009915286, 0.0009398714, 0.0007260416, 0.0006323906, 0.0005646637, 
    0.0005747885, 0.0008597467, 0.0008999279, 0.0008056255, 0.0005731513, 
    0.000335607, 0.0002316725, 0.0001214433, -3.75493e-005, -4.171464e-005, 
    0.0001955279, 0.0003067581, 0.0002394128, 0.0001558871, 0.0001815567, 
    0.0002899258, 0.0004127906, 0.0005080309, 0.0005645519, 0.0005871695, 
    0.0006949827,
  0.0003731181, 0.0003989153, 0.0006420068, 0.0007581483, 0.0006823312, 
    0.0005037235, 0.0006932663, 0.0007846286, 0.0009190482, 0.001003386, 
    0.001018406, 0.0009465623, 0.0008601276, 0.0007726913, 0.0007375486, 
    0.0007441607, 0.0007876332, 0.0008147333, 0.0008090271, 0.0008224584, 
    0.0008174037, 0.0007693225, 0.0007317953, 0.0006898653, 0.0006014123, 
    0.0005775066, 0.0005169641, 0.0005140079, 0.0004844917, 0.0004399233, 
    0.0004082455, 0.000436649, 0.0005110358, 0.0004953002, 0.0004058296, 
    0.0003466383, 0.0003667763, 0.0004127752, 0.000349785, 0.0002515407, 
    0.000213457, 0.0002959976, 0.0003065199, 0.0002701371, 0.0002988905, 
    0.000359115, 0.0004311176, 0.0004853338, 0.000550756, 0.0005890145, 
    0.0006139213, 0.0005423161, 0.0007060138, 0.0007290924, 0.0007822914, 
    0.0008626706, 0.0008198349, 0.0006614146, 0.0006007927, 0.0006079925, 
    0.0006480785, 0.0006711415, 0.00073259, 0.0008016517, 0.0009353249, 
    0.001043408, 0.001044092, 0.0009999205, 0.0009518713, 0.0009156002, 
    0.0008593174, 0.0006273203, 0.000565045, 0.0005189988, 0.0005123706, 
    0.0005457015, 0.000679597, 0.0006189118, 0.0004807087, 0.0003984862, 
    0.0002957119, 0.000189536, 7.705018e-005, -7.794937e-006, 2.782466e-005, 
    4.093791e-005, 0.0001161979, 0.0002362975, 0.0003295671, 0.0003983746, 
    0.0004357109, 0.0003529796, 0.0001964658, 0.0002205302, 0.0003383248, 
    0.0003782995,
  0.00027578, 0.0003345897, 0.0003590672, 0.0006013, 0.0006465525, 
    0.0006769905, 0.0004623979, 0.0007299194, 0.0007683372, 0.0008162751, 
    0.0008412136, 0.0008325032, 0.0007816406, 0.0007553191, 0.0007728192, 
    0.0008039249, 0.0008616061, 0.0008551213, 0.0008447419, 0.0008057842, 
    0.0008097105, 0.0007733915, 0.0006893086, 0.0006165437, 0.0005575749, 
    0.0005203022, 0.0004986539, 0.0005038669, 0.0004654818, 0.0003891084, 
    0.0003890924, 0.0003669355, 0.0003481165, 0.0003524716, 0.000302165, 
    0.0002863817, 0.0003693989, 0.0003157863, 0.0002786089, 0.0002360274, 
    0.0001992474, 0.0002689133, 0.0002709636, 0.0002512704, 0.0002382365, 
    0.0002451031, 0.0002390633, 0.0002411294, 0.0002361548, 0.0002352169, 
    0.0003287566, 0.0002858571, 0.0005119089, 0.0005653948, 0.0006339797, 
    0.0006038593, 0.0005409492, 0.0005296324, 0.0005650457, 0.0006496205, 
    0.0007193971, 0.000786647, 0.0007880302, 0.0008741152, 0.0008867194, 
    0.0008981794, 0.0009203688, 0.0009117064, 0.000890153, 0.0008627188, 
    0.0007916063, 0.0006637659, 0.0005702744, 0.0005194752, 0.0004876386, 
    0.0004730152, 0.0004520188, 0.0004741279, 0.0004176865, 0.0003772189, 
    0.0003296146, 0.0002461048, 0.000233691, 0.0002214839, 0.0002065748, 
    0.0001865316, 0.0001710504, 0.0001249406, 0.0002230264, 0.0004170195, 
    0.0005045983, 0.0005043754, 0.0003481316, 0.0001003514, 4.057167e-005, 
    0.0001167068,
  0.0003079348, 0.0002934546, 0.0002991608, 0.000224933, 0.0001312979, 
    0.0005597046, 0.000613699, 0.0006236646, 0.0006240774, 0.0005878857, 
    0.0005962939, 0.0004555478, 0.0004162404, 0.0003970398, 0.0005385808, 
    0.0005735967, 0.000623839, 0.0006586958, 0.0006598083, 0.000633376, 
    0.000605274, 0.000562025, 0.0005150882, 0.0004710283, 0.0004302589, 
    0.0004143009, 0.000390904, 0.0003884882, 0.0003988352, 0.0004149207, 
    0.000436506, 0.0004018876, 0.0003611499, 0.0003039925, 0.0003271033, 
    0.0002991764, 0.0002432596, 0.0002382686, 0.0001460959, 0.0001559663, 
    0.0001175811, 0.0001407396, 0.0001439024, 0.0001386416, 0.0001860708, 
    0.0001794428, 0.0001994064, 0.0002175421, 0.0002254415, 0.0002128691, 
    0.0002623489, 0.0003307434, 0.0003970873, 0.0005194596, 0.0005764889, 
    0.0006288141, 0.0006759737, 0.0007791291, 0.0009365329, 0.0009255181, 
    0.0009683857, 0.001029675, 0.001080395, 0.001073878, 0.00108475, 
    0.0009922914, 0.0009178729, 0.0008336636, 0.0007769354, 0.0005829742, 
    0.0006298791, 0.0006116639, 0.0005628516, 0.0004916121, 0.0005529651, 
    0.0004844436, 0.0004901498, 0.0004699635, 0.0004577725, 0.0004205792, 
    0.0003629613, 0.0003027208, 0.0003252118, 0.0002914199, 0.0002725529, 
    0.0002483772, 0.0002513974, 0.0002764629, 0.0003464946, 0.0004213739, 
    0.0004465349, 0.0004485224, 0.0004273029, 0.0003653299, 0.0003724191, 
    0.000332746,
  0.0005244822, 0.0004638769, 0.0003963241, 0.0003697169, 0.0003405185, 
    0.0004168288, 0.0005466875, 0.0006255081, 0.0006245065, 0.0006327562, 
    0.0006315003, 0.0006411008, 0.0006064028, 0.0005744386, 0.0005373408, 
    0.0005653627, 0.0005373727, 0.0005363394, 0.0005305858, 0.0005785873, 
    0.000592495, 0.0005929084, 0.0005792866, 0.0005475134, 0.0005154859, 
    0.0005064895, 0.0004971753, 0.0004701067, 0.0004658469, 0.0004288764, 
    0.0004270959, 0.0004223436, 0.0004005681, 0.000356731, 0.0002905617, 
    0.0002878753, 0.0003057248, 0.0003137041, 0.0003330638, 0.0003063928, 
    0.0002555619, 0.0002271582, 0.0002104056, 0.0001984686, 0.0001857688, 
    0.0001700172, 0.0001570155, 0.0001583028, 0.0001732914, 0.0002076236, 
    0.000255657, 0.0003098577, 0.0003581771, 0.0003975956, 0.0004265078, 
    0.0004459627, 0.0004685014, 0.0004965393, 0.0005326201, 0.0005638371, 
    0.0005901742, 0.0006054016, 0.000587997, 0.0007528078, 0.0007066182, 
    0.000721893, 0.0007045039, 0.0006014436, 0.0005577337, 0.0004403681, 
    0.0004739532, 0.0004809787, 0.0004673412, 0.0004917231, 0.0004965867, 
    0.0004921841, 0.00047861, 0.0004715212, 0.0004601886, 0.0004441192, 
    0.0004122664, 0.000466419, 0.0003425367, 0.0003118921, 0.0002811041, 
    0.000264399, 0.0002524462, 0.0002602029, 0.0002896239, 0.0003468759, 
    0.0004394779, 0.0004930586, 0.0005568436, 0.0005631379, 0.0005136898, 
    0.0004971912,
  0.000555747, 0.0005426817, 0.0005278043, 0.0005561921, 0.0005741846, 
    0.000552743, 0.0005773157, 0.0005535532, 0.0005298069, 0.0004933447, 
    0.0004830926, 0.0004752405, 0.0004693597, 0.0004536875, 0.0004379519, 
    0.0004299571, 0.0004254429, 0.0004257134, 0.0004339467, 0.0004492373, 
    0.0004672775, 0.0004799931, 0.000480915, 0.0004637807, 0.0004355998, 
    0.0005020865, 0.0004834264, 0.0004501113, 0.0004422276, 0.0004268894, 
    0.0004036516, 0.000376901, 0.0003617057, 0.0003502934, 0.0003402799, 
    0.0003333814, 0.0003258474, 0.0003107633, 0.0002918011, 0.0002637631, 
    0.0002376165, 0.0002163654, 0.0002025849, 0.0001966722, 0.0001961157, 
    0.0002016471, 0.0002131548, 0.00023288, 0.0002611405, 0.0002965697, 
    0.0003370532, 0.0003771551, 0.0004137604, 0.0004430859, 0.0004619686, 
    0.000477418, 0.0004949495, 0.0005153423, 0.0005401064, 0.0005721658, 
    0.0006040661, 0.0006352355, 0.0006572177, 0.0006649424, 0.000653244, 
    0.0006070859, 0.0005746293, 0.0005494048, 0.0005255945, 0.000528074, 
    0.0005141025, 0.0005113529, 0.0005009102, 0.0005099382, 0.0005070136, 
    0.0004644161, 0.0004479971, 0.0004499363, 0.0004337396, 0.0004225499, 
    0.0004040328, 0.0003712901, 0.0003336676, 0.0002978888, 0.0002726801, 
    0.0002604412, 0.0002624281, 0.0002830751, 0.0003304887, 0.0003964195, 
    0.0004749702, 0.0005744386, 0.0006158758, 0.0006404012, 0.000651448, 
    0.0006351401,
  0.0005564141, 0.0005664756, 0.0005826245, 0.0005966752, 0.0005825926, 
    0.000587504, 0.0005858032, 0.0005984235, 0.000580129, 0.0005611983, 
    0.0005437462, 0.0005263735, 0.0005108443, 0.0004986372, 0.0004899269, 
    0.0004850155, 0.0004859533, 0.0004910557, 0.0005020866, 0.0005158989, 
    0.0005262144, 0.0005332876, 0.0005360692, 0.0005279946, 0.0005059649, 
    0.0004878768, 0.0004714259, 0.0004597276, 0.0004393348, 0.0004187037, 
    0.0003933995, 0.0003688264, 0.0003502457, 0.000334939, 0.0003181384, 
    0.000305407, 0.000292421, 0.0002827729, 0.000271774, 0.0002640014, 
    0.0002576755, 0.0002551483, 0.0002555614, 0.0002547668, 0.0002537973, 
    0.0002533363, 0.0002522077, 0.000253988, 0.0002545284, 0.0002563245, 
    0.0002626982, 0.0002725051, 0.0002827571, 0.0002940899, 0.0003090785, 
    0.0003268329, 0.0003458268, 0.0003665534, 0.0003852614, 0.0004044462, 
    0.0004179565, 0.0004287171, 0.0004340417, 0.0004328338, 0.0004324365, 
    0.0004278587, 0.0004267143, 0.0004281924, 0.0004334694, 0.0004407491, 
    0.0004511283, 0.0004778472, 0.0004483152, 0.0004195777, 0.0004060675, 
    0.0003890443, 0.0003676342, 0.0003467488, 0.0003289151, 0.000312941, 
    0.0002990651, 0.0002873507, 0.0002792445, 0.0002753185, 0.0002767014, 
    0.0002827572, 0.0002966332, 0.0003170578, 0.0003466852, 0.0003814466, 
    0.000419848, 0.0004545138, 0.0005068867, 0.0005172977, 0.0005278517, 
    0.0005410918,
  0.0004451044, 0.0004364101, 0.0004310855, 0.0004239646, 0.0004123456, 
    0.0004010764, 0.0003899025, 0.000376853, 0.0003653773, 0.0003539807, 
    0.0003424729, 0.0003335879, 0.0003270075, 0.0003238287, 0.0003268328, 
    0.0003320302, 0.000338547, 0.0003494667, 0.0003609108, 0.0003737694, 
    0.0003889805, 0.0004023003, 0.0004102157, 0.0004162715, 0.0004183378, 
    0.0004131561, 0.0004081811, 0.0003987239, 0.000383783, 0.0003707972, 
    0.0003525502, 0.0003334131, 0.0003169782, 0.0003011631, 0.0002872553, 
    0.0002763198, 0.0002705024, 0.0002692945, 0.000268452, 0.0002697076, 
    0.0002732998, 0.0002778934, 0.0002828684, 0.0002884791, 0.0002959337, 
    0.0003024028, 0.000307505, 0.0003140853, 0.0003199665, 0.0003256249, 
    0.0003342079, 0.0003446665, 0.0003573028, 0.0003716715, 0.000387423, 
    0.0004028726, 0.0004198798, 0.0004343755, 0.0004469958, 0.0004584877, 
    0.000467309, 0.000474525, 0.0004784988, 0.0004797544, 0.0004765437, 
    0.0004721569, 0.0004667686, 0.0004611737, 0.0004561828, 0.000451033, 
    0.000446932, 0.0004415439, 0.0004387306, 0.0004347886, 0.000431117, 
    0.0004300204, 0.0004302429, 0.0004248548, 0.0004229156, 0.0004251725, 
    0.0004230109, 0.0004285423, 0.0004348205, 0.000440177, 0.0004488078, 
    0.0004561511, 0.0004633514, 0.0004654018, 0.0004668798, 0.0004706945, 
    0.000471076, 0.0004730627, 0.0004702178, 0.0004605857, 0.0004556425, 
    0.0004512396,
  0.0004557854, 0.0004578676, 0.0004589008, 0.0004571524, 0.0004572001, 
    0.0004573591, 0.0004570889, 0.0004566121, 0.0004564848, 0.0004569618, 
    0.0004570095, 0.0004578518, 0.0004600135, 0.0004608083, 0.0004607287, 
    0.0004604108, 0.0004611579, 0.0004606175, 0.000460236, 0.0004597751, 
    0.0004586625, 0.0004566757, 0.0004535444, 0.000447568, 0.000442768, 
    0.0004364578, 0.0004303383, 0.0004221845, 0.0004145869, 0.0004051137, 
    0.0003961014, 0.0003867553, 0.0003772663, 0.0003657109, 0.0003549822, 
    0.0003454455, 0.0003333815, 0.0003237812, 0.0003155159, 0.0003064243, 
    0.0002989061, 0.000292755, 0.0002877958, 0.0002839334, 0.0002805956, 
    0.0002773054, 0.0002754775, 0.0002744603, 0.0002741741, 0.0002743966, 
    0.0002767968, 0.0002778617, 0.000282026, 0.0002855387, 0.0002896396, 
    0.0002932476, 0.0002963153, 0.0002987153, 0.0003025301, 0.0003038335, 
    0.0003053594, 0.0003072984, 0.0003074416, 0.0003074574, 0.0003082837, 
    0.0003087923, 0.0003086494, 0.0003082997, 0.0003084586, 0.0003092374, 
    0.0003109063, 0.0003129409, 0.0003142761, 0.0003157702, 0.0003172484, 
    0.0003210789, 0.0003241625, 0.0003281202, 0.0003343191, 0.0003401842, 
    0.0003477978, 0.0003556972, 0.000364789, 0.000374135, 0.0003842122, 
    0.0003935104, 0.0004015532, 0.0004092144, 0.0004176543, 0.0004271592, 
    0.0004344867, 0.0004404471, 0.0004441505, 0.0004477905, 0.0004510011, 
    0.0004534648,
  1.456728e-005, 1.396328e-005, 1.339108e-005, 1.285067e-005, 1.229435e-005, 
    1.173804e-005, 1.126121e-005, 1.059363e-005, 1.002143e-005, 
    9.544594e-006, 9.099545e-006, 8.686286e-006, 8.257134e-006, 7.85977e-006, 
    7.525985e-006, 7.271672e-006, 6.969673e-006, 6.810728e-006, 
    6.715361e-006, 6.588203e-006, 6.508732e-006, 6.445153e-006, 
    6.461047e-006, 6.57231e-006, 6.683572e-006, 6.810726e-006, 7.033253e-006, 
    7.176303e-006, 7.525984e-006, 7.764402e-006, 8.193556e-006, 
    8.543235e-006, 9.020072e-006, 9.512805e-006, 9.926063e-006, 
    1.053005e-005, 1.105458e-005, 1.165857e-005, 1.250098e-005, 
    1.308908e-005, 1.385202e-005, 1.464675e-005, 1.53938e-005, 1.615674e-005, 
    1.696736e-005, 1.780978e-005, 1.86204e-005, 1.922439e-005, 1.976481e-005, 
    2.025755e-005, 2.073438e-005, 2.095691e-005, 2.102049e-005, 
    2.111585e-005, 2.090922e-005, 2.082975e-005, 2.040059e-005, 
    2.017807e-005, 1.970123e-005, 1.928797e-005, 1.897008e-005, 
    1.846145e-005, 1.828662e-005, 1.788925e-005, 1.760315e-005, 
    1.739652e-005, 1.738063e-005, 1.723757e-005, 1.731705e-005, 
    1.750778e-005, 1.766673e-005, 1.787336e-005, 1.817535e-005, 
    1.822304e-005, 1.869988e-005, 1.898598e-005, 1.927208e-005, 
    1.954229e-005, 2.000323e-005, 2.017806e-005, 2.025754e-005, 2.03688e-005, 
    2.032112e-005, 2.027344e-005, 1.998734e-005, 1.971712e-005, 
    1.941513e-005, 1.903366e-005, 1.855682e-005, 1.812767e-005, 
    1.769851e-005, 1.717399e-005, 1.674484e-005, 1.615674e-005, 
    1.563221e-005, 1.506001e-005,
  2.159268e-005, 2.044827e-005, 1.914492e-005, 1.784156e-005, 1.647463e-005, 
    1.504412e-005, 1.36295e-005, 1.231025e-005, 1.087974e-005, 9.544595e-006, 
    8.304817e-006, 7.128619e-006, 6.000104e-006, 5.078219e-006, 
    4.251703e-006, 3.679499e-006, 3.218556e-006, 2.916559e-006, 2.70993e-006, 
    2.614562e-006, 2.694035e-006, 2.694035e-006, 2.85298e-006, 3.107294e-006, 
    3.298029e-006, 3.647709e-006, 4.029179e-006, 4.649066e-006, 
    5.157692e-006, 5.809369e-006, 6.651782e-006, 7.398826e-006, 8.24124e-006, 
    9.35386e-006, 1.046648e-005, 1.199236e-005, 1.36295e-005, 1.575937e-005, 
    1.823893e-005, 2.103638e-005, 2.418352e-005, 2.782337e-005, 
    3.141552e-005, 3.543686e-005, 3.920386e-005, 4.219206e-005, 
    4.632465e-005, 4.990092e-005, 5.350897e-005, 5.702167e-005, 6.04867e-005, 
    6.460338e-005, 6.721009e-005, 7.043668e-005, 6.89903e-005, 7.404476e-005, 
    7.325003e-005, 7.127909e-005, 6.870418e-005, 6.474643e-005, 
    6.034362e-005, 5.554347e-005, 5.029827e-005, 4.545042e-005, 
    4.131783e-005, 3.812303e-005, 3.585011e-005, 3.41176e-005, 3.289372e-005, 
    3.217848e-005, 3.219437e-005, 3.225795e-005, 3.267121e-005, 
    3.324342e-005, 3.419709e-005, 3.557992e-005, 3.694685e-005, 
    3.864757e-005, 3.99986e-005, 4.106353e-005, 4.316161e-005, 4.370203e-005, 
    4.43537e-005, 4.37974e-005, 4.394046e-005, 4.227153e-005, 4.082513e-005, 
    3.858397e-005, 3.594548e-005, 3.32434e-005, 3.057313e-005, 2.815716e-005, 
    2.632927e-005, 2.486697e-005, 2.369077e-005, 2.256225e-005,
  2.173573e-005, 1.750777e-005, 1.412223e-005, 1.15791e-005, 9.751222e-006, 
    8.193555e-006, 7.112722e-006, 6.270313e-006, 5.841158e-006, 
    5.507373e-006, 5.396112e-006, 5.412006e-006, 5.60274e-006, 5.84116e-006, 
    6.33389e-006, 6.890201e-006, 7.557775e-006, 7.859773e-006, 8.034613e-006, 
    7.764404e-006, 7.287565e-006, 6.476942e-006, 5.332533e-006, 
    4.188125e-006, 3.345712e-006, 3.011925e-006, 2.964242e-006, 
    3.329817e-006, 3.886128e-006, 4.569594e-006, 5.28485e-006, 5.920633e-006, 
    6.508732e-006, 6.906096e-006, 7.255776e-006, 7.986928e-006, 9.33796e-006, 
    1.164267e-005, 1.506001e-005, 1.976481e-005, 2.51054e-005, 3.022345e-005, 
    3.507128e-005, 3.790051e-005, 3.799587e-005, 3.882239e-005, 
    3.842503e-005, 3.797998e-005, 3.874292e-005, 4.114301e-005, 
    4.498949e-005, 5.034598e-005, 5.783229e-005, 6.624052e-005, 
    7.480769e-005, 8.089533e-005, 8.46464e-005, 8.536165e-005, 8.43921e-005, 
    8.191257e-005, 7.81773e-005, 7.375859e-005, 6.867237e-005, 6.390402e-005, 
    6.051848e-005, 5.899261e-005, 5.923102e-005, 5.983502e-005, 
    5.937406e-005, 5.760977e-005, 5.465337e-005, 5.10294e-005, 4.692863e-005, 
    4.390866e-005, 4.184235e-005, 4.107942e-005, 4.034829e-005, 
    4.333645e-005, 4.778695e-005, 5.354077e-005, 6.039132e-005, 
    6.728955e-005, 7.310697e-005, 7.886082e-005, 8.364508e-005, 
    8.679221e-005, 8.714189e-005, 8.698294e-005, 8.320002e-005, 
    7.661968e-005, 6.872007e-005, 5.932639e-005, 4.980555e-005, 
    4.141322e-005, 3.372025e-005, 2.721937e-005,
  2.259404e-005, 1.89065e-005, 1.677662e-005, 1.540969e-005, 1.423349e-005, 
    1.334339e-005, 1.288245e-005, 1.232614e-005, 1.15791e-005, 1.048237e-005, 
    8.988285e-006, 7.287563e-006, 5.714001e-006, 4.903377e-006, 
    4.537805e-006, 4.474226e-006, 4.521913e-006, 4.887486e-006, 
    5.602735e-006, 7.223989e-006, 8.972394e-006, 9.798907e-006, 
    9.449228e-006, 8.431971e-006, 7.176304e-006, 6.524625e-006, 
    6.222629e-006, 6.413365e-006, 7.065043e-006, 8.129977e-006, 
    9.226703e-006, 1.04029e-005, 1.12771e-005, 1.178573e-005, 1.232614e-005, 
    1.348645e-005, 1.47898e-005, 1.634747e-005, 1.850913e-005, 2.179932e-005, 
    2.621801e-005, 3.135196e-005, 3.721706e-005, 4.174699e-005, 
    4.494181e-005, 4.864525e-005, 6.991217e-005, 6.60021e-005, 7.250298e-005, 
    8.207151e-005, 9.216458e-005, 0.0001030682, 0.0001149732, 0.0001248597, 
    0.0001322189, 0.0001359064, 0.0001423118, 0.0001166263, 0.0001143374, 
    0.0001148143, 0.0001148779, 0.0001140673, 0.0001067875, 9.550242e-005, 
    8.324769e-005, 7.220102e-005, 6.57319e-005, 6.358614e-005, 6.325237e-005, 
    6.391991e-005, 6.473053e-005, 6.498485e-005, 6.323644e-005, 
    6.233048e-005, 6.349078e-005, 6.733726e-005, 7.229636e-005, 
    7.970323e-005, 8.696706e-005, 9.465999e-005, 0.0001240331, 0.0001231113, 
    0.0001236994, 0.000125114, 0.0001272756, 0.0001314241, 0.0001360971, 
    0.0001422006, 0.0001533746, 0.00011003, 9.470768e-005, 7.86224e-005, 
    6.272782e-005, 4.872471e-005, 3.726473e-005, 2.858631e-005,
  6.407886e-005, 5.632233e-005, 4.932872e-005, 4.335236e-005, 3.804357e-005, 
    3.38633e-005, 3.157449e-005, 3.155859e-005, 3.257584e-005, 3.254406e-005, 
    2.904725e-005, 2.284836e-005, 1.604547e-005, 1.094331e-005, 
    8.384292e-006, 8.38429e-006, 9.973746e-006, 1.297782e-005, 1.726936e-005, 
    1.995555e-005, 2.33411e-005, 2.639286e-005, 2.639286e-005, 2.251457e-005, 
    1.792104e-005, 1.442423e-005, 1.294603e-005, 1.345466e-005, 
    1.523485e-005, 1.776208e-005, 1.881113e-005, 1.873166e-005, 
    1.874755e-005, 2.025754e-005, 2.404045e-005, 2.876114e-005, 
    3.186058e-005, 3.297321e-005, 3.316395e-005, 3.405404e-005, 3.76621e-005, 
    4.241459e-005, 4.786641e-005, 5.11248e-005, 5.190363e-005, 5.431961e-005, 
    7.189899e-005, 8.569549e-005, 0.0001020828, 0.0001182793, 0.0001290558, 
    0.0001358746, 0.0001411356, 0.000143345, 0.0001401502, 0.00013295, 
    0.0001283088, 0.0001275618, 0.0001335857, 0.0001515148, 0.0001744825, 
    0.0001935401, 0.0002040782, 0.0002036967, 0.0001963375, 0.0001929202, 
    0.0001957336, 0.0002083062, 0.0002344529, 0.0002533357, 0.0002393006, 
    0.0002672274, 0.0002677678, 0.0002681334, 0.0002701997, 0.0002702633, 
    0.0002431312, 0.0002362806, 0.0002286989, 0.0002248206, 0.000252509, 
    0.000244816, 0.0002432425, 0.0002440372, 0.0002495526, 0.0002583105, 
    0.0002628723, 0.0002566734, 0.0002383787, 0.0002094347, 0.0001901863, 
    0.0001164515, 9.733028e-005, 8.593389e-005, 7.663557e-005, 7.073869e-005,
  0.0003135124, 0.0002923249, 0.0001597483, 0.000124367, 9.704422e-005, 
    8.378812e-005, 8.286623e-005, 9.458055e-005, 0.0001171031, 0.0001411039, 
    0.0001508473, 0.0001404046, 0.0001087267, 7.010291e-005, 4.17788e-005, 
    2.755316e-005, 2.318215e-005, 2.361131e-005, 2.844323e-005, 
    3.057311e-005, 3.421295e-005, 3.863167e-005, 4.104762e-005, 
    4.168339e-005, 4.08887e-005, 4.065027e-005, 4.386096e-005, 5.236456e-005, 
    6.320466e-005, 7.126322e-005, 6.964196e-005, 6.166287e-005, 
    5.562295e-005, 5.449443e-005, 5.966017e-005, 6.728955e-005, 
    7.334541e-005, 7.350433e-005, 6.846576e-005, 6.71942e-005, 7.142215e-005, 
    7.890849e-005, 8.711009e-005, 9.027313e-005, 0.0001041967, 0.0001048166, 
    0.0001137334, 0.0001257974, 0.0001263061, 0.00011065, 9.240309e-005, 
    7.398124e-005, 6.46034e-005, 6.881554e-005, 7.301173e-005, 8.084788e-005, 
    9.844324e-005, 0.0001300097, 0.0001680455, 0.0002031565, 0.0002290647, 
    0.0002510787, 0.0002845845, 0.0003249567, 0.000365313, 0.0003992162, 
    0.0004239642, 0.0004476788, 0.0004782282, 0.0005053761, 0.0005259755, 
    0.0005056465, 0.0005086982, 0.0005190773, 0.0005337162, 0.0005316976, 
    0.0005142293, 0.000491993, 0.0004500629, 0.0004408438, 0.0004939954, 
    0.0004856348, 0.0004727124, 0.0004501104, 0.0004310051, 0.0004244566, 
    0.0004308144, 0.0004296541, 0.0004137913, 0.0003817159, 0.0003530103, 
    0.00033284, 0.0003230649, 0.0003235736, 0.0003257353, 0.0003198384,
  0.001021504, 0.001027878, 0.0009769204, 0.0008718253, 0.0007889032, 
    0.0007396619, 0.0007030407, 0.0006731748, 0.0006594897, 0.0006759246, 
    0.000709335, 0.0006988128, 0.0006075937, 0.0004565952, 0.0003262438, 
    0.000230193, 0.0001806655, 0.0001617033, 0.0001623708, 0.0001704453, 
    0.000179696, 0.0001812218, 0.0001822868, 0.000176819, 0.0001755951, 
    0.0001799025, 0.0001857834, 0.0001894393, 0.0001950024, 0.0002025047, 
    0.0002131383, 0.000210341, 0.0002057632, 0.0001807291, 0.0001833199, 
    0.0001946845, 0.0002313058, 0.0002426228, 0.0002262197, 0.0001990241, 
    0.0001791081, 0.0001626095, 0.0001499894, 0.0001384817, 0.0001300577, 
    0.0001227303, 9.07029e-005, 2.447015e-005, -6.577931e-005, -0.0001284196, 
    -0.000149782, -0.0001375591, -0.0001077091, -6.770249e-005, 
    -5.870615e-005, -3.826548e-005, 3.871182e-005, 0.0001292313, 
    0.0002015675, 0.0002619349, 0.0002871596, 0.0003392301, 0.0004167161, 
    0.0005065047, 0.0005647263, 0.0005939247, 0.0006084363, 0.000625809, 
    0.0006462175, 0.0006673571, 0.0007063784, 0.0007682561, 0.0008152567, 
    0.0008575839, 0.0008848433, 0.000897988, 0.0008937283, 0.0008757039, 
    0.0009008489, 0.0008932829, 0.0007790647, 0.0007469259, 0.0007119102, 
    0.0006718242, 0.0006412904, 0.0006370309, 0.0006416243, 0.0006421489, 
    0.0006339473, 0.0006264452, 0.0006270967, 0.0006408137, 0.0006744306, 
    0.0007403932, 0.0008316122, 0.000937486,
  0.001257841, 0.001279744, 0.001280808, 0.001263483, 0.001245729, 
    0.001225575, 0.001190067, 0.00115459, 0.001125153, 0.001103235, 
    0.001082603, 0.001082937, 0.001104713, 0.00114313, 0.001174426, 
    0.001206088, 0.001210268, 0.001198093, 0.001143559, 0.001016434, 
    0.0009041394, 0.0008341394, 0.0007876637, 0.0007715625, 0.0007579568, 
    0.0006853028, 0.0006036683, 0.000534956, 0.0004963002, 0.0004672292, 
    0.0004136167, 0.0003472567, 0.0002971089, 0.0002642549, 0.0002670048, 
    0.0002888916, 0.0003560937, 0.0003778217, 0.0003597494, 0.0003470974, 
    0.0003756282, 0.0003964026, 0.0003763593, 0.0003385143, 0.0003007015, 
    0.0002224206, 8.976436e-005, -6.358651e-005, -0.0001288657, 
    -0.0001410886, -0.0001518175, -0.0001706521, -0.0001810312, -0.00014565, 
    -9.717164e-005, -7.102499e-005, -6.397488e-006, 6.830692e-005, 
    0.0001249553, 0.0001604001, 0.0001777411, 0.0002013126, 0.000234246, 
    0.0002837419, 0.0003312666, 0.0003879941, 0.0004576442, 0.000522081, 
    0.0005741674, 0.0006072437, 0.0006222005, 0.0006362514, 0.0006789286, 
    0.0007177591, 0.0007323499, 0.0007200001, 0.0006949182, 0.0006779749, 
    0.0006620327, 0.0006530045, 0.0007402818, 0.000790159, 0.0007858677, 
    0.0007936083, 0.0008361578, 0.0008768798, 0.0009195727, 0.0009263436, 
    0.0009257556, 0.0009522835, 0.0009819428, 0.0009939432, 0.000993371, 
    0.001022665, 0.001093777, 0.001183247,
  0.0008501294, 0.0008350774, 0.0007966124, 0.0007666349, 0.0007539191, 
    0.0007196821, 0.0006748913, 0.0006262539, 0.0006054163, 0.0006086431, 
    0.0006154617, 0.000623568, 0.00063959, 0.0006630979, 0.0006856525, 
    0.0007125137, 0.0007419663, 0.0007792232, 0.0008042254, 0.0007863122, 
    0.0007453202, 0.000685811, 0.0006242674, 0.000580128, 0.0005464947, 
    0.0005110819, 0.0004748581, 0.0004423214, 0.0004104851, 0.0003894565, 
    0.0003804283, 0.0003629443, 0.0003213165, 0.0002868411, 0.0002651291, 
    0.0002558148, 0.0002780354, 0.0003270062, 0.0003537731, 0.0003604961, 
    0.000390267, 0.0004493468, 0.0005090311, 0.0005407408, 0.0005419804, 
    0.0005086176, 0.0004002643, 0.0002541775, 0.0001281016, 5.106069e-005, 
    1.467858e-005, -1.458405e-005, -5.384348e-005, -7.069157e-005, 
    -6.806874e-005, -8.53464e-005, -8.05303e-005, -1.291488e-005, 
    6.825873e-005, 0.0001131608, 0.0001476044, 0.0002004222, 0.0002418594, 
    0.0002698814, 0.0003120336, 0.000388328, 0.0004749694, 0.0005278182, 
    0.0005487837, 0.0005700025, 0.0005938765, 0.0006194026, 0.0006412901, 
    0.0006768624, 0.0007085879, 0.0006963965, 0.0006630807, 0.0006353445, 
    0.0006324677, 0.0006354088, 0.0006479817, 0.0006967937, 0.0006848734, 
    0.000624601, 0.000570178, 0.0005796989, 0.0006237268, 0.0006887352, 
    0.0007588943, 0.0007886172, 0.0007880926, 0.0007821957, 0.0007759968, 
    0.0007937511, 0.0008240463, 0.0008422297,
  0.0005208096, 0.0005406304, 0.0005532664, 0.0005586387, 0.0005657116, 
    0.0005738023, 0.0005795078, 0.0005740402, 0.0005674281, 0.000560625, 
    0.0005575414, 0.000572657, 0.0006035403, 0.0006287966, 0.0006329929, 
    0.0006461218, 0.0006856038, 0.0007283285, 0.0007361805, 0.0007021341, 
    0.0006483793, 0.0006014109, 0.0005563975, 0.0005192987, 0.0005026415, 
    0.00052518, 0.000576583, 0.0005895689, 0.0005582408, 0.0005386269, 
    0.0005472733, 0.000538484, 0.000500178, 0.000453718, 0.0004185429, 
    0.0003823671, 0.000353042, 0.0003633574, 0.0003884868, 0.0004193536, 
    0.000476304, 0.0005658381, 0.0006851903, 0.000769956, 0.0008017938, 
    0.0007964214, 0.0006774175, 0.0004602186, 0.0003034184, 0.0002029329, 
    0.000153183, 0.000146444, 0.0001156717, 8.477271e-005, 9.020837e-005, 
    0.0001158789, 0.0001508943, 0.0001988327, 0.0002478673, 0.0002782098, 
    0.0002885894, 0.0003082189, 0.0003262279, 0.0003486709, 0.0003987863, 
    0.000469517, 0.0005302182, 0.0005583833, 0.0005550771, 0.00055255, 
    0.0005614194, 0.0005778703, 0.0005826387, 0.0006043664, 0.0006197048, 
    0.0006080861, 0.0006102161, 0.0006319596, 0.0006316416, 0.000614793, 
    0.0006033652, 0.0006262846, 0.0007003383, 0.0006212625, 0.0005638991, 
    0.0005697168, 0.000594194, 0.0006086268, 0.0006034288, 0.0005988039, 
    0.0005983268, 0.0005851509, 0.0005690497, 0.0005536003, 0.0005339861, 
    0.0005175353,
  0.0005678572, 0.0005777911, 0.0006001545, 0.0006270639, 0.0006506837, 
    0.0006715371, 0.0006916597, 0.0007069027, 0.0007000519, 0.0006875428, 
    0.0006666416, 0.000662731, 0.0006780694, 0.0006957757, 0.0007179333, 
    0.0007710368, 0.0008650371, 0.0009252299, 0.0008874331, 0.0008283528, 
    0.0008416567, 0.0008865749, 0.0008965405, 0.0008686767, 0.000845185, 
    0.0008578529, 0.0008916128, 0.0008901665, 0.0008573285, 0.0008161296, 
    0.0007769335, 0.0007217634, 0.000679675, 0.0006831554, 0.0006805491, 
    0.0006319592, 0.000562659, 0.0005357661, 0.0005648057, 0.0006545307, 
    0.0007704338, 0.0008411971, 0.0008368734, 0.0008269073, 0.0008797408, 
    0.0008774842, 0.0007840553, 0.0005671582, 0.0004535913, 0.0003744205, 
    0.0003636917, 0.0003935578, 0.0004110895, 0.0003906805, 0.0003826381, 
    0.0004080534, 0.0004413049, 0.0004781964, 0.0005108118, 0.0005261181, 
    0.0005340171, 0.0005483073, 0.000563581, 0.0005713855, 0.0005841167, 
    0.0006093262, 0.0006212941, 0.0006210566, 0.0006136498, 0.0005835448, 
    0.0005622143, 0.0005762498, 0.0005873283, 0.0006021261, 0.0006208499, 
    0.0006717765, 0.0006212625, 0.0005933996, 0.0006848085, 0.0007475931, 
    0.000676068, 0.0006156513, 0.0006070207, 0.0005682376, 0.0005781245, 
    0.000620245, 0.0006742706, 0.000700783, 0.0006849519, 0.0006557857, 
    0.0006400342, 0.000635393, 0.0006273345, 0.0006234082, 0.0006016169, 
    0.0005754861,
  0.0007543792, 0.0007717041, 0.0007885052, 0.0008061319, 0.0008401787, 
    0.0008984804, 0.000990923, 0.001070571, 0.001087293, 0.001096591, 
    0.001124644, 0.001137217, 0.001126981, 0.001085575, 0.001062432, 
    0.001088405, 0.001155496, 0.001229643, 0.001251085, 0.001394407, 
    0.001610684, 0.001672626, 0.001554323, 0.001385744, 0.00129346, 
    0.001250338, 0.001176937, 0.001059842, 0.0009601042, 0.0008594277, 
    0.0007513128, 0.0007000524, 0.0007196348, 0.0007473235, 0.0007461794, 
    0.0007056314, 0.000657741, 0.0006697257, 0.0007310472, 0.000831787, 
    0.001049113, 0.001128284, 0.001057188, 0.001032312, 0.001133196, 
    0.001056965, 0.0009834208, 0.0008496684, 0.0007035811, 0.0006142855, 
    0.0006420691, 0.0007169326, 0.000748897, 0.0007323823, 0.0007227659, 
    0.0007003224, 0.000685541, 0.0007208427, 0.0007556202, 0.0007811468, 
    0.0007787626, 0.0007706727, 0.000767637, 0.0007508197, 0.0007388354, 
    0.0007539671, 0.0007391693, 0.0006972551, 0.0006720466, 0.0006701709, 
    0.0006853184, 0.0006900234, 0.0006825686, 0.0006806133, 0.0006953957, 
    0.0007094145, 0.0006125998, 0.0005674595, 0.0006256974, 0.0007908111, 
    0.0007705931, 0.0006824574, 0.000647855, 0.0006374912, 0.0006374274, 
    0.0006858739, 0.0007949588, 0.0008701086, 0.0008726353, 0.0008556289, 
    0.0008499217, 0.0008289726, 0.0008070855, 0.0007919222, 0.0007710685, 
    0.0007544109,
  0.001125089, 0.001132623, 0.001091647, 0.001063386, 0.001131304, 
    0.00131247, 0.001557183, 0.001754958, 0.001886407, 0.002018984, 
    0.002111555, 0.002067145, 0.001910471, 0.001739223, 0.001641917, 
    0.001632412, 0.001628486, 0.001628295, 0.001667905, 0.00170486, 
    0.00167385, 0.001545548, 0.001353351, 0.001190289, 0.001086115, 
    0.0009975675, 0.0009302376, 0.0008714595, 0.0008366504, 0.0008433261, 
    0.0008563916, 0.0008379221, 0.0008238712, 0.0007849932, 0.000769353, 
    0.0007948796, 0.0008084695, 0.0008834279, 0.0009496766, 0.001036159, 
    0.001234078, 0.001307813, 0.001316635, 0.001320815, 0.001396982, 
    0.001468905, 0.00118506, 0.001177764, 0.001140825, 0.001148439, 
    0.00122931, 0.001189494, 0.001039417, 0.0009799716, 0.0009781914, 
    0.0008960804, 0.0008515436, 0.0008873702, 0.0009341156, 0.0009793201, 
    0.0009565591, 0.0009077471, 0.0009228629, 0.0009082239, 0.0008773883, 
    0.0008705538, 0.0008509238, 0.0008346797, 0.0008497159, 0.0008518775, 
    0.0008647996, 0.0008377153, 0.0008135396, 0.0008236165, 0.0008127452, 
    0.0008073729, 0.0007460201, 0.0005635815, 0.0006067981, 0.0008468549, 
    0.0009039324, 0.0008647679, 0.000893712, 0.0009892699, 0.001031804, 
    0.001051577, 0.001080934, 0.001082047, 0.001054836, 0.001059381, 
    0.001092299, 0.001115393, 0.001126266, 0.00109071, 0.001073099, 
    0.001098005,
  0.001254915, 0.001186585, 0.001145561, 0.001176588, 0.001327618, 
    0.001537998, 0.001608173, 0.001719849, 0.001828854, 0.001897519, 
    0.001743659, 0.001605075, 0.001515429, 0.001442553, 0.001393994, 
    0.001371218, 0.001352827, 0.001328429, 0.001295654, 0.001249766, 
    0.00114065, 0.001003051, 0.0009178407, 0.0008980185, 0.0009070002, 
    0.0009152652, 0.000945067, 0.001003321, 0.001053024, 0.00115931, 
    0.001135325, 0.001040323, 0.001019057, 0.0009507732, 0.000945162, 
    0.001035141, 0.001040259, 0.001081077, 0.001090645, 0.0009489139, 
    0.001412097, 0.001688505, 0.001727922, 0.001669701, 0.001665632, 
    0.00166088, 0.001619648, 0.001217517, 0.00138832, 0.001321499, 
    0.001201924, 0.001129301, 0.00102915, 0.001037336, 0.001054453, 
    0.001001636, 0.0009986153, 0.001031914, 0.00104158, 0.001071142, 
    0.001064419, 0.001039687, 0.001070475, 0.00107634, 0.001058919, 
    0.001043231, 0.001000062, 0.001031916, 0.001068187, 0.001032853, 
    0.001025716, 0.0009965021, 0.0009363098, 0.000893903, 0.0008419277, 
    0.0008679312, 0.0007877741, 0.0006477432, 0.0006444524, 0.0007160106, 
    0.0008754334, 0.001037097, 0.001362745, 0.001551684, 0.001554878, 
    0.001445809, 0.001332783, 0.00132916, 0.001322786, 0.001252564, 
    0.001185345, 0.001173297, 0.001208678, 0.001210935, 0.00125536, 
    0.001312009,
  0.001206661, 0.001177509, 0.001179401, 0.001206169, 0.001309689, 
    0.001385269, 0.001600544, 0.001643413, 0.001717863, 0.001782361, 
    0.001388097, 0.001361045, 0.001356754, 0.001317224, 0.001305271, 
    0.001254393, 0.001217326, 0.001190258, 0.00112633, 0.001068586, 
    0.001049703, 0.001102328, 0.00116082, 0.001171629, 0.001249147, 
    0.001289106, 0.001260829, 0.001296417, 0.001323088, 0.00129432, 
    0.001121276, 0.001047223, 0.001053134, 0.0010391, 0.001068823, 
    0.001110419, 0.001060716, 0.0009670178, 0.0009989501, 0.0009611845, 
    0.001235462, 0.001969107, 0.002234244, 0.002174703, 0.002006364, 
    0.001923808, 0.001781058, 0.001538349, 0.001328191, 0.001086197, 
    0.0009764284, 0.0009949608, 0.001019009, 0.001095144, 0.001141906, 
    0.001148613, 0.001188493, 0.00122238, 0.001233808, 0.001214052, 
    0.001184456, 0.001183487, 0.001219059, 0.001249719, 0.001305509, 
    0.001344833, 0.001283257, 0.001197681, 0.001148202, 0.001064564, 
    0.0009974577, 0.0009316374, 0.0009121345, 0.0009270757, 0.0008954769, 
    0.0008258754, 0.0006710608, 0.0006371578, 0.0007149447, 0.0007386608, 
    0.0008449159, 0.001150553, 0.001659593, 0.00187773, 0.001763034, 
    0.001592151, 0.001404295, 0.001373173, 0.001416486, 0.001412368, 
    0.001386905, 0.001317605, 0.001286405, 0.001252279, 0.001252485, 
    0.001264914,
  0.001099102, 0.001106081, 0.001081238, 0.001177845, 0.001246398, 
    0.001013732, 0.001043169, 0.001251244, 0.001642855, 0.001904114, 
    0.001808317, 0.001827772, 0.001871848, 0.001763129, 0.00169855, 
    0.001670449, 0.00165724, 0.001649261, 0.001605297, 0.001615152, 
    0.001613006, 0.001623401, 0.001634003, 0.001600767, 0.001582392, 
    0.001556707, 0.001512934, 0.001473149, 0.001415039, 0.001285531, 
    0.001209714, 0.0009081759, 0.0008853199, 0.0009956439, 0.001166002, 
    0.001261067, 0.00110403, 0.001149711, 0.001405105, 0.001515492, 
    0.001673531, 0.002123795, 0.002112716, 0.002141913, 0.002110537, 
    0.001958872, 0.001766706, 0.001523837, 0.00135003, 0.001299836, 
    0.001339858, 0.001384124, 0.001377941, 0.001374587, 0.001393724, 
    0.00142572, 0.001368103, 0.001306273, 0.001365575, 0.001381612, 
    0.001397333, 0.001444842, 0.001504811, 0.001598701, 0.001615088, 
    0.001527159, 0.001341891, 0.001087292, 0.0009002769, 0.0008094544, 
    0.0007663965, 0.000811697, 0.0008396404, 0.0008556135, 0.0008063568, 
    0.0007633455, 0.0007889047, 0.0007929727, 0.0008342336, 0.00103147, 
    0.001182691, 0.001401814, 0.001582567, 0.00193317, 0.001908644, 
    0.001642935, 0.001461545, 0.001503348, 0.001526348, 0.001467713, 
    0.001489728, 0.001423098, 0.00137446, 0.001369676, 0.001295623, 
    0.001194963,
  0.001101582, 0.001086355, 0.001218279, 0.001527207, 0.001707038, 
    0.001316524, 0.001266805, 0.0014426, 0.001895484, 0.002212898, 
    0.002131996, 0.002143995, 0.002237345, 0.002190615, 0.002092989, 
    0.002105991, 0.002101811, 0.00198443, 0.001932184, 0.001986528, 
    0.001991327, 0.00192581, 0.001865921, 0.001841999, 0.001751718, 
    0.001653633, 0.001626214, 0.001527764, 0.001517448, 0.001521039, 
    0.001505748, 0.00119555, 0.001396219, 0.001659131, 0.00160145, 
    0.001543053, 0.001650215, 0.00188485, 0.001918563, 0.001956248, 
    0.002038138, 0.002122426, 0.002031287, 0.002000833, 0.002033655, 
    0.002012325, 0.00198799, 0.001946759, 0.001886661, 0.001882672, 
    0.001856732, 0.001741163, 0.001632873, 0.001605026, 0.001605073, 
    0.001622638, 0.001561189, 0.001540049, 0.001578578, 0.001664137, 
    0.001752575, 0.001811178, 0.00184435, 0.001842395, 0.001682401, 
    0.001362522, 0.001122545, 0.0008506859, 0.0006787861, 0.0006599501, 
    0.0007413626, 0.0009033289, 0.0008632578, 0.0008577909, 0.0008254461, 
    0.0009469278, 0.001377051, 0.0008457093, 0.0009058551, 0.001468682, 
    0.001677616, 0.0017205, 0.001649085, 0.001834879, 0.002161114, 
    0.001898075, 0.001716637, 0.001750239, 0.001740495, 0.001660164, 
    0.001633048, 0.00155197, 0.001495576, 0.001399207, 0.001255393, 
    0.001144117,
  0.001390242, 0.001505573, 0.001813722, 0.002116164, 0.00152514, 
    0.001344673, 0.001456141, 0.001590816, 0.001871196, 0.002188945, 
    0.002419623, 0.002425727, 0.002549594, 0.002455417, 0.002406907, 
    0.002357508, 0.002357732, 0.002284265, 0.002216918, 0.002208527, 
    0.002124063, 0.002072008, 0.002037406, 0.001972826, 0.001874661, 
    0.001828551, 0.001845749, 0.00185678, 0.001893559, 0.002007413, 
    0.002159715, 0.001942913, 0.002052443, 0.002298617, 0.002177501, 
    0.002042557, 0.002163625, 0.002419797, 0.002320504, 0.002270373, 
    0.002301129, 0.00236013, 0.002495376, 0.002576057, 0.002551707, 
    0.002444704, 0.002365629, 0.002325559, 0.002249838, 0.002168458, 
    0.002054079, 0.001919501, 0.001861024, 0.00190696, 0.001970569, 
    0.001978437, 0.001989435, 0.002037883, 0.002095039, 0.002241858, 
    0.002280306, 0.002211944, 0.002109122, 0.001853363, 0.001563652, 
    0.001227958, 0.001024669, 0.0009522839, 0.0008991482, 0.0009613745, 
    0.001000809, 0.0009995224, 0.0009414116, 0.0009793835, 0.0009856457, 
    0.001299581, 0.002118325, 0.001234475, 0.0008668024, 0.002025676, 
    0.002085949, 0.001836038, 0.001816949, 0.001832002, 0.002075538, 
    0.002132504, 0.002008685, 0.001918166, 0.001898027, 0.001856764, 
    0.00177292, 0.001622573, 0.001505447, 0.001415753, 0.001323898, 
    0.001285115,
  0.001938049, 0.002105483, 0.002424439, 0.00250369, 0.001825102, 
    0.001649722, 0.001899949, 0.001929434, 0.001919087, 0.002142693, 
    0.002552629, 0.002524734, 0.002182746, 0.002248725, 0.002469896, 
    0.002439745, 0.002384973, 0.002347779, 0.002357475, 0.002428222, 
    0.00242765, 0.002443862, 0.002450871, 0.002349861, 0.002296249, 
    0.002287301, 0.002289829, 0.002324144, 0.002410991, 0.002648011, 
    0.0028452, 0.002596751, 0.002065078, 0.001877728, 0.002028568, 
    0.001729321, 0.001871388, 0.002431989, 0.002723082, 0.002629749, 
    0.002725101, 0.002954571, 0.003064705, 0.003047553, 0.00291973, 
    0.002754888, 0.00261484, 0.002536749, 0.002417366, 0.00227619, 
    0.002184814, 0.002211612, 0.002304278, 0.002405813, 0.002503818, 
    0.002590617, 0.002642449, 0.002710097, 0.002760816, 0.002791191, 
    0.00269735, 0.002544764, 0.0023361, 0.002007875, 0.001792581, 
    0.001548186, 0.001420776, 0.001394201, 0.001325727, 0.001293905, 
    0.001178305, 0.001151809, 0.001208679, 0.001228499, 0.001306606, 
    0.001835655, 0.002385005, 0.001240166, 0.001139298, 0.002372305, 
    0.002036151, 0.002050743, 0.002402537, 0.00182229, 0.001885026, 
    0.002100873, 0.002186736, 0.002224104, 0.002195111, 0.002051043, 
    0.001921887, 0.001824483, 0.001748602, 0.001737189, 0.001740321, 
    0.001779549,
  0.002475509, 0.002595814, 0.002816605, 0.002761975, 0.002094292, 
    0.001763017, 0.001834098, 0.001805488, 0.002026947, 0.002034673, 
    0.002350386, 0.002744285, 0.002288748, 0.002201915, 0.002444196, 
    0.002545144, 0.002534337, 0.002578616, 0.00267311, 0.002748498, 
    0.002847505, 0.002886303, 0.002858218, 0.002852781, 0.002839081, 
    0.002847761, 0.002977381, 0.003072366, 0.003174553, 0.00337241, 
    0.003483223, 0.003322482, 0.003027494, 0.003214257, 0.003079661, 
    0.00253214, 0.00269878, 0.003263353, 0.002943953, 0.00297436, 0.00320944, 
    0.003383692, 0.003337726, 0.003190892, 0.002998587, 0.002856804, 
    0.002736481, 0.00267683, 0.002631927, 0.002633853, 0.002690978, 
    0.002782736, 0.002921432, 0.003029371, 0.003100196, 0.003143335, 
    0.003141094, 0.003108226, 0.003069555, 0.002932161, 0.002799647, 
    0.002724085, 0.002552249, 0.002345728, 0.002212659, 0.002064236, 
    0.00195717, 0.001892478, 0.001774686, 0.001733981, 0.00170006, 
    0.00171217, 0.001766419, 0.001811178, 0.001950209, 0.002253365, 
    0.001776544, 0.001344816, 0.00180738, 0.002549433, 0.002036626, 
    0.002029554, 0.001983492, 0.001933616, 0.001790675, 0.00190289, 
    0.002344283, 0.002467417, 0.002471376, 0.00242258, 0.002384273, 
    0.002361305, 0.00236687, 0.002360637, 0.00238092, 0.002387326,
  0.002909636, 0.002960705, 0.003034728, 0.003052037, 0.002151895, 
    0.001583537, 0.002017856, 0.001868748, 0.002050169, 0.001974719, 
    0.002165119, 0.002842022, 0.00267807, 0.002501734, 0.002491055, 
    0.00251429, 0.00261271, 0.002703533, 0.002897779, 0.003009615, 
    0.00310147, 0.003132926, 0.003114933, 0.003185298, 0.0032281, 
    0.003345275, 0.003465408, 0.003502045, 0.003628742, 0.003761461, 
    0.003774891, 0.003867857, 0.003846798, 0.003661862, 0.003474055, 
    0.003341253, 0.003473036, 0.003492936, 0.003138105, 0.003300009, 
    0.003473897, 0.003495639, 0.003381021, 0.003164012, 0.002991095, 
    0.002939153, 0.002852367, 0.002865864, 0.002919493, 0.002965683, 
    0.003026702, 0.003111755, 0.003179958, 0.003240166, 0.003300026, 
    0.003257046, 0.003209235, 0.003131349, 0.003126884, 0.003092822, 
    0.002994627, 0.002936024, 0.002857948, 0.002762424, 0.002664875, 
    0.002571004, 0.002460758, 0.002400645, 0.00241746, 0.002397576, 
    0.002376756, 0.002354376, 0.00237275, 0.002363277, 0.002405158, 
    0.002566949, 0.002100365, 0.001964339, 0.002179615, 0.001914286, 
    0.001590069, 0.001484435, 0.001954659, 0.002237979, 0.001823163, 
    0.001965818, 0.002560798, 0.002737245, 0.002724307, 0.002818624, 
    0.002851922, 0.0028449, 0.002893044, 0.002860808, 0.002871585, 0.002842133,
  0.003140748, 0.003086004, 0.003156941, 0.003220232, 0.002531203, 
    0.002109123, 0.002422898, 0.002358492, 0.0021765, 0.002256308, 
    0.002264046, 0.002854532, 0.002713913, 0.00259478, 0.002634408, 
    0.00272499, 0.002942413, 0.003011188, 0.003133068, 0.003166988, 
    0.003199905, 0.003274275, 0.003296958, 0.003299899, 0.003326824, 
    0.003414972, 0.003480395, 0.003557086, 0.003564922, 0.003608394, 
    0.003771076, 0.003762744, 0.003793504, 0.003837453, 0.00375687, 
    0.003558341, 0.003510628, 0.003400143, 0.00307308, 0.003327949, 
    0.003583407, 0.003496164, 0.003347233, 0.003211318, 0.003071364, 
    0.003011584, 0.002904853, 0.002929902, 0.002873637, 0.00281368, 
    0.00281891, 0.002866674, 0.002891611, 0.002948975, 0.003076147, 
    0.003057105, 0.003099544, 0.00310104, 0.003065342, 0.003038447, 
    0.002977157, 0.002964983, 0.002962139, 0.002891503, 0.002858026, 
    0.002842339, 0.0028439, 0.002848905, 0.00288821, 0.002902165, 
    0.002881804, 0.002868915, 0.002859857, 0.002865912, 0.002904136, 
    0.002643212, 0.001836037, 0.001448242, 0.001462373, 0.001312375, 
    0.001217612, 0.001430997, 0.001651836, 0.002297139, 0.002324479, 
    0.002173845, 0.002361942, 0.002903741, 0.002984535, 0.003086768, 
    0.003129095, 0.003137121, 0.003125453, 0.003053229, 0.003090629, 
    0.003063209,
  0.003191225, 0.003139013, 0.003243281, 0.003166193, 0.003342, 0.002873889, 
    0.002913292, 0.002887481, 0.002631975, 0.00221417, 0.002288112, 
    0.002680758, 0.002791589, 0.002638685, 0.002785008, 0.002868691, 
    0.002989175, 0.003147565, 0.003178433, 0.003154749, 0.003205245, 
    0.003299976, 0.003297212, 0.003281744, 0.00328335, 0.003237639, 
    0.003326854, 0.003243247, 0.003047856, 0.003353206, 0.003422253, 
    0.00339237, 0.003363743, 0.00339593, 0.003459351, 0.003470207, 
    0.003289819, 0.003046393, 0.002783959, 0.003063703, 0.003526822, 
    0.003354987, 0.003201526, 0.003129905, 0.002894808, 0.0027893, 
    0.002743617, 0.002746621, 0.00274465, 0.002832802, 0.002870996, 
    0.002888782, 0.002954919, 0.003047585, 0.003134036, 0.003138026, 
    0.003162201, 0.003156129, 0.003154667, 0.003148692, 0.003155433, 
    0.003106557, 0.003083698, 0.003047349, 0.00308203, 0.003054406, 
    0.003070906, 0.003057219, 0.003058506, 0.003089152, 0.003052801, 
    0.003000364, 0.002977539, 0.002986442, 0.003004482, 0.002665051, 
    0.001631094, 0.002107216, 0.001940974, 0.001404675, 0.001438245, 
    0.001782425, 0.00222253, 0.002513655, 0.002692342, 0.002631163, 
    0.002410917, 0.002835456, 0.003034664, 0.003206501, 0.003238147, 
    0.003269697, 0.003269363, 0.003265802, 0.003292806, 0.003246125,
  0.003231391, 0.003256602, 0.0031626, 0.002640512, 0.003346928, 0.003312707, 
    0.003060094, 0.002841625, 0.002886748, 0.002490989, 0.002466194, 
    0.002771975, 0.002704723, 0.00277709, 0.002834249, 0.00304088, 
    0.003182482, 0.003331829, 0.003341157, 0.003362775, 0.00339655, 
    0.003408391, 0.003413446, 0.003372105, 0.003368037, 0.003249271, 
    0.003141729, 0.002550896, 0.002806006, 0.003356829, 0.001870656, 
    0.002472539, 0.002758894, 0.003153777, 0.003250511, 0.003203845, 
    0.002733544, 0.002704997, 0.002950361, 0.003282698, 0.003507622, 
    0.003169704, 0.003051654, 0.003027145, 0.002920236, 0.00287934, 
    0.002977697, 0.002977284, 0.002992462, 0.003128886, 0.003228737, 
    0.003363522, 0.003439942, 0.003512772, 0.003545197, 0.003493987, 
    0.003457857, 0.003348885, 0.003289774, 0.003187096, 0.003147675, 
    0.003057169, 0.00304204, 0.003025716, 0.003029468, 0.003007088, 
    0.003056217, 0.003098864, 0.00311622, 0.003068537, 0.003079295, 
    0.003017133, 0.003001969, 0.002921656, 0.002943605, 0.003037794, 
    0.002388199, 0.00287699, 0.002465719, 0.002195351, 0.002620816, 
    0.002532268, 0.002329884, 0.002967479, 0.003004083, 0.002879361, 
    0.002745384, 0.002871016, 0.003061542, 0.003212634, 0.003175789, 
    0.003212653, 0.003287833, 0.003280094, 0.003201224, 0.00323109,
  0.003105426, 0.003265452, 0.003205849, 0.002619499, 0.003037954, 
    0.003241641, 0.002793988, 0.002550231, 0.002922115, 0.003014875, 
    0.002834359, 0.002757018, 0.002631087, 0.002744015, 0.002837397, 
    0.003014192, 0.003225779, 0.003280727, 0.003283987, 0.003247285, 
    0.003260843, 0.003235348, 0.003315743, 0.003308639, 0.003432646, 
    0.003286211, 0.003042404, 0.002540007, 0.003104918, 0.003301168, 
    0.002604399, 0.002379222, 0.002816655, 0.003040258, 0.00305113, 
    0.003006894, 0.002967142, 0.002966857, 0.003113708, 0.003238272, 
    0.003119001, 0.002999313, 0.003037779, 0.003029687, 0.003034251, 
    0.002996547, 0.003003987, 0.002927771, 0.00292399, 0.002975233, 
    0.003052592, 0.003178908, 0.003253039, 0.003311152, 0.00336354, 
    0.003316078, 0.003323866, 0.003245234, 0.00323678, 0.00318253, 
    0.003153205, 0.003087688, 0.003055329, 0.003017196, 0.003091136, 
    0.003083762, 0.003094411, 0.003104456, 0.003105842, 0.00301473, 
    0.003012395, 0.002887225, 0.002768476, 0.002679452, 0.002712099, 
    0.002864879, 0.002628716, 0.002793068, 0.002933752, 0.002854053, 
    0.002874083, 0.002017728, 0.001850886, 0.002843786, 0.002741521, 
    0.002812713, 0.002805196, 0.002824634, 0.00302276, 0.003120957, 
    0.003084382, 0.003035394, 0.003069839, 0.003109479, 0.003078962, 
    0.003128823,
  0.002952585, 0.003297608, 0.002851542, 0.002868202, 0.0031121, 0.003171818, 
    0.00297118, 0.002816416, 0.003091456, 0.003146863, 0.002959546, 
    0.002750055, 0.002433436, 0.002851367, 0.00299523, 0.003002143, 
    0.003300533, 0.003369657, 0.003310975, 0.003141887, 0.003147515, 
    0.003034631, 0.003031882, 0.003175776, 0.00341359, 0.003278581, 
    0.002607895, 0.002914738, 0.003076784, 0.003052194, 0.002989411, 
    0.002898844, 0.00292011, 0.003049303, 0.002984548, 0.002969097, 
    0.003033996, 0.003049906, 0.003065022, 0.002972165, 0.002966112, 
    0.003070187, 0.003103932, 0.003121495, 0.003138946, 0.00308721, 
    0.003050748, 0.003037222, 0.00300594, 0.002991287, 0.003001794, 
    0.002951041, 0.00299472, 0.002938945, 0.002920795, 0.002936928, 
    0.002981719, 0.002937755, 0.002964569, 0.003021838, 0.003067249, 
    0.003098497, 0.003116062, 0.003091503, 0.003218152, 0.003201971, 
    0.003281457, 0.003316252, 0.003322657, 0.003229579, 0.003108144, 
    0.003058314, 0.002949961, 0.002800506, 0.002743538, 0.002825286, 
    0.002615554, 0.002815047, 0.003042899, 0.002019572, 0.002347017, 
    0.002630148, 0.002733747, 0.002766412, 0.002811741, 0.002934242, 
    0.002860095, 0.00294777, 0.002998678, 0.003067564, 0.003214242, 
    0.003190238, 0.003151521, 0.003141601, 0.002727645, 0.002763536,
  0.003018832, 0.002926994, 0.003008025, 0.003020789, 0.003089469, 
    0.003278837, 0.003156433, 0.003046442, 0.0033239, 0.003196074, 
    0.002838778, 0.003205324, 0.002410328, 0.00250835, 0.003174409, 
    0.002927553, 0.003243264, 0.003409935, 0.003469093, 0.003408456, 
    0.003229849, 0.003059333, 0.003204353, 0.003305046, 0.003325311, 
    0.003365843, 0.003164997, 0.003136724, 0.003191464, 0.003226655, 
    0.003310831, 0.003009278, 0.003057599, 0.002976552, 0.002947705, 
    0.00297452, 0.002960164, 0.003015462, 0.00307955, 0.003119191, 
    0.003083635, 0.003067199, 0.003121305, 0.003199918, 0.003203591, 
    0.003160659, 0.0031293, 0.003112165, 0.003096892, 0.0030514, 0.00306035, 
    0.003004927, 0.003032615, 0.002964856, 0.002971945, 0.00293852, 
    0.002941603, 0.002931811, 0.002932526, 0.002944622, 0.0029705, 
    0.002959881, 0.003019612, 0.003014447, 0.003162615, 0.003172675, 
    0.003248619, 0.003310338, 0.003354192, 0.0032463, 0.003141666, 
    0.003173534, 0.002797039, 0.002664732, 0.002545524, 0.002629464, 
    0.002651939, 0.002715183, 0.002855755, 0.002576839, 0.002777714, 
    0.002758687, 0.002703885, 0.002670249, 0.002636062, 0.002704775, 
    0.002685968, 0.002789507, 0.002781004, 0.002862765, 0.002982751, 
    0.002971103, 0.003029134, 0.002929697, 0.003011061, 0.003047856,
  0.003189223, 0.003129825, 0.003249779, 0.003314836, 0.002652429, 
    0.002575913, 0.002548925, 0.003109798, 0.003541144, 0.003133863, 
    0.002849126, 0.001743485, 0.001941419, 0.001967011, 0.003627928, 
    0.0030655, 0.003090486, 0.0033681, 0.003479123, 0.003493747, 0.003067026, 
    0.003014063, 0.003330491, 0.003508462, 0.003427353, 0.00338717, 
    0.003392925, 0.003016289, 0.002993356, 0.003067803, 0.003278024, 
    0.003153173, 0.003036365, 0.003088119, 0.002835536, 0.002973486, 
    0.002978936, 0.003083745, 0.003104663, 0.003171848, 0.003095396, 
    0.003099354, 0.003188744, 0.003193069, 0.003192879, 0.003165541, 
    0.003101423, 0.002992354, 0.002994595, 0.00299488, 0.002978828, 
    0.002953919, 0.002917076, 0.002890676, 0.002941111, 0.00289988, 
    0.002876848, 0.002833804, 0.002831534, 0.002819708, 0.002835061, 
    0.002812728, 0.002881648, 0.00290517, 0.003011694, 0.002998712, 
    0.003012156, 0.003257457, 0.003458254, 0.003291123, 0.003249303, 
    0.002996229, 0.002597565, 0.002319343, 0.00250574, 0.002550421, 
    0.002644088, 0.00263509, 0.002710065, 0.002732366, 0.002703771, 
    0.00259761, 0.00257043, 0.002539596, 0.002529694, 0.002499573, 
    0.002513196, 0.002551246, 0.002558606, 0.002600996, 0.002610819, 
    0.002885098, 0.002800805, 0.003470922, 0.00346908, 0.00323702,
  0.002342535, 0.002129229, 0.00193584, 0.001470256, 0.0004686275, 
    0.0009620897, 0.001330877, 0.001546358, 0.002040442, 0.001998162, 
    0.002143772, 0.002165962, 0.001105969, 0.001497944, 0.002723511, 
    0.003378892, 0.003132813, 0.003296955, 0.003376683, 0.003455313, 
    0.003102707, 0.003277898, 0.003480041, 0.003732467, 0.003714407, 
    0.003421677, 0.002986044, 0.003018498, 0.003063655, 0.002960466, 
    0.002988378, 0.003047729, 0.002907379, 0.002746813, 0.002809532, 
    0.002978761, 0.003054278, 0.003133288, 0.003098814, 0.003040275, 
    0.00289177, 0.002880154, 0.002954638, 0.00294742, 0.002968622, 
    0.002965841, 0.002987426, 0.00291579, 0.002851576, 0.002826288, 
    0.002786711, 0.002732143, 0.00265949, 0.002588058, 0.0025378, 
    0.002457039, 0.002434311, 0.002368474, 0.002386609, 0.002385464, 
    0.002423629, 0.002466607, 0.002509508, 0.002445342, 0.002311891, 
    0.002198465, 0.002452223, 0.003017448, 0.00331614, 0.002990399, 
    0.00288303, 0.002346653, 0.001785556, 0.00241301, 0.002494883, 
    0.002524847, 0.002564091, 0.002539692, 0.00252901, 0.002527738, 
    0.002513528, 0.002471043, 0.002466228, 0.002408704, 0.002441144, 
    0.0023645, 0.002320074, 0.002244719, 0.002243686, 0.002157124, 
    0.002242429, 0.0024743, 0.002145919, 0.0009107199, 0.0006829016, 
    0.001768391,
  0.0006464571, 0.001181467, 0.0008926787, 0.001187746, 0.0002694684, 
    0.001131114, 0.0008551665, 0.0006832196, 0.0009428104, 0.001320196, 
    0.002539737, 0.001822243, 0.001282335, 0.0009544443, 0.002012928, 
    0.004067318, 0.003528461, 0.003343351, 0.003440516, 0.003552476, 
    0.003205992, 0.003784822, 0.00382866, 0.003397934, 0.003613938, 
    0.003357703, 0.003184501, 0.002947498, 0.002789998, 0.002876639, 
    0.0028538, 0.002882123, 0.002867231, 0.002769621, 0.002735861, 
    0.002944143, 0.002939407, 0.002905011, 0.00286804, 0.002795786, 
    0.00268613, 0.002653576, 0.002687303, 0.002675908, 0.002603253, 
    0.002600251, 0.00262147, 0.002627382, 0.002569811, 0.002500035, 
    0.002477815, 0.002414824, 0.002344729, 0.002294436, 0.002264031, 
    0.002183637, 0.002122155, 0.002041301, 0.001957583, 0.001904543, 
    0.001889476, 0.001859213, 0.001895881, 0.001914827, 0.001712187, 
    0.001512535, 0.001712572, 0.002305422, 0.002286522, 0.002555807, 
    0.002740903, 0.002247676, 0.001654699, 0.002503514, 0.002492182, 
    0.0025141, 0.002512766, 0.002398452, 0.002348863, 0.002425155, 
    0.002452748, 0.002346032, 0.002325512, 0.002268991, 0.002228347, 
    0.002194365, 0.002149113, 0.002031892, 0.001980218, 0.001849344, 
    0.001855145, 0.002124366, 0.001117143, -0.0005465904, -0.001893498, 
    -0.000804448,
  0.001001732, 0.001123151, 0.0002901317, 0.0001006355, 0.0003944626, 
    0.0006222646, 0.0001223488, 0.0005121629, 0.0007176322, 0.001427134, 
    0.001989117, 0.00131956, 0.001525124, 0.001409682, 0.001730307, 
    0.00369742, 0.004054952, 0.003736153, 0.003526777, 0.003417484, 
    0.003695307, 0.004536748, 0.004783304, 0.003621113, 0.003034744, 
    0.003262782, 0.003156003, 0.002539629, 0.002617177, 0.002672633, 
    0.002708856, 0.003061289, 0.002718234, 0.002782177, 0.002824539, 
    0.002902057, 0.002814937, 0.002721572, 0.002662746, 0.002568491, 
    0.002512621, 0.002533382, 0.002554251, 0.002532808, 0.002477255, 
    0.002449919, 0.00238774, 0.002366791, 0.002368731, 0.002319725, 
    0.002287444, 0.002238329, 0.002145155, 0.00202771, 0.001972382, 
    0.00194862, 0.001855589, 0.001802199, 0.001713348, 0.001642823, 
    0.001587097, 0.001546328, 0.001613561, 0.001548108, 0.001400447, 
    0.001367243, 0.001571566, 0.002373911, 0.002710352, 0.002755252, 
    0.002853639, 0.002723144, 0.002473524, 0.002499525, 0.002445452, 
    0.002321126, 0.002244433, 0.002382921, 0.002454432, 0.002351424, 
    0.002357494, 0.002410514, 0.002409085, 0.002323364, 0.002216442, 
    0.002161749, 0.002082244, 0.001997734, 0.001902193, 0.001765657, 
    0.001703143, 0.001778674, 0.001314712, 0.001477965, 0.001060319, 
    0.0003534714,
  0.0003284053, 0.001085925, 0.001041404, 0.0004960457, 0.001358008, 
    0.001231567, 0.0005512624, 0.0004734267, 0.0009745997, 0.001107844, 
    0.001426196, 0.0009979638, 0.001414959, 0.001385156, 0.00208196, 
    0.00298164, 0.003076863, 0.003053341, 0.003632474, 0.004191358, 
    0.004955858, 0.004230127, 0.003801959, 0.0033273, 0.002781097, 
    0.002690196, 0.0024074, 0.00237787, 0.002874319, 0.00322729, 0.003097717, 
    0.003043627, 0.003183948, 0.002946654, 0.003087752, 0.003067775, 
    0.002891278, 0.002752379, 0.002616735, 0.002392842, 0.002269752, 
    0.002258515, 0.002259582, 0.002258852, 0.002251556, 0.002249647, 
    0.002178406, 0.002089715, 0.002082865, 0.002105117, 0.002125477, 
    0.002102272, 0.002057894, 0.00197877, 0.001879733, 0.001808159, 
    0.001707594, 0.001662898, 0.001627374, 0.001546455, 0.001462547, 
    0.00140458, 0.001397029, 0.001286101, 0.001310213, 0.001505859, 
    0.001759839, 0.002724085, 0.002958753, 0.002876559, 0.002960341, 
    0.002791686, 0.002677452, 0.002539011, 0.002528137, 0.002063472, 
    0.002044734, 0.002152232, 0.002229923, 0.002227204, 0.002312684, 
    0.002363754, 0.002336605, 0.002356235, 0.002287873, 0.002142786, 
    0.00205095, 0.002023929, 0.001967454, 0.00181299, 0.001653806, 
    0.001610065, 0.0018032, 0.001373029, 0.001256156, 1.339056e-005,
  0.001152031, 0.0007794932, -0.0004362194, 0.001082667, 0.001474357, 
    0.001720834, 0.00158786, 0.0009028036, 0.002234832, 0.001911538, 
    0.001645875, 0.001360439, 0.00179608, 0.002080878, 0.00162979, 
    0.001618457, 0.00197734, 0.002090843, 0.002306882, 0.003614432, 
    0.00348084, 0.002789729, 0.001999848, 0.002018761, 0.002209608, 
    0.002042667, 0.00219667, 0.002159159, 0.002585769, 0.00322888, 
    0.003440149, 0.003402864, 0.003249494, 0.002013771, 0.002496584, 
    0.002738547, 0.002706298, 0.002577997, 0.002541916, 0.002486443, 
    0.002318898, 0.002209083, 0.002160111, 0.00211068, 0.002073074, 
    0.002082562, 0.002064252, 0.002000373, 0.001977324, 0.00193131, 
    0.001910694, 0.00190305, 0.001897058, 0.001885565, 0.001844446, 
    0.001751017, 0.001643602, 0.001553273, 0.001465535, 0.001391991, 
    0.001369612, 0.00130562, 0.001274054, 0.001325917, 0.001450849, 
    0.002026487, 0.002317945, 0.002458311, 0.002766808, 0.002760151, 
    0.003039306, 0.002533445, 0.002646009, 0.002659488, 0.002677751, 
    0.002405478, 0.002198864, 0.002079273, 0.002106277, 0.002084486, 
    0.002072914, 0.002064331, 0.002063444, 0.002121427, 0.002050521, 
    0.001976626, 0.001960889, 0.001900475, 0.00186592, 0.001819095, 
    0.001687995, 0.001565194, 0.001608856, 0.001864282, 0.002193587, 
    0.001439405,
  0.002420211, 0.002298443, 0.001729689, 0.001753878, 0.001802819, 
    0.001747695, 0.001543769, 0.001603993, 0.002123761, 0.002028584, 
    0.002331551, 0.001987975, 0.001758536, 0.001983303, 0.00163966, 
    0.001487707, 0.002329517, 0.002184669, 0.002115878, 0.00181307, 
    0.001714874, 0.001496864, 0.001446446, 0.001406296, 0.001223302, 
    0.001705543, 0.001821954, 0.002154645, 0.002206796, 0.002392554, 
    0.002493772, 0.002692821, 0.002686589, 0.001938702, 0.00244135, 
    0.002373274, 0.002683885, 0.002784037, 0.002490054, 0.002451414, 
    0.002266002, 0.002089445, 0.002010989, 0.002025501, 0.001978341, 
    0.001926605, 0.001878142, 0.001858735, 0.001875059, 0.001819571, 
    0.001747617, 0.0017147, 0.001674597, 0.001677474, 0.001673151, 
    0.001647132, 0.001601467, 0.00150052, 0.001393486, 0.001314983, 
    0.00124422, 0.001202958, 0.001252501, 0.001358042, 0.002146062, 
    0.002221433, 0.002561641, 0.002489211, 0.002742649, 0.003148519, 
    0.003244916, 0.002880153, 0.002823233, 0.002829385, 0.002887003, 
    0.002795846, 0.002361719, 0.002166724, 0.002018651, 0.00185128, 
    0.001763497, 0.001738112, 0.001678221, 0.001659147, 0.00163068, 
    0.001523439, 0.00153571, 0.001564734, 0.001585873, 0.001553304, 
    0.001547646, 0.001502221, 0.001458765, 0.001613181, 0.001718831, 0.0025333,
  0.002441477, 0.001589308, 0.001569948, 0.001649753, 0.001635432, 
    0.001447304, 0.00227015, 0.002041077, 0.001508372, 0.0015277, 
    0.001988595, 0.001940181, 0.00179333, 0.002188372, 0.001814897, 
    0.001943247, 0.001203116, 0.001361982, 0.002344617, 0.002320441, 
    0.002119612, 0.001719356, 0.0008611598, 0.001138265, 0.001823258, 
    0.001642473, 0.001758091, 0.002153611, 0.002210259, 0.002172464, 
    0.002035626, 0.002010449, 0.002037501, 0.002009067, 0.002033114, 
    0.001784175, 0.001747172, 0.00206527, 0.002000293, 0.00208091, 
    0.002122665, 0.002006237, 0.001876013, 0.00185249, 0.001811084, 
    0.001760205, 0.001730228, 0.001707355, 0.001695291, 0.001633604, 
    0.001590753, 0.001530004, 0.00142467, 0.001421332, 0.001424829, 
    0.001405597, 0.001378037, 0.001307544, 0.001247351, 0.001168753, 
    0.001112024, 0.001140444, 0.001238117, 0.001811672, 0.001914763, 
    0.001838279, 0.001648832, 0.002099887, 0.002466481, 0.003117886, 
    0.003285654, 0.003164347, 0.00303727, 0.002985121, 0.002835361, 
    0.00284574, 0.002676575, 0.002304276, 0.002027027, 0.001693749, 
    0.001609937, 0.001613419, 0.00149761, 0.001305254, 0.00101049, 
    0.0006012367, 0.0005686209, 0.0009317799, 0.001175093, 0.001190051, 
    0.001252628, 0.001339381, 0.001360759, 0.001565291, 0.002171461, 
    0.002363913,
  0.001663201, 0.001429916, 0.001204913, 0.001740051, 0.001245284, 
    0.001403118, 0.001467634, 0.001530338, 0.001711329, 0.001569899, 
    0.001623305, 0.001655492, 0.001630791, 0.001656652, 0.001812593, 
    0.001567911, 0.001509674, 0.001079376, 0.001577608, 0.001810876, 
    0.002014375, 0.002091798, 0.001991502, 0.002091289, 0.001888967, 
    0.001451548, 0.001449911, 0.001721057, 0.001988626, 0.002008017, 
    0.001920327, 0.001931883, 0.001863377, 0.001861931, 0.001845051, 
    0.001714302, 0.001452104, 0.001486707, 0.001676138, 0.001689315, 
    0.001651422, 0.00147326, 0.001343655, 0.001260717, 0.001162298, 
    0.001094874, 0.001103679, 0.001147978, 0.001164555, 0.001165923, 
    0.001192164, 0.001190766, 0.001160884, 0.001166892, 0.00118606, 
    0.00119318, 0.001155496, 0.001070746, 0.001022569, 0.001045092, 
    0.001062942, 0.001097941, 0.001158944, 0.001404008, 0.001869924, 
    0.001844208, 0.001872913, 0.00228765, 0.002446963, 0.003106968, 
    0.003305872, 0.003209917, 0.003174313, 0.002985947, 0.002426664, 
    0.002811219, 0.002633389, 0.002229, 0.002052776, 0.00185163, 0.001481747, 
    0.001332116, 0.001215052, 0.0009827847, 0.0007583061, 0.0006132852, 
    0.0005618818, 0.0006523859, 0.0007266449, 0.0008194214, 0.0009844862, 
    0.00111417, 0.001165272, 0.001323804, 0.001639693, 0.001757519,
  0.001388829, 0.001260178, 0.001129366, 0.001126457, 0.001172614, 
    0.001301505, 0.001382455, 0.001496578, 0.001541592, 0.001629758, 
    0.001781106, 0.001636593, 0.001693908, 0.00192694, 0.001869036, 
    0.002109473, 0.002191806, 0.002145043, 0.002184749, 0.002227489, 
    0.002115576, 0.001900427, 0.00189499, 0.001914271, 0.001813198, 
    0.001994412, 0.001868097, 0.001818729, 0.001961382, 0.001998257, 
    0.001873358, 0.001945487, 0.00196844, 0.001899441, 0.001879589, 
    0.001972031, 0.001817791, 0.001371201, 0.001246492, 0.0009053778, 
    0.000920732, 0.0009660954, 0.0009421427, 0.0009240867, 0.0009213053, 
    0.0008859243, 0.000849653, 0.0008742101, 0.0009001335, 0.0009095431, 
    0.0009270748, 0.0009585777, 0.0009814501, 0.001018818, 0.001020456, 
    0.001023444, 0.001004752, 0.0009552082, 0.0009354833, 0.0009911773, 
    0.001021726, 0.00102206, 0.001031295, 0.001315284, 0.001522008, 
    0.001540415, 0.001722439, 0.002065699, 0.002414457, 0.002817862, 
    0.00284795, 0.002890993, 0.002710366, 0.001936666, 0.002195843, 
    0.002328165, 0.002217014, 0.002013708, 0.00182062, 0.001777021, 
    0.001369707, 0.0009432076, 0.000691724, 0.0006145397, 0.0005666018, 
    0.0006265086, 0.0005630571, 0.0004425123, 0.0003748341, 0.0004602838, 
    0.0007488504, 0.0009390274, 0.0009709122, 0.001002654, 0.001127474, 
    0.001335709,
  0.001050196, 0.001014258, 0.0009499472, 0.001000636, 0.001014083, 
    0.00115235, 0.001236813, 0.00125994, 0.001389639, 0.001526237, 
    0.001621621, 0.001881735, 0.002115179, 0.002283932, 0.002275603, 
    0.002366583, 0.002423566, 0.002313034, 0.002257801, 0.002253065, 
    0.002228555, 0.002139132, 0.001954722, 0.001735283, 0.001643618, 
    0.001764878, 0.001659147, 0.001558216, 0.00140264, 0.001486786, 
    0.001523312, 0.001595681, 0.001703637, 0.00169011, 0.001589513, 
    0.001755722, 0.001854889, 0.001630378, 0.000910162, 0.0008607139, 
    0.00103352, 0.001010028, 0.0009661117, 0.0008985912, 0.0008998634, 
    0.0008877832, 0.0008611442, 0.0008443757, 0.0008390509, 0.0008200095, 
    0.00082384, 0.0008551199, 0.0009059827, 0.0009641727, 0.001009472, 
    0.001015623, 0.0009961845, 0.0009743292, 0.0009781756, 0.001008248, 
    0.001004418, 0.001000618, 0.001055948, 0.001148343, 0.001285719, 
    0.001320132, 0.001600766, 0.001966485, 0.002206158, 0.002161956, 
    0.002233593, 0.00230461, 0.002341994, 0.002312397, 0.002325734, 
    0.002222927, 0.00197289, 0.001784205, 0.001737396, 0.001636657, 
    0.001246397, 0.001226354, 0.0007305848, 0.0007433798, 0.0006817738, 
    0.0005470039, 0.00028317, 1.591817e-005, -7.814541e-005, 3.04142e-005, 
    0.0003520092, 0.000675479, 0.0008383514, 0.0008707922, 0.000875337, 
    0.0009131664,
  0.0008933935, 0.0007970734, 0.0007954836, 0.0008754656, 0.001048303, 
    0.001208124, 0.001352383, 0.001399478, 0.001475024, 0.001549411, 
    0.00185767, 0.002032653, 0.002182777, 0.002324334, 0.002286681, 
    0.002226949, 0.002215743, 0.002164515, 0.002099776, 0.001973526, 
    0.001958982, 0.001947729, 0.001775941, 0.001815119, 0.00162677, 
    0.001530433, 0.001423796, 0.001398842, 0.001472736, 0.001412272, 
    0.001184583, 0.001157022, 0.001277661, 0.001414672, 0.00135208, 
    0.001263896, 0.001346294, 0.001383376, 0.000867533, 0.0008170516, 
    0.001067026, 0.001147023, 0.001286261, 0.0009236885, 0.0008971291, 
    0.0008780714, 0.0008714749, 0.0008497792, 0.0008447571, 0.0008595865, 
    0.0008866391, 0.0009244685, 0.0009778584, 0.001044329, 0.00109551, 
    0.001091345, 0.00104638, 0.001007136, 0.0009858687, 0.0009702127, 
    0.0009212727, 0.0009774286, 0.001066089, 0.001307463, 0.001387143, 
    0.001517542, 0.001674883, 0.001784603, 0.001958886, 0.002183461, 
    0.00232443, 0.002423865, 0.002535669, 0.002554727, 0.002344188, 
    0.001036365, 0.001610255, 0.001598048, 0.001615389, 0.001538077, 
    0.001316873, 0.0006449139, 0.0005413764, 0.0005223025, 0.0004940578, 
    0.0004814225, 0.0003088554, 1.211884e-005, -0.0001789969, -0.0001137815, 
    0.0001761992, 0.0004603937, 0.0006210725, 0.0006980342, 0.0008332971, 
    0.0009156307,
  0.0005201581, 0.0006305613, 0.0007383106, 0.001085622, 0.00122896, 
    0.001340159, 0.001268028, 0.001562811, 0.001721772, 0.001833733, 
    0.00198346, 0.002114272, 0.00213848, 0.002297298, 0.002246833, 
    0.00213573, 0.00196572, 0.00200371, 0.002053508, 0.001944709, 
    0.001733819, 0.001633668, 0.00162189, 0.001534597, 0.001424431, 
    0.001389353, 0.001311518, 0.001401336, 0.001443108, 0.001309864, 
    0.00112741, 0.0009874906, 0.00100712, 0.001089485, 0.001152253, 
    0.00109044, 0.001033569, 0.001034729, 0.0007415842, 0.0006522411, 
    0.0007164069, 0.0007933211, 0.001037145, 0.0009941338, 0.0007758527, 
    0.0008506211, 0.0009038677, 0.0009724367, 0.001072462, 0.001145307, 
    0.00120879, 0.00116891, 0.001107144, 0.001124518, 0.001201653, 
    0.0009879987, 0.0009588478, 0.0009553512, 0.0009759027, 0.0009747264, 
    0.001018277, 0.001147183, 0.001270652, 0.001352175, 0.001396235, 
    0.001560394, 0.001666744, 0.001681495, 0.00189383, 0.002035658, 
    0.001970554, 0.00169731, 0.0007812097, 0.000516359, 0.0003900609, 
    0.000449125, 0.001188873, 0.001323485, 0.001208265, 0.001043072, 
    0.0004347244, 0.0004241222, 0.0003103646, 0.0001478745, 0.0001291987, 
    0.0003248286, 0.0003891224, 0.0002845041, 0.0001726858, 0.0001938739, 
    0.0002816441, 0.0003723064, 0.0004699626, 0.0005351142, 0.0006040335, 
    0.0006528613,
  0.0003236691, 0.0004359805, 0.0009022634, 0.001224128, 0.001419346, 
    0.001032694, 0.001384679, 0.001595871, 0.001717432, 0.001853092, 
    0.001985827, 0.002056257, 0.00208474, 0.002022401, 0.001939273, 
    0.001889475, 0.001783999, 0.001736791, 0.001661833, 0.001545295, 
    0.001439929, 0.001319909, 0.001229978, 0.001210491, 0.001198618, 
    0.001201431, 0.001122912, 0.001067169, 0.001056075, 0.001062544, 
    0.001057331, 0.001096463, 0.001129589, 0.00113814, 0.001096892, 
    0.00104301, 0.001040738, 0.000940585, 0.0008622566, 0.0007805573, 
    0.0007734857, 0.0008129836, 0.0009031375, 0.0009674625, 0.0009982022, 
    0.001002256, 0.001032773, 0.0008017616, 0.0008401945, 0.0008993852, 
    0.0009480701, 0.0009827842, 0.001255282, 0.001322563, 0.001345833, 
    0.001294939, 0.001145657, 0.00104053, 0.000971531, 0.0009062202, 
    0.0009538406, 0.001024826, 0.001156656, 0.001348647, 0.001449132, 
    0.001535407, 0.001617932, 0.001578816, 0.001656954, 0.00159851, 
    0.001356372, 0.0006630812, 0.0003914433, 0.0001986425, 0.0001639447, 
    0.0002849975, 0.0007854369, 0.0008771964, 0.0004782917, 0.0003157696, 
    0.0002078773, 0.0002538282, 0.0002094184, 0.0001072325, 0.0001171825, 
    8.822232e-005, 0.0001725587, 0.000307186, 0.0004158258, 0.0004642406, 
    0.0004536235, 0.000316882, 0.0001446963, 0.0001552659, 0.0002849498, 
    0.0003259261,
  0.0001811101, 0.0002834238, 0.000442815, 0.0009399974, 0.00112919, 
    0.001208027, 0.000800984, 0.00134027, 0.00141561, 0.00152115, 
    0.001569184, 0.001624306, 0.001625626, 0.001655587, 0.00169135, 
    0.001635258, 0.001525458, 0.001362412, 0.00118905, 0.0010789, 
    0.001056933, 0.001018246, 0.0009723422, 0.0009431923, 0.0009538569, 
    0.0009528715, 0.0009319065, 0.0008686939, 0.0007350841, 0.0006740647, 
    0.000710798, 0.0008130791, 0.0008935528, 0.0009013731, 0.000932558, 
    0.0009247861, 0.0009088754, 0.0009863772, 0.001011188, 0.0009703077, 
    0.0009251833, 0.0009315256, 0.0009888881, 0.0011046, 0.00119992, 
    0.001213843, 0.001086528, 0.0009657773, 0.001009884, 0.0007317453, 
    0.0006733327, 0.0004331665, 0.0008902946, 0.001062211, 0.001128411, 
    0.001077898, 0.0009573703, 0.0008708872, 0.000850352, 0.0008806633, 
    0.0009463555, 0.001064038, 0.001178432, 0.001308211, 0.001393104, 
    0.001412749, 0.001396331, 0.001334342, 0.001272083, 0.001168752, 
    0.001127044, 0.001109019, 0.001045011, 0.0009630434, 0.0005095876, 
    0.0004668473, 0.0004400965, 0.0007102725, 0.000624489, 0.0005282641, 
    0.0003155153, 0.0003147202, 0.0003803647, 0.0003121453, 0.00028193, 
    0.0002331177, 0.0001530724, 0.0001187716, 0.0001905994, 0.0003833049, 
    0.0004964899, 0.0005572708, 0.000350514, 8.996995e-005, -9.370968e-006, 
    2.480252e-005,
  0.0001790118, 0.00018537, 0.0002183835, 0.0002172701, 0.0002359147, 
    0.0008748774, 0.001035063, 0.001126186, 0.001138138, 0.001065023, 
    0.0009888876, 0.0006438803, 0.0006085471, 0.0006103751, 0.001071381, 
    0.001173535, 0.001226067, 0.001211476, 0.001154605, 0.001123865, 
    0.001083811, 0.00106043, 0.0009951834, 0.000909606, 0.0008507967, 
    0.001005434, 0.0008320878, 0.0006465344, 0.0005356702, 0.0004536235, 
    0.0004216908, 0.0004040156, 0.0004534163, 0.0005160253, 0.000558591, 
    0.0006115832, 0.0006365855, 0.0006226934, 0.0006954432, 0.0007419037, 
    0.0008091531, 0.0009091459, 0.0008720327, 0.000926137, 0.001004894, 
    0.001118985, 0.001145672, 0.00109233, 0.0009220042, 0.0005037701, 
    0.0003706531, 0.0002884148, 0.0002865391, 0.0006319922, 0.0007689083, 
    0.0008256044, 0.0008209306, 0.0007358477, 0.0006808206, 0.0007495964, 
    0.0007158993, 0.0008221706, 0.0008546435, 0.0009474992, 0.001010299, 
    0.001048812, 0.001069347, 0.00100669, 0.0009657778, 0.0005839264, 
    0.0008854456, 0.0009172028, 0.0009758228, 0.0006416559, 0.000781782, 
    0.0004892107, 0.0007099702, 0.0007138008, 0.0007107493, 0.0005508021, 
    0.0004983502, 0.0004021088, 0.0005025303, 0.0004935029, 0.0005063456, 
    0.0004821701, 0.000422772, 0.0003378633, 0.000264748, 0.0002455632, 
    0.0002211968, 0.0002246457, 0.0002612029, 0.0002603924, 0.0002604718, 
    0.0002227537,
  0.0004467405, 0.0004348983, 0.00037194, 0.0003474304, 0.000324876, 
    0.000444483, 0.0006379201, 0.000733987, 0.0006840145, 0.0005898073, 
    0.0004811364, 0.0004164772, 0.0003657101, 0.0003086643, 0.0003339369, 
    0.0006537039, 0.000489481, 0.0005126393, 0.0005067107, 0.000756335, 
    0.0007646787, 0.0007967069, 0.0007497701, 0.0007362911, 0.0007227017, 
    0.0006708694, 0.0006181309, 0.0005374504, 0.000471917, 0.000395163, 
    0.0003912845, 0.00035762, 0.000332729, 0.0002927538, 0.0002883668, 
    0.0003322517, 0.0003579534, 0.0003795065, 0.0004785922, 0.0005155634, 
    0.0004296058, 0.0004138066, 0.0004050967, 0.0004126467, 0.0004316089, 
    0.0004476306, 0.0004403354, 0.0004066864, 0.0003522793, 0.0002863486, 
    0.0002343415, 0.0002070665, 0.0002121846, 0.000239555, 0.0002670847, 
    0.0002796573, 0.0002744913, 0.0002568325, 0.0002372502, 0.0002295892, 
    0.0002355336, 0.0002490275, 0.0002941047, 0.000686605, 0.0008200239, 
    0.0008873059, 0.0009107501, 0.0008715703, 0.0008322946, 0.0004952354, 
    0.0007732308, 0.0007969455, 0.000552837, 0.0008208826, 0.0007340347, 
    0.0006762582, 0.0005894895, 0.0003738799, 0.000377981, 0.000362881, 
    0.0003267366, 0.0005559039, 0.0004408283, 0.0004776878, 0.0005057736, 
    0.000521859, 0.0005227808, 0.0004930579, 0.0004280012, 0.0003522479, 
    0.0003781714, 0.000208592, 0.0001536764, 0.0001549004, 0.0002737441, 
    0.0003664407,
  0.0002753655, 0.0003611164, 0.0004068131, 0.0004818672, 0.0005153732, 
    0.0004177648, 0.000384704, 0.0003492909, 0.0003101267, 0.0002936916, 
    0.0002911487, 0.000295599, 0.0003040233, 0.0003183761, 0.0003330945, 
    0.0003439505, 0.0003525175, 0.0003604013, 0.0003706531, 0.0003795545, 
    0.000377059, 0.0003874858, 0.0003989774, 0.0003962279, 0.0003817321, 
    0.0007029609, 0.0007285036, 0.0005418696, 0.0005227006, 0.0005040877, 
    0.0004358999, 0.0002923093, 0.0002413832, 0.000199517, 0.000183336, 
    0.0001897733, 0.0002046507, 0.000232164, 0.0002552271, 0.0002662421, 
    0.0002621729, 0.0002611396, 0.0002592164, 0.0002578972, 0.0002635557, 
    0.0002763984, 0.0002915619, 0.0003071227, 0.0003220476, 0.0003340957, 
    0.0003482101, 0.0003635804, 0.000379316, 0.0003910619, 0.0003949562, 
    0.0003888204, 0.0003729262, 0.0003470019, 0.0003176134, 0.0002913871, 
    0.0002703904, 0.0002562918, 0.0002542415, 0.0002482014, 0.0002366938, 
    0.0006983201, 0.0007177908, 0.0007313648, 0.000738692, 0.000767811, 
    0.0007465282, 0.000696158, 0.0007132129, 0.0007370231, 0.0006480613, 
    0.0003797766, 0.0003634212, 0.0003524544, 0.0004595998, 0.0004949966, 
    0.0005244655, 0.000533128, 0.0005255624, 0.000511877, 0.0005083483, 
    0.0005203011, 0.0005368473, 0.0005481484, 0.000534336, 0.0004945202, 
    0.0004320543, 0.0005215721, 0.0002703904, 0.0002432745, 0.0001810468, 
    0.000163547,
  0.00028913, 0.0002886213, 0.0002738873, 0.0002637627, 0.000360878, 
    0.0003665369, 0.0003715435, 0.0003439663, 0.0003484965, 0.0003490208, 
    0.0003532809, 0.0003608784, 0.0003724017, 0.0003799833, 0.0003850379, 
    0.0003850218, 0.0003764706, 0.0003630875, 0.0003450788, 0.0003234781, 
    0.0003006377, 0.0002786079, 0.0002572613, 0.0002409536, 0.0002146321, 
    0.0003099041, 0.0003197112, 0.0002983648, 0.0003044682, 0.0003062165, 
    0.0002956945, 0.0002765891, 0.000255672, 0.0002381401, 0.0002239624, 
    0.0002141397, 0.0002121369, 0.0002195439, 0.0002338011, 0.0002558467, 
    0.0002773998, 0.0003019886, 0.0003200448, 0.0003352242, 0.0003475107, 
    0.0003546316, 0.000352009, 0.0003466208, 0.0003368296, 0.0003294225, 
    0.0003208555, 0.0003117479, 0.0003075679, 0.0003062324, 0.0003102697, 
    0.0003183284, 0.0003264982, 0.0003316479, 0.0003310121, 0.0003275154, 
    0.0003195524, 0.0003061057, 0.0002981902, 0.0002986987, 0.0003058515, 
    0.0003230174, 0.0003448564, 0.0003735938, 0.0004046836, 0.0004306715, 
    0.000441893, 0.0007010696, 0.0007632489, 0.0005469404, 0.0005415361, 
    0.0005261505, 0.0005072518, 0.0004944883, 0.0004810255, 0.0004726175, 
    0.0004608238, 0.0004459941, 0.0004334374, 0.0004263644, 0.0004270637, 
    0.0004256967, 0.0004257603, 0.0004206898, 0.0004156512, 0.000404668, 
    0.0004012031, 0.0003886141, 0.0003272134, 0.0003103493, 0.0003043411, 
    0.0002967275,
  0.0003476699, 0.0003442683, 0.0003450315, 0.0003466208, 0.0003506104, 
    0.0003575562, 0.0003684759, 0.0003807626, 0.0003941774, 0.0004069407, 
    0.0004176379, 0.0004268566, 0.000435408, 0.0004386345, 0.0004403193, 
    0.0004385074, 0.0004322608, 0.0004240274, 0.0004117887, 0.000399089, 
    0.0003854036, 0.0003751358, 0.0003628333, 0.000356046, 0.000350022, 
    0.0003432669, 0.0003393092, 0.0003349222, 0.0003305988, 0.0003251312, 
    0.0003183442, 0.000310238, 0.0003001448, 0.0002897659, 0.0002817712, 
    0.0002743483, 0.0002676088, 0.0002666553, 0.0002714237, 0.0002790689, 
    0.0002881289, 0.0002975543, 0.0003095069, 0.0003159125, 0.0003215233, 
    0.0003254176, 0.000329566, 0.0003326654, 0.0003341117, 0.0003332854, 
    0.0003322521, 0.0003316798, 0.0003299157, 0.0003314731, 0.0003350335, 
    0.000338403, 0.0003410734, 0.0003414231, 0.0003408827, 0.0003405649, 
    0.0003385302, 0.0003341595, 0.000332427, 0.000327579, 0.0003228583, 
    0.0003229536, 0.0003256716, 0.0003298838, 0.0003385462, 0.0003456988, 
    0.0003548542, 0.0003653921, 0.000382209, 0.0004004398, 0.0004209599, 
    0.0004367433, 0.0004567544, 0.0004733959, 0.0004878601, 0.0005022287, 
    0.0005096039, 0.0005174559, 0.0005212387, 0.0005226214, 0.0005178372, 
    0.0005065203, 0.0004930415, 0.0004778784, 0.0004533369, 0.0004349311, 
    0.0004152376, 0.0003952105, 0.0003813819, 0.0003677923, 0.0003574765, 
    0.000350849,
  0.0003987865, 0.0003963388, 0.0003963229, 0.0003961322, 0.0003961003, 
    0.0003973085, 0.0003987867, 0.0004005828, 0.0004032848, 0.0004077828, 
    0.0004117568, 0.0004143792, 0.0004171131, 0.0004203238, 0.0004233439, 
    0.0004237252, 0.0004244724, 0.0004232961, 0.0004231371, 0.0004226284, 
    0.0004209755, 0.0004180826, 0.0004157142, 0.0004126152, 0.0004097542, 
    0.0004056692, 0.0004009644, 0.0003976743, 0.0003937643, 0.0003888367, 
    0.0003848316, 0.0003803652, 0.000377472, 0.0003769156, 0.0003754376, 
    0.0003741819, 0.0003745791, 0.0003748811, 0.0003775514, 0.0003787754, 
    0.000381398, 0.0003851491, 0.0003880896, 0.0003915862, 0.0003958938, 
    0.0004015204, 0.0004034119, 0.0004045723, 0.0004098015, 0.00041306, 
    0.0004148402, 0.0004183687, 0.0004199264, 0.0004215317, 0.0004227397, 
    0.0004223105, 0.0004211662, 0.0004204826, 0.0004184325, 0.0004157939, 
    0.0004139182, 0.0004122653, 0.0004126625, 0.0004111684, 0.0004105009, 
    0.0004094518, 0.0004063046, 0.000404143, 0.0004035232, 0.0004024263, 
    0.0004033167, 0.0004063365, 0.0004078466, 0.0004115817, 0.0004155077, 
    0.000419402, 0.0004237252, 0.0004276987, 0.0004309255, 0.0004341363, 
    0.0004371244, 0.0004410185, 0.0004416066, 0.0004417815, 0.0004409549, 
    0.0004390315, 0.0004360275, 0.0004327216, 0.0004285572, 0.0004239795, 
    0.0004218337, 0.000417558, 0.0004112481, 0.0004066704, 0.0004027763, 
    0.0004001854,
  6.982305e-006, 6.712098e-006, 6.267053e-006, 5.822005e-006, 5.45643e-006, 
    5.043164e-006, 4.693482e-006, 4.327909e-006, 4.010019e-006, 
    3.692126e-006, 3.39013e-006, 3.15171e-006, 3.008658e-006, 2.738449e-006, 
    2.627188e-006, 2.436453e-006, 2.372874e-006, 2.229826e-006, 
    2.150353e-006, 2.134457e-006, 2.166245e-006, 2.134456e-006, 
    2.229824e-006, 2.341086e-006, 2.420558e-006, 2.515928e-006, 
    2.674872e-006, 2.833818e-006, 3.040447e-006, 3.231182e-006, 
    3.453704e-006, 3.692125e-006, 3.962333e-006, 4.312014e-006, 
    4.693482e-006, 5.02727e-006, 5.424634e-006, 5.869686e-006, 6.29884e-006, 
    6.871045e-006, 7.31609e-006, 7.920084e-006, 8.428711e-006, 9.000914e-006, 
    9.58901e-006, 1.014532e-005, 1.066984e-005, 1.111489e-005, 1.168709e-005, 
    1.19732e-005, 1.245003e-005, 1.262487e-005, 1.264076e-005, 1.27997e-005, 
    1.270434e-005, 1.283149e-005, 1.25295e-005, 1.246592e-005, 1.205267e-005, 
    1.198909e-005, 1.178246e-005, 1.144868e-005, 1.140099e-005, 
    1.105131e-005, 1.084468e-005, 1.059037e-005, 1.036785e-005, 
    1.009764e-005, 9.700274e-006, 9.477753e-006, 9.191648e-006, 
    8.937335e-006, 8.539973e-006, 8.094925e-006, 8.126714e-006, 
    7.999555e-006, 7.777027e-006, 7.681658e-006, 7.729341e-006, 
    7.792914e-006, 7.840605e-006, 7.951865e-006, 8.063129e-006, 
    8.126703e-006, 8.28565e-006, 8.444596e-006, 8.539966e-006, 8.555857e-006, 
    8.667121e-006, 8.619434e-006, 8.539966e-006, 8.365128e-006, 
    8.206185e-006, 7.96777e-006, 7.697559e-006, 7.411461e-006,
  1.200499e-005, 1.033606e-005, 8.826079e-006, 7.411458e-006, 6.346518e-006, 
    5.281581e-006, 4.343802e-006, 3.612653e-006, 3.024551e-006, 
    2.515926e-006, 2.150351e-006, 1.896038e-006, 1.62583e-006, 1.482781e-006, 
    1.466885e-006, 1.466884e-006, 1.419201e-006, 1.387411e-006, 
    1.323833e-006, 1.435094e-006, 1.371517e-006, 1.371516e-006, 
    1.450989e-006, 1.562251e-006, 1.689408e-006, 1.927826e-006, 
    2.150351e-006, 2.293402e-006, 2.674872e-006, 2.94508e-006, 3.310654e-006, 
    3.803385e-006, 4.423275e-006, 5.186214e-006, 6.012733e-006, 
    7.173041e-006, 8.539975e-006, 1.035195e-005, 1.273613e-005, 
    1.567663e-005, 1.893502e-005, 2.267024e-005, 2.646905e-005, 
    3.076057e-005, 3.433685e-005, 3.697535e-005, 4.071058e-005, 
    4.334908e-005, 4.549485e-005, 4.698894e-005, 4.848303e-005, 
    5.113742e-005, 5.115333e-005, 5.310835e-005, 5.050164e-005, 
    5.511106e-005, 5.44276e-005, 5.32514e-005, 5.191626e-005, 5.002481e-005, 
    4.814925e-005, 4.627368e-005, 4.404844e-005, 4.217289e-005, 
    4.044038e-005, 3.916882e-005, 3.781777e-005, 3.65462e-005, 3.524285e-005, 
    3.354214e-005, 3.157122e-005, 2.926649e-005, 2.656441e-005, 
    2.392591e-005, 2.154172e-005, 1.979333e-005, 1.866481e-005, 
    1.812439e-005, 1.710714e-005, 1.699587e-005, 1.740913e-005, 
    1.651905e-005, 1.834692e-005, 1.836281e-005, 2.022248e-005, 
    2.122384e-005, 2.25113e-005, 2.324245e-005, 2.348087e-005, 2.327423e-005, 
    2.25113e-005, 2.119204e-005, 1.941185e-005, 1.761576e-005, 1.559715e-005, 
    1.368982e-005,
  7.02999e-006, 5.822005e-006, 4.979591e-006, 4.423277e-006, 4.105383e-006, 
    3.994122e-006, 4.089489e-006, 4.200751e-006, 4.343801e-006, 
    4.439168e-006, 4.423275e-006, 4.502746e-006, 4.55043e-006, 4.788851e-006, 
    5.233898e-006, 5.567684e-006, 6.04452e-006, 6.346516e-006, 6.298833e-006, 
    5.774313e-006, 4.916008e-006, 3.644441e-006, 2.420559e-006, 
    1.435094e-006, 8.469951e-007, 7.675226e-007, 9.900464e-007, 
    1.371517e-006, 1.975511e-006, 2.643083e-006, 3.167605e-006, 
    3.549074e-006, 3.787494e-006, 3.96233e-006, 4.455066e-006, 5.20211e-006, 
    6.569047e-006, 8.778392e-006, 1.190961e-005, 1.608989e-005, 
    2.092183e-005, 2.522928e-005, 3.012481e-005, 3.341498e-005, 
    3.486139e-005, 3.621243e-005, 3.643495e-005, 3.668925e-005, 
    3.761114e-005, 4.048807e-005, 4.544718e-005, 5.264742e-005, 
    6.124638e-005, 7.054468e-005, 7.95728e-005, 8.661411e-005, 9.106456e-005, 
    9.236793e-005, 8.963404e-005, 8.462729e-005, 7.81423e-005, 7.07672e-005, 
    6.312193e-005, 5.655746e-005, 5.159837e-005, 4.870554e-005, 
    4.722735e-005, 4.695713e-005, 4.67505e-005, 4.617831e-005, 4.465243e-005, 
    4.209341e-005, 3.845355e-005, 3.500444e-005, 3.230235e-005, 
    3.066521e-005, 2.912344e-005, 2.987049e-005, 3.180962e-005, 
    3.419381e-005, 3.734093e-005, 4.102847e-005, 4.350803e-005, 
    4.533591e-005, 4.598759e-005, 4.592401e-005, 4.525644e-005, 4.44617e-005, 
    4.214111e-005, 3.83264e-005, 3.413023e-005, 2.824923e-005, 2.216161e-005, 
    1.672567e-005, 1.216393e-005, 9.032694e-006,
  1.198909e-005, 1.084469e-005, 9.875115e-006, 9.080384e-006, 8.539969e-006, 
    8.142603e-006, 8.222077e-006, 8.285652e-006, 8.174392e-006, 
    7.649874e-006, 6.664411e-006, 5.329266e-006, 4.0577e-006, 3.183498e-006, 
    2.77024e-006, 2.817926e-006, 3.119927e-006, 4.073599e-006, 5.647165e-006, 
    7.745231e-006, 9.000909e-006, 8.794286e-006, 7.220724e-006, 
    5.297481e-006, 3.406023e-006, 2.277507e-006, 1.784776e-006, 
    1.927827e-006, 2.341086e-006, 2.770238e-006, 3.040445e-006, 
    2.976869e-006, 2.722558e-006, 2.91329e-006, 3.390131e-006, 4.280224e-006, 
    5.85379e-006, 7.618093e-006, 9.541332e-006, 1.216393e-005, 1.553357e-005, 
    1.942775e-005, 2.511802e-005, 3.176194e-005, 3.786546e-005, 
    4.374645e-005, 6.846248e-005, 6.556967e-005, 7.156192e-005, 
    8.024036e-005, 9.416402e-005, 0.0001098202, 0.0001242206, 0.0001369522, 
    0.0001447246, 0.0001448836, 0.0001432464, 0.0001183396, 0.0001102175, 
    0.0001047338, 9.858265e-005, 9.441828e-005, 8.979299e-005, 8.332389e-005, 
    7.582165e-005, 6.779493e-005, 6.111922e-005, 5.744759e-005, 
    5.555613e-005, 5.460245e-005, 5.35375e-005, 5.128048e-005, 4.67982e-005, 
    4.061522e-005, 3.51316e-005, 3.130101e-005, 2.880556e-005, 2.858303e-005, 
    2.963208e-005, 3.300172e-005, 4.873733e-005, 5.436399e-005, 
    5.865553e-005, 6.277222e-005, 6.558557e-005, 6.970225e-005, 
    7.540842e-005, 8.182981e-005, 9.362359e-005, 7.413687e-005, 
    6.660284e-005, 5.536538e-005, 4.18709e-005, 2.977512e-005, 2.061986e-005, 
    1.478653e-005,
  3.695946e-005, 3.285867e-005, 2.851945e-005, 2.362392e-005, 2.036553e-005, 
    1.917344e-005, 2.081058e-005, 2.457759e-005, 2.905986e-005, 
    3.177784e-005, 3.123742e-005, 2.735914e-005, 2.19391e-005, 1.658262e-005, 
    1.305403e-005, 1.094005e-005, 1.033606e-005, 1.057448e-005, 
    1.070162e-005, 9.763848e-006, 1.178246e-005, 1.448453e-005, 
    1.448453e-005, 1.178245e-005, 8.015457e-006, 4.979594e-006, 
    3.167612e-006, 2.531828e-006, 2.658986e-006, 3.07224e-006, 3.564975e-006, 
    4.232548e-006, 4.995487e-006, 6.235259e-006, 8.55586e-006, 1.256129e-005, 
    1.732966e-005, 2.225698e-005, 2.491138e-005, 2.529285e-005, 
    2.500675e-005, 2.767703e-005, 3.358982e-005, 4.15371e-005, 5.131226e-005, 
    6.177089e-005, 8.569221e-005, 0.0001035418, 0.0001264777, 0.0001507964, 
    0.0001695361, 0.0001830941, 0.0001917249, 0.0001972721, 0.0001951581, 
    0.000184636, 0.000166707, 0.0001512574, 0.0001438187, 0.0001462824, 
    0.000153419, 0.0001596656, 0.0001599677, 0.0001571225, 0.000152672, 
    0.0001501766, 0.0001519091, 0.0001604763, 0.000168805, 0.0001710621, 
    0.0001387166, 0.0001303243, 0.0001172907, 0.0001046227, 9.594433e-005, 
    9.479991e-005, 6.704789e-005, 6.207291e-005, 6.011783e-005, 6.30742e-005, 
    7.256333e-005, 9.127118e-005, 0.0001103129, 0.0001241094, 0.0001321679, 
    0.0001376039, 0.0001414662, 0.0001445339, 0.0001456465, 0.000138192, 
    0.0001274631, 7.795155e-005, 5.992712e-005, 4.94367e-005, 4.230004e-005, 
    4.031323e-005,
  0.0001932508, 0.0001860664, 0.0001023338, 8.416634e-005, 7.229309e-005, 
    6.78108e-005, 6.863735e-005, 7.423222e-005, 8.502467e-005, 9.448195e-005, 
    9.66595e-005, 8.853739e-005, 7.216593e-005, 5.264741e-005, 3.811978e-005, 
    2.953671e-005, 2.573791e-005, 2.376697e-005, 2.478423e-005, 
    2.616704e-005, 2.967977e-005, 3.363751e-005, 3.366929e-005, 
    2.942544e-005, 2.354445e-005, 1.950723e-005, 1.728199e-005, 1.64237e-005, 
    1.49932e-005, 1.519981e-005, 1.659853e-005, 1.77906e-005, 1.980925e-005, 
    2.440278e-005, 3.147587e-005, 3.964567e-005, 4.872147e-005, 
    5.658927e-005, 6.425046e-005, 7.380312e-005, 8.710688e-005, 0.0001028425, 
    0.0001189437, 0.0001301811, 0.0001585211, 0.0001687095, 0.000180996, 
    0.0001987981, 0.0002139775, 0.0002294905, 0.0002489295, 0.0002652691, 
    0.0002759662, 0.0002758548, 0.0002633458, 0.0002431915, 0.0002248652, 
    0.0002182848, 0.0002283144, 0.0002420633, 0.000250376, 0.0002551127, 
    0.0002577194, 0.0002586094, 0.0002684959, 0.0002883959, 0.0003065474, 
    0.0003261453, 0.0003393379, 0.0003419604, 0.0003270673, 0.0003061975, 
    0.0002988703, 0.0002987908, 0.0003075328, 0.000313382, 0.0003101715, 
    0.0002911139, 0.00023499, 0.0002156463, 0.0002258825, 0.0002323197, 
    0.0002435572, 0.0002520767, 0.0002572424, 0.0002557165, 0.0002487865, 
    0.0002380418, 0.0002251037, 0.000205299, 0.0001889116, 0.0001803126, 
    0.0001782622, 0.0001837458, 0.000192154, 0.0001949038,
  0.0003770398, 0.0003704595, 0.0003489223, 0.0003287521, 0.0003201691, 
    0.0003233002, 0.0003279733, 0.0003254619, 0.0003195174, 0.0003142721, 
    0.0003084706, 0.0002986478, 0.0002820221, 0.0002518859, 0.0002111957, 
    0.0001702195, 0.0001442319, 0.0001355694, 0.0001427219, 0.0001567727, 
    0.0001603172, 0.0001525765, 0.0001336302, 0.0001132057, 0.0001050041, 
    0.0001086122, 0.0001146998, 0.0001125541, 9.890055e-005, 8.217955e-005, 
    7.084676e-005, 6.892352e-005, 6.364641e-005, 4.075823e-005, 
    4.902342e-005, 6.402784e-005, 8.815603e-005, 0.0001133487, 0.0001376357, 
    0.0001646087, 0.0001897381, 0.0002041229, 0.0002094316, 0.0002143588, 
    0.0002280601, 0.0002478331, 0.0002667952, 0.0002614545, 0.0002268204, 
    0.0001767843, 0.0001480469, 0.0001599836, 0.0001517821, 0.0001518298, 
    0.0001696476, 0.0001684873, 0.0001959054, 0.0001958419, 0.0002247859, 
    0.00027541, 0.0003015408, 0.0003521332, 0.0004164584, 0.0005036403, 
    0.0005831288, 0.0006688004, 0.0007521515, 0.0007717336, 0.0008162542, 
    0.0008371398, 0.0008624282, 0.0008988424, 0.0009132111, 0.000901735, 
    0.0008500301, 0.0007699218, 0.0006612669, 0.0005929357, 0.000541247, 
    0.0005001434, 0.0004515854, 0.0004303503, 0.0004186677, 0.0004108636, 
    0.0004098146, 0.0004134225, 0.0004178254, 0.0004132796, 0.0003967808, 
    0.0003731297, 0.0003488745, 0.0003242221, 0.0003063884, 0.0003083911, 
    0.0003294515, 0.0003572988,
  0.0006618868, 0.0007136869, 0.0007472879, 0.0007690478, 0.0008134573, 
    0.0008792608, 0.0009380708, 0.0009592102, 0.0009530907, 0.0009419172, 
    0.0009557612, 0.0009754704, 0.0009777275, 0.0009701933, 0.0009266263, 
    0.0008803735, 0.0007928103, 0.000719727, 0.000644784, 0.0005609242, 
    0.0004833426, 0.0004258998, 0.0004013586, 0.0003805367, 0.0003867674, 
    0.0003797102, 0.0003834772, 0.0003775008, 0.0003910112, 0.0003705549, 
    0.0003263681, 0.0003697763, 0.0003323599, 0.0002736454, 0.0002038365, 
    0.0002369608, 0.0003644512, 0.0004116739, 0.000414853, 0.0003926323, 
    0.0003927117, 0.0004046327, 0.000390264, 0.0003799647, 0.0003609385, 
    0.0002990768, 0.0001949673, 4.323805e-005, -7.603504e-005, -0.0001178377, 
    -0.0001347177, -0.0001559847, -0.0001717047, -0.0001698448, 
    -0.0001009421, -3.628246e-005, 2.548378e-005, 7.588509e-005, 
    0.0001665796, 0.0002864725, 0.000372939, 0.0004156639, 0.0004145191, 
    0.0004051095, 0.0004339265, 0.0004779224, 0.0005135739, 0.000541898, 
    0.000559716, 0.0005718435, 0.0005890415, 0.0006173973, 0.0006602171, 
    0.0007077262, 0.0007392927, 0.0007341271, 0.0007130825, 0.0006788142, 
    0.0006490755, 0.0006557989, 0.0006906714, 0.0006498698, 0.0006374565, 
    0.0006288259, 0.000624137, 0.0006384262, 0.0006508557, 0.0006282855, 
    0.0005958127, 0.000582382, 0.0005851952, 0.0005655974, 0.000537909, 
    0.0005307246, 0.0005448232, 0.0005991668,
  0.0007647878, 0.0007619106, 0.0007697624, 0.0007832572, 0.0008083864, 
    0.0008201802, 0.0008090544, 0.000749259, 0.0006968388, 0.0007022428, 
    0.0007054692, 0.0007110641, 0.0007251466, 0.0007442678, 0.0007901238, 
    0.0008263474, 0.0008619989, 0.0009038015, 0.0009414402, 0.0009112244, 
    0.0008169693, 0.0008002643, 0.0007958933, 0.0007668539, 0.000715276, 
    0.0006742999, 0.0006343885, 0.0006275061, 0.0006075108, 0.0005873251, 
    0.0005320278, 0.0004423349, 0.0003869578, 0.0003506704, 0.0003306274, 
    0.0003331548, 0.0003208206, 0.0003155277, 0.0003225531, 0.000365373, 
    0.0004236426, 0.0004811808, 0.0005604948, 0.000635454, 0.0006371385, 
    0.0006181765, 0.0005139709, 0.0002888883, 0.0001310715, 6.353529e-005, 
    4.031323e-005, 1.478614e-005, -2.638041e-005, -6.25567e-005, 
    -9.487034e-005, -0.0001175676, -8.827401e-005, -1.453888e-005, 
    9.071478e-005, 0.0001747494, 0.0002399809, 0.0002962318, 0.0003487633, 
    0.0003749095, 0.0003989742, 0.0004510127, 0.0005192487, 0.0005493369, 
    0.0005487008, 0.0005511802, 0.0005609395, 0.0005839071, 0.0006204972, 
    0.0006358034, 0.0006310979, 0.0005936984, 0.000534412, 0.0005398002, 
    0.0005674884, 0.0005677589, 0.0005788852, 0.0006329268, 0.0006099432, 
    0.0006494883, 0.0007290728, 0.0007834481, 0.0008446102, 0.0008696122, 
    0.0008406523, 0.0008632862, 0.0008988106, 0.0008656069, 0.0008168903, 
    0.0007566339, 0.0007266885, 0.0007444904,
  0.000582048, 0.000603792, 0.0006247726, 0.0006314006, 0.0006138689, 
    0.0006045073, 0.0006065096, 0.0005829537, 0.0005507513, 0.0005404835, 
    0.0005306767, 0.0005232061, 0.0005308671, 0.0005637533, 0.0005972749, 
    0.0006280467, 0.0006896541, 0.0007717179, 0.0008085612, 0.0007663611, 
    0.0006887324, 0.0006259808, 0.0005801723, 0.0005653109, 0.0005638804, 
    0.0005969729, 0.0006401106, 0.0006485984, 0.0006440049, 0.0006501242, 
    0.0006414298, 0.0005968611, 0.0005766274, 0.0005954306, 0.0006190499, 
    0.0006010893, 0.00054282, 0.0004682743, 0.0004345141, 0.0004619327, 
    0.0005573644, 0.0006648912, 0.0007889327, 0.0008137119, 0.0007965458, 
    0.000768492, 0.000718201, 0.0005722102, 0.000377994, 0.0002472927, 
    0.0001872745, 0.0001501292, 0.0001079924, 8.534314e-005, 0.0001112353, 
    0.0001373501, 0.0001713005, 0.0002112119, 0.0002514096, 0.0002846448, 
    0.0003459346, 0.0004061111, 0.0004311451, 0.0004241834, 0.0004302394, 
    0.0004687994, 0.0005009701, 0.0005297712, 0.0005503548, 0.000568077, 
    0.0005926182, 0.0006216099, 0.0006297166, 0.0006025368, 0.000552326, 
    0.000520187, 0.0005500684, 0.0005882627, 0.0005894704, 0.0005605752, 
    0.0005763746, 0.0006328318, 0.000763071, 0.0006748089, 0.0006275063, 
    0.0006382032, 0.0006746177, 0.0006832485, 0.0006760962, 0.0006656372, 
    0.0006331329, 0.0005959081, 0.0005677906, 0.0005506244, 0.0005541372, 
    0.0005662807,
  0.0005968774, 0.0006031715, 0.0006374882, 0.0006691816, 0.000666416, 
    0.0006583417, 0.0006780992, 0.0006884143, 0.0006906711, 0.0007042296, 
    0.0006935964, 0.000681214, 0.0006943117, 0.0006966477, 0.0006999536, 
    0.0007334757, 0.00081786, 0.0009008457, 0.000852796, 0.0008081638, 
    0.0008261723, 0.0009135134, 0.0009553642, 0.000942776, 0.0009145788, 
    0.0009193476, 0.0009613731, 0.0009782366, 0.0009510415, 0.0009063934, 
    0.0008438644, 0.0007753745, 0.0007403903, 0.0007555694, 0.000798326, 
    0.0007988503, 0.0007195203, 0.0006325771, 0.000589042, 0.0006496636, 
    0.0008009486, 0.000908793, 0.000919681, 0.000922638, 0.0009589409, 
    0.0009532347, 0.000895171, 0.0007366389, 0.0005375277, 0.0004458795, 
    0.0004290789, 0.0004732502, 0.0004859655, 0.0004770965, 0.0004684338, 
    0.0004551937, 0.0004432253, 0.0004436225, 0.0004440518, 0.0004434637, 
    0.000484535, 0.0005346984, 0.0005254797, 0.0005041808, 0.0005076141, 
    0.0004836768, 0.000460153, 0.0004911949, 0.0005318057, 0.0005379724, 
    0.000541247, 0.0005733538, 0.0005945736, 0.0005675843, 0.0005319011, 
    0.0005945577, 0.000632911, 0.000615204, 0.0006396822, 0.0006481381, 
    0.0006067641, 0.0005634525, 0.0006348025, 0.0005919663, 0.0005777087, 
    0.0006196229, 0.0006748408, 0.0006907505, 0.0006739974, 0.0006415891, 
    0.0005997701, 0.0005812533, 0.000591696, 0.0005891055, 0.0005741958, 
    0.0005862759,
  0.0007167868, 0.0007616733, 0.0008036345, 0.00083412, 0.0008510007, 
    0.0008958071, 0.0009803185, 0.001062859, 0.001104535, 0.001136975, 
    0.001156574, 0.001168574, 0.001153442, 0.001078754, 0.001005925, 
    0.0009848801, 0.001044405, 0.001169257, 0.001225731, 0.001372931, 
    0.001627196, 0.001755784, 0.001675977, 0.00151568, 0.001406596, 
    0.001342652, 0.001298544, 0.001237382, 0.001169417, 0.001071856, 
    0.0009646947, 0.0009047878, 0.0008658781, 0.0008307667, 0.0007981188, 
    0.0007436485, 0.0006729653, 0.0006515565, 0.0006705178, 0.0007413123, 
    0.0009672539, 0.001099084, 0.00107203, 0.001076831, 0.00116859, 
    0.001110543, 0.001032692, 0.0009479257, 0.0008542594, 0.0007567937, 
    0.0007788721, 0.0008880994, 0.0009486419, 0.000895808, 0.0008365852, 
    0.0007800162, 0.0007094918, 0.0006657182, 0.0006345012, 0.0006116442, 
    0.0006247256, 0.0006345958, 0.0006311946, 0.0006332602, 0.0006232471, 
    0.0005961629, 0.0005867532, 0.0005919668, 0.0005907905, 0.0005836221, 
    0.0005786149, 0.0006000884, 0.0006147595, 0.0006195279, 0.0006103893, 
    0.0006202916, 0.0006185742, 0.0005418342, 0.0005755306, 0.0006847433, 
    0.0006795139, 0.0006399998, 0.0006256471, 0.0005902979, 0.0005887402, 
    0.0006388398, 0.0007358445, 0.0007965295, 0.0007864367, 0.0007442525, 
    0.0006768592, 0.0006342465, 0.0006397143, 0.0006414945, 0.0006428934, 
    0.0006774957,
  0.0009439206, 0.0009878217, 0.001010853, 0.001006435, 0.001045725, 
    0.001187886, 0.001451481, 0.001702758, 0.001876486, 0.002028264, 
    0.002121041, 0.002087836, 0.001886739, 0.001663945, 0.001543193, 
    0.001517746, 0.001525979, 0.001579639, 0.001648129, 0.001692967, 
    0.001693191, 0.001626592, 0.001454581, 0.001296462, 0.001227749, 
    0.001166699, 0.001082791, 0.0009870259, 0.0009249575, 0.0008796742, 
    0.0008770199, 0.0008862545, 0.000856325, 0.0007749922, 0.0007344456, 
    0.0007395796, 0.0007664091, 0.0008385228, 0.0008878759, 0.0009482438, 
    0.001116789, 0.001189237, 0.001222265, 0.001286654, 0.001400889, 
    0.001526551, 0.001294857, 0.001239003, 0.001246632, 0.001293425, 
    0.001385089, 0.001416752, 0.001340855, 0.001214653, 0.001140997, 
    0.001033104, 0.0008672602, 0.0007813503, 0.0007674904, 0.0007604808, 
    0.0007706373, 0.0007660757, 0.0007715272, 0.0007811277, 0.000747479, 
    0.0007480192, 0.0007507852, 0.0007137028, 0.0006833607, 0.0006829789, 
    0.0006929287, 0.0006974745, 0.0007182648, 0.0007358915, 0.0006909897, 
    0.0006128838, 0.0005934285, 0.0005363361, 0.0005453159, 0.0007026098, 
    0.0007611653, 0.000766919, 0.0007733088, 0.000835822, 0.0008890047, 
    0.0009110034, 0.0009415052, 0.0009508035, 0.0009148815, 0.0008935356, 
    0.0008700429, 0.0008507469, 0.0008584876, 0.0008580745, 0.0008739531, 
    0.0009127362,
  0.001059489, 0.001047458, 0.001015445, 0.00101961, 0.001153284, 
    0.001437493, 0.001604418, 0.001713946, 0.001801653, 0.001873687, 
    0.001752475, 0.00155241, 0.00134977, 0.001212345, 0.001175359, 
    0.001175168, 0.001183323, 0.001202047, 0.001186867, 0.00112739, 
    0.0009925561, 0.0008747317, 0.000805256, 0.0007760101, 0.0007839249, 
    0.0007820339, 0.00080756, 0.0008660844, 0.0009420286, 0.001124896, 
    0.001172421, 0.001045534, 0.000973992, 0.0008369819, 0.0007515, 
    0.0008409866, 0.0009124493, 0.0009461134, 0.0009490061, 0.0008171932, 
    0.001148928, 0.001344511, 0.001509513, 0.001576811, 0.001659143, 
    0.001748201, 0.001714631, 0.001378971, 0.00146383, 0.00139577, 
    0.001283729, 0.001256978, 0.001216114, 0.001151281, 0.001115693, 
    0.001064321, 0.001002619, 0.0009573349, 0.0009314744, 0.0009110975, 
    0.0009421399, 0.0009748512, 0.0009923829, 0.00102743, 0.001026794, 
    0.001016558, 0.0009905868, 0.0009698919, 0.0009588771, 0.0009115264, 
    0.0008804216, 0.0008716313, 0.0008271742, 0.0007815408, 0.0006749365, 
    0.0006103888, 0.0005978951, 0.0004962655, 0.00052416, 0.0006104838, 
    0.0008088481, 0.0009558727, 0.001211219, 0.001430914, 0.001640419, 
    0.001578605, 0.00143565, 0.001349152, 0.001295524, 0.001234186, 
    0.001179223, 0.001137945, 0.001109335, 0.001040957, 0.00101926, 
    0.001061127,
  0.001157559, 0.001102054, 0.001029146, 0.001057041, 0.001211535, 
    0.00133335, 0.001535609, 0.001568464, 0.001677277, 0.001722943, 
    0.001301165, 0.001180778, 0.00114802, 0.001085682, 0.00108174, 
    0.001065385, 0.001079896, 0.001058264, 0.0009133527, 0.0007645646, 
    0.0006522378, 0.000653049, 0.0007147351, 0.0007722909, 0.0009161355, 
    0.001004542, 0.001078786, 0.001224491, 0.001341745, 0.001382434, 
    0.001182066, 0.001049904, 0.0009904429, 0.000952757, 0.0009731026, 
    0.001031674, 0.0009704162, 0.000836377, 0.0008396362, 0.0007672203, 
    0.0009046602, 0.001669618, 0.002085848, 0.002075517, 0.00198433, 
    0.00196338, 0.001769149, 0.001552076, 0.001375948, 0.001092326, 
    0.0009811269, 0.001031243, 0.001079325, 0.001136005, 0.001146416, 
    0.001143984, 0.001099336, 0.001063971, 0.001090134, 0.001102674, 
    0.001103452, 0.001133589, 0.001188012, 0.001231372, 0.001239033, 
    0.001249842, 0.00124075, 0.001195926, 0.001104691, 0.0009855293, 
    0.0009084251, 0.0008274587, 0.0007280707, 0.0007064864, 0.0006876346, 
    0.0006556399, 0.0006132182, 0.0005808403, 0.0006650337, 0.0008122493, 
    0.0009619291, 0.001275131, 0.001827131, 0.002142941, 0.002036495, 
    0.001910642, 0.001747579, 0.001548119, 0.001414159, 0.001347625, 
    0.001307506, 0.001254863, 0.001230449, 0.001194894, 0.001174899, 
    0.001190777,
  0.001202698, 0.001162468, 0.001083059, 0.001165949, 0.001256374, 
    0.0009112088, 0.0008239956, 0.001178031, 0.001678662, 0.00184142, 
    0.001694301, 0.001653928, 0.001661272, 0.001463765, 0.001405815, 
    0.001402237, 0.001365093, 0.001385071, 0.001278006, 0.00120478, 
    0.001200107, 0.001264178, 0.001338897, 0.001338437, 0.001400966, 
    0.001450208, 0.001456375, 0.001512975, 0.001502087, 0.001362152, 
    0.001237968, 0.0009374507, 0.0009447951, 0.0009772829, 0.001013109, 
    0.001155255, 0.001052751, 0.001053561, 0.001224778, 0.001103868, 
    0.00117223, 0.001857871, 0.001868553, 0.001877375, 0.001840706, 
    0.00176527, 0.001557162, 0.00135697, 0.001244882, 0.001111336, 
    0.001140566, 0.001174437, 0.001206178, 0.001280819, 0.001312434, 
    0.001345065, 0.001314182, 0.001277179, 0.001299305, 0.001312243, 
    0.001294584, 0.001296842, 0.001368827, 0.001452179, 0.00148907, 
    0.001461668, 0.001374359, 0.001168525, 0.0009667901, 0.0008152677, 
    0.0007246844, 0.0007024482, 0.0007147975, 0.000690368, 0.0006383145, 
    0.0005523879, 0.000601518, 0.0008151261, 0.0009716088, 0.001159738, 
    0.001238653, 0.00153159, 0.001880379, 0.002160346, 0.002106002, 
    0.001807104, 0.001601413, 0.001491772, 0.001444279, 0.001370226, 
    0.001364791, 0.001342173, 0.001349897, 0.001377919, 0.001342888, 
    0.001277084,
  0.001245803, 0.001225283, 0.001282489, 0.00151269, 0.001639847, 
    0.0008956012, 0.0009100488, 0.001301215, 0.001882256, 0.002186046, 
    0.002080904, 0.001949393, 0.001934913, 0.001840483, 0.001844964, 
    0.001916014, 0.001844647, 0.001778971, 0.001720098, 0.001718746, 
    0.001713883, 0.001682714, 0.001685671, 0.001683222, 0.00166461, 
    0.001641372, 0.001607325, 0.001533511, 0.001534529, 0.001573645, 
    0.001481377, 0.001055962, 0.001139901, 0.001237954, 0.000958432, 
    0.001181575, 0.001413891, 0.001501693, 0.001500485, 0.001549011, 
    0.001613574, 0.001792355, 0.001614701, 0.001581719, 0.001604767, 
    0.001604591, 0.001624078, 0.001640577, 0.001636921, 0.001588745, 
    0.001531286, 0.001415955, 0.001379445, 0.001436125, 0.001426334, 
    0.001402111, 0.001398169, 0.001425794, 0.001465737, 0.001524181, 
    0.001567207, 0.0015955, 0.001606943, 0.001647634, 0.001672191, 
    0.001547291, 0.001408898, 0.001215271, 0.0009929687, 0.0008504568, 
    0.000707374, 0.0007052291, 0.0006574821, 0.0005827462, 0.0005748151, 
    0.0006376151, 0.001114292, 0.001148706, 0.001192177, 0.001512278, 
    0.001538996, 0.001773917, 0.001886992, 0.002003196, 0.002145167, 
    0.001869459, 0.001601079, 0.001521558, 0.001498876, 0.001449763, 
    0.001441657, 0.0014195, 0.001421582, 0.001395276, 0.001382513, 0.00132197,
  0.001385406, 0.001536245, 0.001811873, 0.002065756, 0.001206165, 
    0.0008683731, 0.001261652, 0.001497878, 0.001821825, 0.002117367, 
    0.00231101, 0.002210175, 0.002255029, 0.002206647, 0.002095575, 
    0.00203578, 0.001992706, 0.00196036, 0.001920878, 0.001903521, 
    0.001901153, 0.001849622, 0.001778717, 0.001761104, 0.001743939, 
    0.001777635, 0.001871844, 0.001884192, 0.001847618, 0.001821711, 
    0.0017063, 0.001127121, 0.00110614, 0.001093059, 0.0009909999, 
    0.001565462, 0.001746994, 0.001597568, 0.001585218, 0.001844332, 
    0.001951841, 0.001925184, 0.001954573, 0.002088167, 0.002115601, 
    0.002036224, 0.001985203, 0.001936136, 0.001837049, 0.001663974, 
    0.001546927, 0.001461349, 0.00138574, 0.001346845, 0.001404035, 
    0.001458998, 0.001500228, 0.001588125, 0.001701309, 0.001853356, 
    0.001958658, 0.002012763, 0.002028308, 0.001945688, 0.001837176, 
    0.001630547, 0.001394894, 0.001203444, 0.001003427, 0.0009266092, 
    0.0008540032, 0.0007872758, 0.0006836122, 0.0006820066, 0.0006876336, 
    0.0009579686, 0.00189702, 0.001426702, 0.001005352, 0.001879934, 
    0.001761837, 0.001699006, 0.001898451, 0.001795835, 0.002047827, 
    0.002003687, 0.001763791, 0.001636396, 0.001617006, 0.001578015, 
    0.001510638, 0.001443865, 0.001412013, 0.001360165, 0.001371419, 
    0.001341632,
  0.001824412, 0.002018359, 0.002309054, 0.002453918, 0.001510578, 
    0.001398234, 0.001860178, 0.00188804, 0.001849353, 0.002039229, 
    0.002467586, 0.00233129, 0.001837113, 0.001994327, 0.002209379, 
    0.002111151, 0.002025574, 0.002015338, 0.002037718, 0.002055663, 
    0.002093985, 0.002136582, 0.002138235, 0.002157467, 0.002255855, 
    0.002331847, 0.002330051, 0.00226234, 0.002159932, 0.002095081, 
    0.002050959, 0.001838385, 0.001300308, 0.0008712336, 0.0013842, 
    0.001346959, 0.001423777, 0.001779641, 0.002181676, 0.002277568, 
    0.002332373, 0.002435862, 0.002564068, 0.002675314, 0.002625913, 
    0.002451278, 0.002282254, 0.002122737, 0.001973265, 0.001817022, 
    0.001732176, 0.001691154, 0.001619834, 0.001635299, 0.001809392, 
    0.001943177, 0.002016197, 0.00209718, 0.00216834, 0.002282891, 
    0.002378721, 0.002445971, 0.002383282, 0.002166702, 0.001988764, 
    0.001811044, 0.001563742, 0.001388775, 0.001264702, 0.001169414, 
    0.001057199, 0.0009701913, 0.0009110318, 0.0009266399, 0.001020735, 
    0.001564029, 0.002421129, 0.001593229, 0.001255898, 0.00218886, 
    0.001805738, 0.002187239, 0.00246158, 0.001747293, 0.001873385, 
    0.002103507, 0.002002431, 0.001991274, 0.001913946, 0.001784137, 
    0.001743526, 0.00168114, 0.001631485, 0.001603669, 0.001597438, 
    0.001639336,
  0.002349538, 0.002464488, 0.002799197, 0.002865045, 0.001967784, 
    0.001518047, 0.001764794, 0.001751444, 0.001958166, 0.002009888, 
    0.002278187, 0.002507259, 0.002117239, 0.002107766, 0.002182709, 
    0.002156212, 0.002163412, 0.002222175, 0.002302378, 0.002397364, 
    0.002504668, 0.002562572, 0.002610384, 0.002648165, 0.002718259, 
    0.002716481, 0.00265314, 0.002580803, 0.00258093, 0.00266549, 
    0.002731547, 0.002637484, 0.002381263, 0.002390594, 0.002447275, 
    0.002091905, 0.002159407, 0.002821782, 0.002745122, 0.002832322, 
    0.003020353, 0.003188804, 0.003165565, 0.003110252, 0.002963512, 
    0.002713175, 0.002507387, 0.002309546, 0.002154829, 0.00204514, 
    0.002006454, 0.001985153, 0.002020488, 0.002176335, 0.002375161, 
    0.002530022, 0.002649311, 0.002724921, 0.002725653, 0.002723759, 
    0.002759315, 0.002761271, 0.002605567, 0.002422287, 0.002263024, 
    0.002169197, 0.001985805, 0.00186426, 0.001779575, 0.001679057, 
    0.001582594, 0.001573057, 0.00160065, 0.001571849, 0.001729841, 
    0.002158723, 0.002153432, 0.00171956, 0.001846191, 0.002318338, 
    0.001971534, 0.002192612, 0.002124646, 0.002142511, 0.001827132, 
    0.001945165, 0.002172457, 0.002174128, 0.002135708, 0.002090488, 
    0.002125202, 0.002094701, 0.002051118, 0.002034842, 0.002095289, 
    0.00218398,
  0.002798765, 0.002864935, 0.003131169, 0.003097615, 0.001836239, 
    0.001379177, 0.001826575, 0.001808886, 0.002022604, 0.001988255, 
    0.002191563, 0.002573413, 0.002453568, 0.002309245, 0.002320133, 
    0.002340462, 0.002442043, 0.00251635, 0.002632778, 0.0027075, 
    0.002799036, 0.002868829, 0.002919804, 0.003032403, 0.003090052, 
    0.003015809, 0.003028013, 0.003066735, 0.003180174, 0.003262762, 
    0.003239572, 0.00333548, 0.003306041, 0.003130168, 0.002969379, 
    0.002954183, 0.003191027, 0.003293977, 0.003217859, 0.003229158, 
    0.003494788, 0.003495157, 0.003394257, 0.003253449, 0.00305769, 
    0.002794569, 0.002600132, 0.002473054, 0.002435988, 0.002489442, 
    0.002544135, 0.002589989, 0.002696341, 0.002826963, 0.002955232, 
    0.003006173, 0.003088301, 0.003159573, 0.003124762, 0.003097519, 
    0.003057389, 0.003030304, 0.002943074, 0.002852838, 0.002726477, 
    0.002614546, 0.002495608, 0.002442298, 0.002356293, 0.002250832, 
    0.002226211, 0.002197411, 0.002197426, 0.002176525, 0.002227864, 
    0.002529195, 0.002267729, 0.001970613, 0.002028611, 0.001631725, 
    0.001607007, 0.001365729, 0.001968355, 0.002434081, 0.001711436, 
    0.00186016, 0.002325568, 0.002422494, 0.002430694, 0.002491381, 
    0.00251411, 0.002513713, 0.002566085, 0.002580645, 0.00265821, 0.002713587,
  0.003040426, 0.003073789, 0.003333049, 0.00334907, 0.002329464, 
    0.002119274, 0.002349205, 0.002166767, 0.00198932, 0.002067744, 
    0.002323964, 0.002749332, 0.002551079, 0.002540208, 0.002620714, 
    0.00265586, 0.002784526, 0.002845528, 0.003024263, 0.003075983, 
    0.003150353, 0.00324332, 0.003295027, 0.003293674, 0.003326749, 
    0.003345298, 0.003398642, 0.003473043, 0.003530232, 0.00358998, 
    0.003597498, 0.003569795, 0.003564281, 0.003563564, 0.003530076, 
    0.003335528, 0.003383782, 0.003391812, 0.003126529, 0.003437173, 
    0.003656548, 0.003571145, 0.003457943, 0.0032763, 0.003031906, 
    0.002838675, 0.002653567, 0.002569262, 0.002509659, 0.002592262, 
    0.002670573, 0.002691237, 0.00281194, 0.002963575, 0.003083451, 
    0.003100887, 0.003162131, 0.003250852, 0.003204603, 0.003226981, 
    0.003177088, 0.003160048, 0.003163436, 0.003122509, 0.003077321, 
    0.002979519, 0.002896739, 0.002835577, 0.002760285, 0.00272228, 
    0.002718863, 0.002663231, 0.002634557, 0.002610525, 0.002635369, 
    0.002587353, 0.001752237, 0.001654644, 0.00166461, 0.001324355, 
    0.00135554, 0.001470267, 0.001611586, 0.002390991, 0.002339669, 
    0.002241074, 0.002388607, 0.002688726, 0.002684975, 0.002771283, 
    0.002835322, 0.002844017, 0.002869019, 0.002910439, 0.002980598, 
    0.002954468,
  0.003228668, 0.003297016, 0.003332553, 0.003214506, 0.003074933, 
    0.002595953, 0.002581297, 0.002732136, 0.002408746, 0.002117938, 
    0.002240183, 0.002573619, 0.002664249, 0.002645655, 0.002769249, 
    0.002844812, 0.0030156, 0.003212705, 0.003335906, 0.003346857, 
    0.003334062, 0.003270976, 0.003282659, 0.003316185, 0.003431246, 
    0.003480788, 0.003549499, 0.003493028, 0.003240827, 0.003467308, 
    0.00347797, 0.003414838, 0.003401326, 0.003439823, 0.003485998, 
    0.003423166, 0.003318103, 0.00320085, 0.003047373, 0.003146619, 
    0.003587961, 0.003437329, 0.00326111, 0.00308077, 0.00286144, 0.00275323, 
    0.002652697, 0.002618317, 0.002637455, 0.002688363, 0.002814997, 
    0.002978314, 0.003147369, 0.003299795, 0.003355173, 0.003380463, 
    0.003376976, 0.003401184, 0.003381109, 0.003365677, 0.003278576, 
    0.003244132, 0.003233451, 0.003181826, 0.003124241, 0.003080817, 
    0.003066162, 0.003008369, 0.002974642, 0.002953613, 0.002915163, 
    0.002842352, 0.002826393, 0.002780057, 0.002905292, 0.002991838, 
    0.001867965, 0.002298056, 0.002376941, 0.001727567, 0.00179275, 
    0.001692568, 0.001932225, 0.002202911, 0.002857099, 0.002700649, 
    0.002681606, 0.002804553, 0.003000451, 0.003111046, 0.003140023, 
    0.003163928, 0.003198167, 0.003221914, 0.003166489, 0.003148131,
  0.003366297, 0.003444944, 0.003305692, 0.002583443, 0.003563295, 
    0.002758888, 0.002348061, 0.002674073, 0.002934029, 0.002335122, 
    0.002440329, 0.002561158, 0.002704466, 0.002806015, 0.002935966, 
    0.003086999, 0.003213421, 0.003403271, 0.003392398, 0.003339805, 
    0.003377872, 0.00331364, 0.003366426, 0.003433121, 0.003500003, 
    0.003351709, 0.003373357, 0.003291547, 0.003055926, 0.003465608, 
    0.003053492, 0.003048278, 0.002920549, 0.003376838, 0.00347222, 
    0.003162196, 0.002783064, 0.002753038, 0.003097158, 0.003404759, 
    0.003524197, 0.003172815, 0.003032815, 0.003010403, 0.002970191, 
    0.002972273, 0.002995258, 0.003065463, 0.003289878, 0.003469534, 
    0.003656153, 0.003893537, 0.003929682, 0.003907919, 0.00378553, 
    0.003595877, 0.003432944, 0.003281564, 0.003182031, 0.003086157, 
    0.003021831, 0.002992921, 0.00299521, 0.003005922, 0.003044054, 
    0.003053684, 0.003025234, 0.003036359, 0.003088765, 0.003041446, 
    0.003109444, 0.003010627, 0.003033118, 0.002949448, 0.003009353, 
    0.003296504, 0.002316462, 0.002965531, 0.003094484, 0.002496864, 
    0.002989946, 0.002807572, 0.002341717, 0.002773907, 0.002949779, 
    0.002935316, 0.002894389, 0.003029, 0.003242223, 0.003317118, 
    0.003269451, 0.003342042, 0.003363213, 0.003290974, 0.003204301, 
    0.003294835,
  0.003274918, 0.00345435, 0.003303703, 0.002628057, 0.003308091, 
    0.003686572, 0.003073169, 0.002979455, 0.003112857, 0.002993729, 
    0.002842444, 0.002698852, 0.002560364, 0.002824262, 0.003041476, 
    0.003080877, 0.003225043, 0.003347814, 0.003343031, 0.003203984, 
    0.003205622, 0.003207339, 0.003268786, 0.003288209, 0.003388265, 
    0.003276702, 0.003193462, 0.003170589, 0.003261903, 0.003476497, 
    0.003306217, 0.002847912, 0.002546297, 0.003001742, 0.003119027, 
    0.002946811, 0.002881944, 0.002907677, 0.003189504, 0.003477672, 
    0.003370926, 0.003093215, 0.003103863, 0.00308422, 0.003088335, 
    0.003057817, 0.003120936, 0.003172051, 0.003296793, 0.003463002, 
    0.003642833, 0.00384363, 0.003890958, 0.003883664, 0.003814589, 
    0.003696682, 0.003640559, 0.00348282, 0.003366124, 0.003266655, 
    0.00313767, 0.003047582, 0.003046723, 0.003012899, 0.003036043, 
    0.002995098, 0.002988454, 0.003056897, 0.003018349, 0.002936762, 
    0.002995556, 0.002830507, 0.002751002, 0.002686772, 0.002625277, 
    0.002862425, 0.002788069, 0.003084931, 0.003566856, 0.002997496, 
    0.002843143, 0.002413927, 0.002537396, 0.003198974, 0.00312883, 
    0.003139542, 0.002981313, 0.00294172, 0.002970029, 0.003050169, 
    0.003188912, 0.00328172, 0.003233798, 0.003244957, 0.003236199, 
    0.003238456,
  0.003014393, 0.003377711, 0.002957126, 0.002836835, 0.003160719, 
    0.003379412, 0.003226936, 0.00299303, 0.00322805, 0.00310008, 
    0.002713143, 0.002604963, 0.002184201, 0.002916705, 0.003094563, 
    0.003209751, 0.003384341, 0.003318204, 0.003235137, 0.003198197, 
    0.003233453, 0.003107836, 0.003063366, 0.003207179, 0.003294488, 
    0.003212409, 0.002951993, 0.003183845, 0.003085332, 0.003100891, 
    0.003045183, 0.002831716, 0.002727099, 0.002962941, 0.002964899, 
    0.0029041, 0.003004795, 0.002992826, 0.003092641, 0.003147891, 
    0.003155252, 0.003071567, 0.003064604, 0.00300853, 0.003072837, 
    0.003093502, 0.00308034, 0.003033515, 0.003024504, 0.003055418, 
    0.0030839, 0.003081977, 0.003158065, 0.003177727, 0.003221055, 
    0.003248807, 0.003278149, 0.003259849, 0.00327355, 0.003242653, 
    0.003233338, 0.003323985, 0.003391614, 0.003302097, 0.003334394, 
    0.00330607, 0.003363578, 0.0033271, 0.003256785, 0.003280755, 
    0.003093243, 0.002929384, 0.002828917, 0.002833366, 0.002732517, 
    0.002753783, 0.002722488, 0.002807619, 0.003040476, 0.002252056, 
    0.002546059, 0.002888875, 0.002923446, 0.002901271, 0.003073677, 
    0.003115701, 0.002936255, 0.002975672, 0.002922202, 0.002959553, 
    0.003143104, 0.003246041, 0.003139755, 0.003118424, 0.002819002, 
    0.002807494,
  0.003019271, 0.003068577, 0.003033496, 0.00294867, 0.003022896, 
    0.003120789, 0.003084932, 0.003007066, 0.003412105, 0.003334509, 
    0.002804218, 0.00321123, 0.002404452, 0.002164667, 0.002990931, 
    0.003022004, 0.003325287, 0.003355585, 0.003352378, 0.003317503, 
    0.003150037, 0.002920549, 0.003109979, 0.003186516, 0.003145779, 
    0.003128739, 0.003212646, 0.003242606, 0.003198452, 0.00307573, 
    0.003180889, 0.003137894, 0.003015362, 0.002975561, 0.002963087, 
    0.002836756, 0.002964247, 0.002956871, 0.002984496, 0.003059074, 
    0.003083488, 0.00302266, 0.002998101, 0.003003156, 0.003073983, 
    0.003103593, 0.00309881, 0.003076002, 0.003119426, 0.003116658, 
    0.003122875, 0.003085045, 0.003061442, 0.003030686, 0.003055561, 
    0.002992028, 0.002972161, 0.002999436, 0.003096011, 0.003149912, 
    0.003180522, 0.003214698, 0.003209945, 0.003091227, 0.003142616, 
    0.003165694, 0.003332825, 0.003383562, 0.003430195, 0.003400521, 
    0.003186405, 0.003109284, 0.002693085, 0.002615903, 0.002593488, 
    0.002568582, 0.002777021, 0.002789706, 0.003061347, 0.002732869, 
    0.00291435, 0.002827313, 0.002878953, 0.002806745, 0.002769791, 
    0.002830762, 0.002781203, 0.002862042, 0.002885964, 0.002920169, 
    0.003059864, 0.003081704, 0.003093723, 0.003030384, 0.00309086, 
    0.003098855,
  0.003209496, 0.003115876, 0.003064841, 0.003142469, 0.003249565, 
    0.003162228, 0.002853716, 0.002878301, 0.003353627, 0.00339235, 
    0.003017443, 0.002521676, 0.002352081, 0.001705348, 0.002991347, 
    0.002774321, 0.003015742, 0.003317995, 0.003338261, 0.003366299, 
    0.002872819, 0.002764134, 0.003191808, 0.003176915, 0.003123479, 
    0.003310207, 0.003347987, 0.002971699, 0.002967887, 0.003124129, 
    0.003356334, 0.003295917, 0.003067113, 0.003019573, 0.003033977, 
    0.00285602, 0.002963357, 0.002971144, 0.002925368, 0.002964754, 
    0.003002584, 0.003082708, 0.0031316, 0.003113417, 0.00311375, 
    0.003063507, 0.003062919, 0.003061645, 0.003078811, 0.003062421, 
    0.003097963, 0.00307072, 0.003043398, 0.003081944, 0.003123714, 
    0.003115751, 0.003143584, 0.003123667, 0.003149463, 0.003196035, 
    0.003164977, 0.003090035, 0.003077714, 0.003021447, 0.003020529, 
    0.003045293, 0.003274016, 0.003469454, 0.003505696, 0.003445661, 
    0.003423456, 0.002829762, 0.002750274, 0.00219463, 0.002472529, 
    0.002571838, 0.002719181, 0.002723156, 0.002743881, 0.002774861, 
    0.002733152, 0.00261806, 0.002616281, 0.002576036, 0.002539702, 
    0.002528688, 0.002557853, 0.002621528, 0.00264192, 0.002708025, 
    0.002786685, 0.002802834, 0.003197098, 0.003370255, 0.003360735, 
    0.00322248,
  0.002784653, 0.002322992, 0.002550541, 0.002965452, 0.00304612, 
    0.002999119, 0.002124138, 0.002193058, 0.00286638, 0.00282806, 
    0.003096744, 0.002456571, 0.001759025, 0.002415392, 0.002483292, 
    0.002940675, 0.002696259, 0.003013404, 0.003081867, 0.003196212, 
    0.00279527, 0.002782967, 0.003371464, 0.003382968, 0.003160177, 
    0.003044685, 0.002714112, 0.002690174, 0.002853539, 0.003194861, 
    0.003256865, 0.003303627, 0.003126761, 0.002910981, 0.002906499, 
    0.002886394, 0.002880607, 0.00289903, 0.002911985, 0.002922777, 
    0.002961067, 0.00299737, 0.002995925, 0.003011296, 0.003057532, 
    0.003059754, 0.003037326, 0.002982855, 0.002930215, 0.002899315, 
    0.002885168, 0.002855938, 0.002878018, 0.00289, 0.002896138, 0.002904229, 
    0.002906326, 0.002871184, 0.00288091, 0.002893483, 0.002890702, 
    0.002924891, 0.002785431, 0.002617059, 0.002455316, 0.00238042, 
    0.002808003, 0.003355062, 0.003625285, 0.003124366, 0.002884598, 
    0.002498612, 0.00155476, 0.002576591, 0.002632381, 0.002606014, 
    0.002577499, 0.002594234, 0.002597874, 0.002557693, 0.00251467, 
    0.002553547, 0.002509072, 0.002417566, 0.002448894, 0.002348997, 
    0.00235421, 0.002319131, 0.002308402, 0.002297277, 0.002388416, 
    0.002577052, 0.002098784, 0.00143207, 0.001382479, 0.002718849,
  0.001647444, 0.001603273, 0.001409424, 0.001750425, 0.0008323081, 
    0.001562394, 0.001157368, 0.001235585, 0.001696814, 0.002250802, 
    0.003262011, 0.002183282, 0.001777383, 0.002163034, 0.003724023, 
    0.003619975, 0.002838073, 0.002909647, 0.003030606, 0.003337974, 
    0.003179358, 0.003189549, 0.003324671, 0.003390346, 0.003371745, 
    0.002870787, 0.00272592, 0.002737239, 0.00298173, 0.003112035, 
    0.003107265, 0.003178058, 0.003165798, 0.002876395, 0.002734758, 
    0.002826629, 0.002761684, 0.002815679, 0.002910253, 0.002873249, 
    0.002858516, 0.002856784, 0.002938576, 0.002954943, 0.002868477, 
    0.00286792, 0.002757901, 0.002705909, 0.002658004, 0.002575368, 
    0.002593758, 0.002623195, 0.002661631, 0.002676873, 0.002709724, 
    0.002658004, 0.002627263, 0.002572299, 0.00250721, 0.002506942, 
    0.002412638, 0.002386936, 0.002274213, 0.002103427, 0.001567716, 
    0.001262318, 0.001778476, 0.002335055, 0.002685867, 0.002676663, 
    0.002283527, 0.001797471, 0.00197808, 0.002826579, 0.002618583, 
    0.002625817, 0.002550589, 0.002451008, 0.002454776, 0.002540005, 
    0.002521344, 0.00240439, 0.002391452, 0.002365766, 0.002347026, 
    0.00224379, 0.002195963, 0.002114885, 0.002090773, 0.002034158, 
    0.00196934, 0.00212463, 0.001439828, -0.000128773, -0.001003689, 
    0.0006959178,
  0.00165644, 0.001776492, 0.0009297896, 0.0009589409, 0.001044676, 
    0.001093393, 0.0005956376, 0.0007247811, 0.000740103, 0.001727901, 
    0.002867592, 0.00157886, 0.001789734, 0.00228194, 0.003704362, 
    0.00554635, 0.004009008, 0.003637297, 0.003491994, 0.003402302, 
    0.003369048, 0.003430244, 0.003330311, 0.002988037, 0.003021255, 
    0.003014473, 0.002827471, 0.00283882, 0.003114529, 0.003206512, 
    0.002855172, 0.003011247, 0.0029789, 0.00291273, 0.002718788, 
    0.002717961, 0.00270677, 0.002656937, 0.002719069, 0.00273552, 
    0.002740337, 0.00273994, 0.002797954, 0.002776863, 0.002686042, 
    0.002656525, 0.002513586, 0.002439547, 0.002412574, 0.002363559, 
    0.002363525, 0.002337856, 0.002355896, 0.002352064, 0.002371805, 
    0.002320084, 0.002323295, 0.002293399, 0.002177065, 0.002135088, 
    0.002039022, 0.002020568, 0.00203964, 0.001855043, 0.001381034, 
    0.00128667, 0.001440573, 0.002082875, 0.002170946, 0.002793044, 
    0.002915053, 0.002853155, 0.002738954, 0.002793932, 0.002777927, 
    0.002686407, 0.002524044, 0.00262801, 0.002685167, 0.00255752, 
    0.00252638, 0.002501713, 0.002476884, 0.002393628, 0.00231619, 
    0.002275882, 0.002206614, 0.002139237, 0.002059842, 0.002002193, 
    0.001853198, 0.001908527, 0.001372897, 0.001356795, 0.00137989, 
    0.0009870105,
  0.0006419388, 0.001552632, 0.001622902, 0.001220407, 0.00172051, 
    0.00170948, 0.001004463, 0.0007206011, 0.001113992, 0.001133622, 
    0.001611079, 0.001335802, 0.001902107, 0.001747007, 0.003099635, 
    0.004076087, 0.004360185, 0.00429977, 0.004471308, 0.004004642, 
    0.003815044, 0.003352391, 0.003080482, 0.002827297, 0.002760873, 
    0.00286333, 0.002660673, 0.002701506, 0.003339279, 0.00351561, 
    0.003207048, 0.003102938, 0.003230814, 0.003009101, 0.002901303, 
    0.002732515, 0.002712093, 0.002688123, 0.00266058, 0.002634909, 
    0.002586778, 0.00260199, 0.002598559, 0.002558837, 0.00251667, 
    0.002409207, 0.002289997, 0.002159787, 0.00207836, 0.002120273, 
    0.002187429, 0.002257174, 0.002271034, 0.002182993, 0.002108354, 
    0.002043502, 0.001956353, 0.001921115, 0.001879328, 0.001825605, 
    0.001816133, 0.001818517, 0.001734323, 0.001521464, 0.001401966, 
    0.001684191, 0.001511831, 0.002358614, 0.002619555, 0.002915213, 
    0.002901571, 0.002991803, 0.002883913, 0.002926208, 0.002715765, 
    0.002442377, 0.002420571, 0.002514446, 0.002578977, 0.002526443, 
    0.002506003, 0.002422016, 0.002389766, 0.002406486, 0.002333483, 
    0.002250769, 0.002187541, 0.002138826, 0.002052549, 0.00196891, 
    0.001844345, 0.001793975, 0.002084718, 0.001635379, 0.00160909, 
    8.502509e-005,
  0.001218482, 0.0009084116, 0.0001602059, 0.001280501, 0.001712628, 
    0.002338856, 0.002102885, 0.001550726, 0.00260633, 0.002286961, 
    0.002091316, 0.001816817, 0.002097562, 0.002613055, 0.002261483, 
    0.002002832, 0.002125647, 0.002475027, 0.003622169, 0.004465962, 
    0.004157199, 0.003199245, 0.002938734, 0.002291968, 0.002429998, 
    0.002444254, 0.002250213, 0.00265047, 0.003377647, 0.003701562, 
    0.003652859, 0.003543871, 0.003556093, 0.002413847, 0.002740465, 
    0.002794968, 0.00277343, 0.002657799, 0.002600165, 0.002544867, 
    0.002495181, 0.002505623, 0.002487231, 0.002442664, 0.002411954, 
    0.002375017, 0.002325456, 0.002182756, 0.002066726, 0.00201324, 
    0.002033983, 0.002143782, 0.00220542, 0.002158706, 0.002093761, 
    0.001999824, 0.001869252, 0.001753015, 0.001715203, 0.001700628, 
    0.001691201, 0.001638192, 0.001567191, 0.001537803, 0.001628768, 
    0.002371042, 0.002706578, 0.002846514, 0.002783936, 0.002687139, 
    0.002748827, 0.002770493, 0.002818525, 0.00274959, 0.00265203, 
    0.002552019, 0.002401369, 0.002216185, 0.002274213, 0.002326522, 
    0.002269207, 0.002166655, 0.00215688, 0.002193833, 0.002091267, 
    0.002077807, 0.002099424, 0.002039499, 0.002029373, 0.002002448, 
    0.00192458, 0.001797743, 0.001838957, 0.002126933, 0.002515128, 
    0.001539853,
  0.002577928, 0.00257316, 0.002116874, 0.002176525, 0.002284911, 
    0.002407362, 0.002337983, 0.002333278, 0.002793933, 0.00243416, 
    0.002998894, 0.002594918, 0.002550192, 0.003170891, 0.002893307, 
    0.002326062, 0.002745186, 0.00236742, 0.002038307, 0.002087866, 
    0.002220983, 0.002301871, 0.002152065, 0.001867758, 0.002287423, 
    0.002355213, 0.002088947, 0.002481798, 0.002994779, 0.0031031, 
    0.003102399, 0.003185894, 0.003143074, 0.002292586, 0.002818428, 
    0.002775161, 0.002706068, 0.002709692, 0.002433747, 0.002396824, 
    0.002340939, 0.002262658, 0.002229343, 0.002259606, 0.002239881, 
    0.002195185, 0.002202115, 0.002193183, 0.002112471, 0.002022619, 
    0.001970374, 0.00196748, 0.001984376, 0.002032425, 0.002017929, 
    0.00195025, 0.001926154, 0.001811633, 0.001674019, 0.001649414, 
    0.001617895, 0.001548977, 0.001598425, 0.001508555, 0.00273231, 
    0.003054271, 0.00300187, 0.002733663, 0.003188898, 0.002676062, 
    0.002680717, 0.002712555, 0.003106788, 0.002958078, 0.002841635, 
    0.002884153, 0.002805173, 0.002585908, 0.002432954, 0.002306161, 
    0.002255395, 0.00221127, 0.002049622, 0.001883938, 0.001707143, 
    0.001623871, 0.00160982, 0.001662956, 0.001787489, 0.001829532, 
    0.001861082, 0.001793197, 0.001696717, 0.001908576, 0.001847143, 
    0.002669813,
  0.003162452, 0.002206678, 0.002290378, 0.002374207, 0.002346326, 
    0.002340303, 0.003564551, 0.002828185, 0.002484865, 0.00251063, 
    0.003057547, 0.003137242, 0.003087523, 0.003113987, 0.002697661, 
    0.002353305, 0.001579099, 0.00158924, 0.002572094, 0.001978686, 
    0.002331642, 0.00140143, 0.0007495927, 0.00103827, 0.001489533, 
    0.0015403, 0.001746117, 0.002131417, 0.0027061, 0.002677857, 0.002283908, 
    0.002493335, 0.002757551, 0.002769504, 0.00286805, 0.002504001, 
    0.002317972, 0.002451691, 0.002349219, 0.002321245, 0.002266202, 
    0.002223955, 0.002111073, 0.002085689, 0.002074229, 0.00198746, 
    0.001957118, 0.001988064, 0.001990004, 0.001921752, 0.001874132, 
    0.001828053, 0.001757021, 0.001734927, 0.001703058, 0.00167812, 
    0.001694714, 0.00163166, 0.001535498, 0.001507015, 0.001475575, 
    0.001450812, 0.001560326, 0.00227725, 0.002908043, 0.002538811, 
    0.002146389, 0.002586225, 0.003060836, 0.003236105, 0.002903162, 
    0.002864793, 0.002801741, 0.002785619, 0.002697932, 0.002797034, 
    0.002956043, 0.003019399, 0.002975387, 0.002623528, 0.002482973, 
    0.002434033, 0.002191896, 0.00183991, 0.00138666, 0.000831686, 
    0.0005929973, 0.0008848859, 0.001270456, 0.001456057, 0.001583038, 
    0.001621152, 0.001619213, 0.001809726, 0.002698933, 0.00318332,
  0.002459512, 0.002030359, 0.0019259, 0.002773431, 0.001333748, 0.002401005, 
    0.002031917, 0.002183455, 0.002063022, 0.002084482, 0.002043839, 
    0.001913565, 0.001887229, 0.001817164, 0.001931733, 0.001639972, 
    0.00151134, 0.0009829409, 0.0015029, 0.00187399, 0.002139222, 
    0.002386764, 0.002431538, 0.002278665, 0.001589955, 0.001128281, 
    0.00114788, 0.001398569, 0.002016372, 0.002425658, 0.002312917, 
    0.002486136, 0.002583395, 0.002706259, 0.002673755, 0.002515939, 
    0.001945738, 0.002026513, 0.002371727, 0.001937695, 0.001783947, 
    0.001655806, 0.001526472, 0.001493729, 0.001468806, 0.001412651, 
    0.001350486, 0.001358195, 0.001416529, 0.001453689, 0.001496525, 
    0.001479439, 0.001436666, 0.001375169, 0.001340932, 0.001365236, 
    0.001378348, 0.001357018, 0.001313276, 0.001367763, 0.001378762, 
    0.001362914, 0.001500323, 0.001726344, 0.002408476, 0.002425133, 
    0.002232173, 0.003032815, 0.003155377, 0.003199246, 0.003164213, 
    0.00293635, 0.002788131, 0.002648769, 0.002751242, 0.002761272, 
    0.002894134, 0.00280107, 0.002515224, 0.00230052, 0.001967114, 
    0.001782293, 0.001672843, 0.001410058, 0.001089274, 0.0007289751, 
    0.0004578773, 0.0005097259, 0.0007548034, 0.001028317, 0.001268009, 
    0.001369384, 0.001416082, 0.001658283, 0.002476553, 0.002556709,
  0.002129684, 0.002084973, 0.002165464, 0.002120577, 0.001856776, 
    0.001897862, 0.00191886, 0.001766891, 0.002064008, 0.001979402, 
    0.001911182, 0.001665532, 0.001465833, 0.001501403, 0.001610885, 
    0.002024718, 0.002015737, 0.001845045, 0.001926426, 0.001988286, 
    0.001946039, 0.001930319, 0.001990384, 0.001836542, 0.001759263, 
    0.002206074, 0.001994391, 0.002081953, 0.002329496, 0.002397778, 
    0.002425356, 0.002488217, 0.002531897, 0.002580645, 0.002537794, 
    0.002317384, 0.002059717, 0.001734466, 0.0016518, 0.001265912, 
    0.001122719, 0.001171784, 0.00115821, 0.001132922, 0.001123068, 
    0.001104471, 0.001057233, 0.00104555, 0.001109382, 0.001156113, 
    0.001168161, 0.001172484, 0.001169194, 0.001148865, 0.001119046, 
    0.001164217, 0.001212363, 0.001226874, 0.001207944, 0.001246884, 
    0.001301578, 0.001335036, 0.00140378, 0.001733719, 0.001987603, 
    0.00200024, 0.002332133, 0.002853286, 0.003087158, 0.003232528, 
    0.003078511, 0.002899713, 0.002667492, 0.002176859, 0.002370344, 
    0.002610162, 0.002583412, 0.002582076, 0.002509788, 0.002450421, 
    0.001667393, 0.001220804, 0.0008340413, 0.0007605129, 0.0007428699, 
    0.0007634517, 0.0005730027, 0.0003954442, 0.0003504623, 0.0004442083, 
    0.0008035842, 0.001150674, 0.001259488, 0.001289435, 0.001509352, 
    0.00202974,
  0.00175791, 0.001856314, 0.001942129, 0.001937312, 0.001770929, 
    0.001738567, 0.001539392, 0.001525261, 0.001440321, 0.001566413, 
    0.001645615, 0.001617163, 0.001683715, 0.001859286, 0.001916092, 
    0.002047922, 0.002115221, 0.00211433, 0.002213639, 0.00221356, 
    0.002391436, 0.00246614, 0.002275486, 0.00195699, 0.001968864, 
    0.001814878, 0.002024304, 0.002018535, 0.002084433, 0.002224241, 
    0.002286898, 0.002200162, 0.002234875, 0.002237498, 0.002217837, 
    0.002110023, 0.001859652, 0.001591352, 0.001062001, 0.001001681, 
    0.001166174, 0.001170323, 0.001133209, 0.001069169, 0.001075432, 
    0.001088767, 0.001079341, 0.00106669, 0.001064862, 0.001055039, 
    0.001060904, 0.001087718, 0.001130395, 0.001153426, 0.001179208, 
    0.001185692, 0.001180097, 0.001192193, 0.001203637, 0.001202857, 
    0.001224824, 0.001314357, 0.001478675, 0.001570291, 0.001673622, 
    0.00166817, 0.002234065, 0.002682308, 0.002794985, 0.002792201, 
    0.002650185, 0.002386828, 0.002291365, 0.002186063, 0.002228375, 
    0.002179912, 0.002070033, 0.002015674, 0.002036274, 0.002055554, 
    0.001728556, 0.001803054, 0.0009620399, 0.0008601565, 0.000805812, 
    0.0006345483, 0.0002857898, -5.470403e-005, -0.0001919698, -9.88273e-005, 
    0.0003054822, 0.0008115796, 0.001096586, 0.001120793, 0.001189045, 
    0.001322797,
  0.001617308, 0.001252211, 0.001508922, 0.001488307, 0.001520779, 
    0.001537295, 0.001372531, 0.001233215, 0.001339423, 0.001356319, 
    0.001385025, 0.001329918, 0.001386073, 0.001648906, 0.00174564, 
    0.001715806, 0.001909036, 0.002162619, 0.002267824, 0.00230079, 
    0.002372204, 0.002388258, 0.002330639, 0.002234637, 0.002292127, 
    0.002360379, 0.002386335, 0.002244969, 0.002186175, 0.002154639, 
    0.002288535, 0.002297246, 0.002203833, 0.002101122, 0.002009347, 
    0.00194871, 0.001754986, 0.001406085, 0.000921573, 0.0008948217, 
    0.001198106, 0.001339219, 0.001575777, 0.001138708, 0.001064417, 
    0.001020532, 0.001032151, 0.001042005, 0.001054976, 0.001057058, 
    0.001096667, 0.001168987, 0.001228512, 0.001272238, 0.00130088, 
    0.001303185, 0.001260683, 0.001223871, 0.001181909, 0.001161135, 
    0.001148068, 0.00141969, 0.001534275, 0.00162435, 0.001699706, 
    0.001877581, 0.002091268, 0.002204866, 0.002160759, 0.002178672, 
    0.002193804, 0.00218263, 0.00212765, 0.002078076, 0.002140956, 
    0.0007504351, 0.001588, 0.001671145, 0.001727332, 0.001755703, 
    0.001642772, 0.0009696372, 0.0007267524, 0.0005845437, 0.0005030683, 
    0.0004943106, 0.0003180713, -1.191534e-005, -0.0002388745, -0.0001549353, 
    0.0001861779, 0.0005775811, 0.0008389037, 0.0009741029, 0.001348737, 
    0.001586217,
  0.0008563087, 0.0009093969, 0.0008977465, 0.001226302, 0.001346845, 
    0.001462081, 0.001325547, 0.001142378, 0.001295045, 0.00135279, 
    0.001291183, 0.001419373, 0.001552998, 0.001582578, 0.001785584, 
    0.00185134, 0.001949933, 0.002080031, 0.002336522, 0.002455984, 
    0.002582188, 0.002613659, 0.002632573, 0.002648293, 0.002559935, 
    0.002477824, 0.002501618, 0.002470925, 0.00237629, 0.002269733, 
    0.002240629, 0.002209825, 0.002191928, 0.002162158, 0.00206803, 
    0.001861306, 0.001615735, 0.001356335, 0.0007884237, 0.0007688254, 
    0.000958337, 0.001104058, 0.001690709, 0.001642216, 0.001065403, 
    0.001002794, 0.001031356, 0.00114052, 0.001255025, 0.001343716, 
    0.001422967, 0.001416688, 0.001378526, 0.001377603, 0.001400523, 
    0.001251687, 0.001208485, 0.001180844, 0.001189571, 0.001192877, 
    0.001462654, 0.001491455, 0.001601415, 0.001688865, 0.001786348, 
    0.001944339, 0.002036908, 0.001911802, 0.001917079, 0.001976175, 
    0.001920306, 0.001772345, 0.0006902744, 0.0004057619, 0.0003075486, 
    0.0003943164, 0.00127378, 0.001505109, 0.001494222, 0.001309067, 
    0.0006635245, 0.0005276576, 0.0003548674, 0.0001598573, 0.0001738286, 
    0.0003791703, 0.0004317188, 0.000346364, 0.000235022, 0.0002708323, 
    0.0004124218, 0.0005504498, 0.0006605675, 0.0007577632, 0.0008965544, 
    0.001155651,
  0.0005283407, 0.000575786, 0.0008193855, 0.001013602, 0.001128265, 
    0.001008546, 0.001203255, 0.001180032, 0.001285174, 0.001362502, 
    0.001431961, 0.001508461, 0.001588109, 0.001674449, 0.001825781, 
    0.002012287, 0.002189862, 0.002434558, 0.002633669, 0.002708215, 
    0.002649136, 0.002605886, 0.00261776, 0.002529179, 0.00242313, 
    0.002458639, 0.002359664, 0.002275947, 0.00225468, 0.002239039, 
    0.00218689, 0.002150475, 0.002194805, 0.002182551, 0.002072893, 
    0.001882683, 0.001709719, 0.001569546, 0.00144285, 0.001437653, 
    0.001524438, 0.001570102, 0.001713916, 0.001683924, 0.001675643, 
    0.001547946, 0.001563379, 0.001050573, 0.001099973, 0.001194593, 
    0.001253007, 0.001249955, 0.001411506, 0.001408343, 0.001432836, 
    0.001504919, 0.001558865, 0.001770739, 0.001809411, 0.001752875, 
    0.001719527, 0.001735533, 0.001755973, 0.001848463, 0.001956371, 
    0.002026275, 0.001946039, 0.001714917, 0.001647683, 0.001643916, 
    0.001500103, 0.0008745082, 0.0005870867, 0.0003523396, 0.0002364044, 
    0.0002516787, 0.0009237495, 0.001014285, 0.0004296671, 0.0003861471, 
    0.0003905499, 0.0003505759, 0.000291368, 0.0001844768, 0.0001299107, 
    0.0001157499, 0.0002100673, 0.0003353651, 0.0004398241, 0.0005405792, 
    0.0005938262, 0.0005057068, 0.0003435505, 0.0003015087, 0.0004410795, 
    0.0005156407,
  0.0002749022, 0.000331725, 0.0004345146, 0.0007710988, 0.0008778623, 
    0.0009863749, 0.0008272696, 0.001193083, 0.001293028, 0.001386949, 
    0.001465182, 0.001538695, 0.001637877, 0.001776191, 0.00192541, 
    0.002076234, 0.002256637, 0.002448245, 0.002572286, 0.002673121, 
    0.00269976, 0.002709932, 0.002645098, 0.002542721, 0.002479796, 
    0.002349094, 0.00219142, 0.002031363, 0.001950602, 0.002026306, 
    0.001936328, 0.002067554, 0.002038863, 0.001951761, 0.001906509, 
    0.001810062, 0.001489851, 0.001417022, 0.001319906, 0.001306857, 
    0.001519335, 0.001374933, 0.001403114, 0.001308605, 0.001145701, 
    0.001087941, 0.001186074, 0.001258045, 0.001194864, 0.001309559, 
    0.001295015, 0.001042387, 0.001331653, 0.001390192, 0.001492934, 
    0.001590288, 0.00165064, 0.001689455, 0.001705858, 0.001738139, 
    0.001791244, 0.00187895, 0.001854456, 0.001780689, 0.001776684, 
    0.001736502, 0.001671826, 0.001592832, 0.001524311, 0.001337501, 
    0.001308525, 0.00132458, 0.001174471, 0.0009425213, 0.0004480728, 
    0.000408384, 0.0005123666, 0.0008142041, 0.0007686503, 0.0006541461, 
    0.0004869509, 0.0004614559, 0.0005403566, 0.0003860521, 0.0003349986, 
    0.0002766496, 0.0001880215, 0.0001843823, 0.0002460531, 0.0004586587, 
    0.0005878657, 0.0006751758, 0.0004814197, 0.000206857, 9.254366e-005, 
    0.0001308969,
  0.0003148611, 0.0003182627, 0.0003055949, 0.0002597547, 0.0002314621, 
    0.00074794, 0.00100664, 0.00123104, 0.001359753, 0.001362058, 
    0.001308256, 0.0009345263, 0.0009312681, 0.0009983745, 0.001644235, 
    0.001783789, 0.00197117, 0.002106973, 0.002267382, 0.002463695, 
    0.002585972, 0.002595478, 0.00252829, 0.002374257, 0.002173334, 
    0.001868126, 0.001733324, 0.00179002, 0.001828564, 0.001845253, 
    0.001786713, 0.001693937, 0.001594309, 0.001542987, 0.001311641, 
    0.001279486, 0.001350726, 0.001189237, 0.001153665, 0.00103115, 
    0.0008149678, 0.0007505622, 0.0006383308, 0.0005751816, 0.0006858399, 
    0.0007374017, 0.0007329206, 0.0007577315, 0.0007713209, 0.0005034343, 
    0.0004143608, 0.0004962026, 0.0005981335, 0.001057645, 0.001203081, 
    0.001283095, 0.001273796, 0.001221693, 0.001223092, 0.001197295, 
    0.001108953, 0.001105155, 0.001106283, 0.001208215, 0.001347627, 
    0.001442962, 0.001611269, 0.001481013, 0.001371516, 0.0007123677, 
    0.0010785, 0.001007992, 0.0009666495, 0.0006428612, 0.0008928985, 
    0.0005813963, 0.0008008368, 0.0007568412, 0.0006185737, 0.0005523572, 
    0.0005418509, 0.0005375112, 0.0005870871, 0.0006076379, 0.0006327196, 
    0.000594191, 0.0005003177, 0.0003840807, 0.0003031937, 0.0003220921, 
    0.0003897713, 0.0004606456, 0.0004074466, 0.0003867839, 0.0003576013, 
    0.0003378759,
  0.0006001364, 0.0006088465, 0.0005629114, 0.0004967265, 0.0004368196, 
    0.000517135, 0.0007208874, 0.000856881, 0.0008626035, 0.0007863576, 
    0.0006681648, 0.0005975133, 0.0005503537, 0.0005133834, 0.0004853455, 
    0.0007572388, 0.0005693485, 0.0006355015, 0.0007559503, 0.001513137, 
    0.001919036, 0.002047607, 0.002112139, 0.002135759, 0.002084991, 
    0.002009078, 0.001896927, 0.001853201, 0.001852056, 0.001739204, 
    0.001709037, 0.001503329, 0.001280185, 0.001081583, 0.0009192042, 
    0.000615872, 0.0005903137, 0.0006201961, 0.0008936459, 0.000837808, 
    0.0005684108, 0.000466113, 0.0003658659, 0.0002778894, 0.0002327967, 
    0.0002264548, 0.000241173, 0.0002463546, 0.0002269314, 0.0001854624, 
    0.0001351084, 0.000110806, 0.0001334553, 0.0001879102, 0.0002373583, 
    0.0002650148, 0.0002626146, 0.0002422857, 0.0002324786, 0.0002428736, 
    0.0002958663, 0.0003757202, 0.0004921961, 0.00097838, 0.001171261, 
    0.001285383, 0.001384311, 0.00134262, 0.001224412, 0.0006478676, 
    0.0008508731, 0.0007800786, 0.0006580399, 0.0007918249, 0.0008301949, 
    0.0009324602, 0.0006550048, 0.0005000953, 0.0004423505, 0.0004190016, 
    0.0004430022, 0.0006156815, 0.0005323614, 0.000571446, 0.0005845594, 
    0.0005929837, 0.0006017573, 0.0006171747, 0.0006087667, 0.0005690937, 
    0.0006294453, 0.0003512905, 0.0003607161, 0.0004130728, 0.0004439875, 
    0.000517501,
  0.000426027, 0.0004758402, 0.0005589691, 0.0006410806, 0.0006375518, 
    0.0005872608, 0.000548749, 0.0004468807, 0.0003597941, 0.0002714838, 
    0.0002159481, 0.0001724446, 0.0001374607, 9.815348e-005, 7.704552e-005, 
    8.519948e-005, 9.975885e-005, 0.0001427059, 0.0002032323, 0.0002871717, 
    0.0003786292, 0.0004612808, 0.000534921, 0.0005844003, 0.0006228974, 
    0.001033089, 0.001025714, 0.001104137, 0.001052384, 0.0009150556, 
    0.000796291, 0.0004643011, 0.0003583473, 0.0002797807, 0.0002030891, 
    0.0001831418, 0.0001882121, 0.0002098128, 0.000235721, 0.0002457823, 
    0.000234958, 0.0002061254, 0.0001740183, 0.0001486663, 0.0001350448, 
    0.0001403219, 0.0001560415, 0.0001761641, 0.0001905011, 0.0001927738, 
    0.0001879737, 0.0001827762, 0.0001747336, 0.0001663889, 0.0001569951, 
    0.0001457259, 0.0001342183, 0.0001232671, 0.0001168614, 0.0001212163, 
    0.000142833, 0.0001791681, 0.0002371354, 0.000302033, 0.0003776753, 
    0.0006029662, 0.000695806, 0.0007403586, 0.0008000107, 0.0008490295, 
    0.0008174949, 0.0005600657, 0.0005422961, 0.0005303281, 0.0005364306, 
    0.0003188336, 0.000294531, 0.00027897, 0.000429508, 0.0004736469, 
    0.0005133196, 0.0005328221, 0.0005341896, 0.0005308198, 0.0005307086, 
    0.0005520709, 0.000592618, 0.0006412072, 0.0006736957, 0.000651062, 
    0.0005911556, 0.0005535488, 0.0003556614, 0.0002726917, 0.0002619154, 
    0.0003722711,
  0.0001809483, 0.0001452651, 0.000136825, 0.0001321521, 0.0002667313, 
    0.0002524264, 0.00023828, 0.0001049086, 0.00011346, 0.0001197702, 
    0.0001105512, 0.0001045908, 9.961566e-005, 9.977468e-005, 0.0001076267, 
    0.0001103922, 0.0001166072, 0.0001215662, 0.0001234259, 0.0001195318, 
    0.0001192139, 0.0001163527, 0.0001156055, 0.000113603, 0.0001336776, 
    0.0002703872, 0.0002770629, 0.0002201281, 0.0002279168, 0.0002170769, 
    0.0001982097, 0.0001747813, 0.0001451219, 0.0001126016, 8.715456e-005, 
    7.346924e-005, 7.612375e-005, 8.923677e-005, 0.0001148744, 0.0001444225, 
    0.0001689638, 0.0001870198, 0.0001934415, 0.0001917724, 0.0001869088, 
    0.0001773085, 0.0001691387, 0.0001659915, 0.0001639731, 0.0001656737, 
    0.00017165, 0.0001857325, 0.0001980509, 0.0002114023, 0.0002186978, 
    0.0002262001, 0.0002291724, 0.0002242769, 0.000220017, 0.0002090817, 
    0.0002035345, 0.0002036458, 0.000203884, 0.0002160755, 0.0002383755, 
    0.0002668584, 0.0002995376, 0.0003245717, 0.000344869, 0.0003493989, 
    0.0003449484, 0.000519217, 0.0006774156, 0.000383175, 0.0003800758, 
    0.0003911546, 0.0004018191, 0.0004204158, 0.0004411105, 0.0004653179, 
    0.0004859333, 0.0005098865, 0.0005289124, 0.0005440284, 0.0005619891, 
    0.0005840665, 0.0006023132, 0.0006107374, 0.0005994204, 0.0005657719, 
    0.0005123822, 0.0004546209, 0.0003222192, 0.000280655, 0.0002467996, 
    0.0002140566,
  0.0001867178, 0.0001750197, 0.0001680737, 0.000159872, 0.0001604601, 
    0.0001621291, 0.0001622562, 0.0001609689, 0.0001607782, 0.0001599994, 
    0.0001617477, 0.0001657212, 0.0001700285, 0.0001720632, 0.0001726833, 
    0.0001695838, 0.0001629717, 0.0001551039, 0.0001431194, 0.0001313095, 
    0.0001181646, 0.0001051312, 9.284448e-005, 8.252915e-005, 7.784017e-005, 
    7.769722e-005, 8.07012e-005, 8.891872e-005, 9.502214e-005, 0.0001029854, 
    0.0001114414, 0.000117386, 0.0001222179, 0.0001271134, 0.0001343137, 
    0.0001368884, 0.0001398132, 0.0001447881, 0.0001503194, 0.0001525604, 
    0.0001546904, 0.0001538161, 0.0001554694, 0.0001573926, 0.0001582508, 
    0.0001586482, 0.0001580759, 0.0001606189, 0.0001664364, 0.0001719994, 
    0.0001812503, 0.0001929486, 0.0002037252, 0.0002154235, 0.0002242611, 
    0.0002315091, 0.0002352761, 0.0002391383, 0.0002385026, 0.0002379939, 
    0.0002369131, 0.0002314453, 0.0002289498, 0.0002273447, 0.0002256597, 
    0.0002255167, 0.0002261684, 0.0002292201, 0.000236023, 0.0002460685, 
    0.0002580211, 0.0002710705, 0.0002842948, 0.0002960407, 0.0003157819, 
    0.0003374782, 0.0003628458, 0.000390566, 0.0004201299, 0.0004454975, 
    0.0004666531, 0.0004850591, 0.0004930701, 0.0004943416, 0.0004876817, 
    0.0004748865, 0.0004391398, 0.0004047598, 0.0003694422, 0.0003373667, 
    0.0003028279, 0.0002724852, 0.0002505507, 0.0002342905, 0.0002181258, 
    0.0002020723,
  0.0002697194, 0.0002659047, 0.0002636635, 0.0002603736, 0.0002575284, 
    0.0002536499, 0.0002499307, 0.0002449399, 0.0002399806, 0.0002352919, 
    0.0002317631, 0.000225628, 0.0002189046, 0.0002124673, 0.0002053624, 
    0.0001975421, 0.0001897537, 0.0001831895, 0.0001782463, 0.0001737161, 
    0.0001690113, 0.0001630192, 0.0001594431, 0.0001572177, 0.0001551195, 
    0.0001536414, 0.0001513208, 0.0001496361, 0.0001486982, 0.0001486344, 
    0.0001505737, 0.0001524652, 0.0001548335, 0.000158807, 0.0001631305, 
    0.0001682963, 0.0001734779, 0.0001783099, 0.0001832689, 0.0001872424, 
    0.000192154, 0.0001955871, 0.0001998947, 0.000201659, 0.0002043608, 
    0.0002088591, 0.0002128009, 0.0002162503, 0.0002195244, 0.0002221151, 
    0.0002231644, 0.0002229577, 0.0002214159, 0.0002219405, 0.0002210503, 
    0.0002213998, 0.0002215111, 0.0002196676, 0.0002200648, 0.0002196673, 
    0.0002219405, 0.0002252941, 0.0002273605, 0.0002291724, 0.00022771, 
    0.0002279168, 0.000228171, 0.0002309049, 0.0002322719, 0.0002362456, 
    0.0002412365, 0.0002449399, 0.0002456869, 0.0002493109, 0.0002521083, 
    0.0002526646, 0.0002541109, 0.0002573533, 0.0002616292, 0.0002664609, 
    0.0002695764, 0.0002725963, 0.0002724375, 0.00027444, 0.0002752985, 
    0.0002774759, 0.0002772217, 0.000277333, 0.0002787793, 0.0002811796, 
    0.0002818787, 0.0002793833, 0.0002772377, 0.0002790496, 0.000277492, 
    0.0002750759,
  8.377514e-006, 7.900679e-006, 7.455632e-006, 6.962902e-006, 6.533746e-006, 
    6.168173e-006, 5.707228e-006, 5.357548e-006, 5.08734e-006, 4.769448e-006, 
    4.546922e-006, 4.308505e-006, 4.213137e-006, 4.070082e-006, 
    3.911138e-006, 3.81577e-006, 3.783982e-006, 3.656824e-006, 3.752192e-006, 
    3.783982e-006, 3.768087e-006, 3.879349e-006, 3.879349e-006, 
    4.006505e-006, 4.117767e-006, 4.292608e-006, 4.37208e-006, 4.562815e-006, 
    4.817128e-006, 5.087336e-006, 5.278071e-006, 5.580067e-006, 
    5.850276e-006, 6.231746e-006, 6.597322e-006, 6.994688e-006, 
    7.487421e-006, 7.932469e-006, 8.377521e-006, 8.854355e-006, 
    9.251724e-006, 9.82392e-006, 1.012592e-005, 1.049149e-005, 1.090475e-005, 
    1.119085e-005, 1.131801e-005, 1.152464e-005, 1.16518e-005, 1.176306e-005, 
    1.176306e-005, 1.176306e-005, 1.162001e-005, 1.142927e-005, 
    1.142928e-005, 1.131801e-005, 1.128623e-005, 1.112728e-005, 
    1.109549e-005, 1.109549e-005, 1.119085e-005, 1.119085e-005, 1.13498e-005, 
    1.150874e-005, 1.157233e-005, 1.16677e-005, 1.176306e-005, 1.185843e-005, 
    1.19379e-005, 1.206506e-005, 1.203327e-005, 1.200148e-005, 1.198558e-005, 
    1.176306e-005, 1.190611e-005, 1.192201e-005, 1.174717e-005, 
    1.179485e-005, 1.184253e-005, 1.189022e-005, 1.185842e-005, 
    1.187432e-005, 1.176306e-005, 1.179485e-005, 1.173127e-005, 
    1.168359e-005, 1.155643e-005, 1.141338e-005, 1.122264e-005, 
    1.107959e-005, 1.084118e-005, 1.053918e-005, 1.011003e-005, 
    9.712661e-006, 9.235824e-006, 8.743093e-006,
  9.680873e-006, 8.568253e-006, 7.471524e-006, 6.660905e-006, 5.99333e-006, 
    5.627755e-006, 5.246285e-006, 4.801235e-006, 4.467449e-006, 
    4.149558e-006, 3.942927e-006, 3.593246e-006, 3.418407e-006, 
    3.132303e-006, 3.084619e-006, 2.87799e-006, 2.814412e-006, 2.893886e-006, 
    2.862096e-006, 2.941569e-006, 2.973357e-006, 3.021042e-006, 
    3.068726e-006, 3.195883e-006, 3.116411e-006, 3.338935e-006, 
    3.513774e-006, 3.625036e-006, 3.768087e-006, 3.847559e-006, 
    4.054189e-006, 4.356185e-006, 4.801235e-006, 5.341652e-006, 
    6.104594e-006, 7.05827e-006, 8.234465e-006, 9.649082e-006, 1.13657e-005, 
    1.300284e-005, 1.463998e-005, 1.622945e-005, 1.742153e-005, 
    1.856594e-005, 1.910635e-005, 1.918583e-005, 1.964677e-005, 
    1.975803e-005, 1.980571e-005, 1.977392e-005, 1.990108e-005, 2.04256e-005, 
    2.017129e-005, 2.036202e-005, 1.907456e-005, 1.918584e-005, 
    1.802553e-005, 1.651554e-005, 1.502145e-005, 1.390883e-005, 
    1.325715e-005, 1.295516e-005, 1.308232e-005, 1.357505e-005, 
    1.468766e-005, 1.629302e-005, 1.791426e-005, 1.918582e-005, 
    1.994877e-005, 2.037792e-005, 2.037792e-005, 2.012361e-005, 
    1.978982e-005, 1.940835e-005, 1.910636e-005, 1.931299e-005, 
    1.977393e-005, 2.039381e-005, 2.026666e-005, 2.115675e-005, 
    2.263494e-005, 2.276211e-005, 2.486019e-005, 2.546419e-005, 
    2.713313e-005, 2.751459e-005, 2.767353e-005, 2.713312e-005, 2.59728e-005, 
    2.433568e-005, 2.225348e-005, 1.993287e-005, 1.750101e-005, 
    1.524397e-005, 1.306642e-005, 1.115907e-005,
  6.374801e-006, 5.119129e-006, 4.197243e-006, 3.736299e-006, 3.243569e-006, 
    3.227675e-006, 3.243566e-006, 3.338934e-006, 3.46609e-006, 3.370723e-006, 
    3.243566e-006, 3.052831e-006, 2.846202e-006, 2.846202e-006, 
    3.068725e-006, 3.259463e-006, 3.736299e-006, 3.942929e-006, 
    4.022401e-006, 3.720404e-006, 3.291249e-006, 2.671361e-006, 
    2.194524e-006, 1.924318e-006, 1.797163e-006, 1.876635e-006, 
    2.083264e-006, 2.337577e-006, 2.591891e-006, 2.893888e-006, 
    3.116411e-006, 3.164094e-006, 3.164093e-006, 3.307144e-006, 
    3.656824e-006, 4.578712e-006, 6.072805e-006, 8.091414e-006, 
    1.071402e-005, 1.384525e-005, 1.669038e-005, 1.86613e-005, 1.971035e-005, 
    1.902688e-005, 1.758048e-005, 1.624533e-005, 1.51645e-005, 1.510092e-005, 
    1.589565e-005, 1.754869e-005, 1.993287e-005, 2.36681e-005, 2.821394e-005, 
    3.2728e-005, 3.647913e-005, 3.841828e-005, 3.749637e-005, 3.414261e-005, 
    2.9565e-005, 2.455819e-005, 2.006003e-005, 1.635659e-005, 1.405188e-005, 
    1.284391e-005, 1.327304e-005, 1.494199e-005, 1.748512e-005, 
    2.028257e-005, 2.220581e-005, 2.315947e-005, 2.307999e-005, 
    2.238063e-005, 2.149054e-005, 2.093423e-005, 2.099781e-005, 
    2.199916e-005, 2.368399e-005, 2.733974e-005, 3.196507e-005, 
    3.705133e-005, 4.331379e-005, 4.959214e-005, 5.471017e-005, 
    5.774606e-005, 5.865203e-005, 5.707849e-005, 5.305714e-005, 
    4.865434e-005, 4.310717e-005, 3.68288e-005, 3.132931e-005, 2.54324e-005, 
    1.980572e-005, 1.506913e-005, 1.117496e-005, 8.377519e-006,
  1.147695e-005, 9.315296e-006, 7.598683e-006, 6.231747e-006, 5.373443e-006, 
    4.833025e-006, 4.626394e-006, 4.896602e-006, 4.944286e-006, 
    4.721763e-006, 4.133663e-006, 3.418406e-006, 2.87799e-006, 2.639572e-006, 
    2.719045e-006, 3.243569e-006, 4.292615e-006, 5.595968e-006, 
    6.692695e-006, 7.042374e-006, 6.390695e-006, 4.864818e-006, 
    3.021047e-006, 1.670007e-006, 1.145483e-006, 1.081904e-006, 
    1.368006e-006, 1.813054e-006, 2.464732e-006, 2.973357e-006, 
    3.354829e-006, 3.720404e-006, 3.799878e-006, 3.863455e-006, 
    4.038298e-006, 4.642292e-006, 5.754911e-006, 7.201321e-006, 
    8.965613e-006, 1.131801e-005, 1.424261e-005, 1.710363e-005, 
    1.963088e-005, 2.090244e-005, 2.177664e-005, 2.409725e-005, 
    2.908815e-005, 2.834111e-005, 3.345916e-005, 2.708544e-005, 
    3.002591e-005, 3.237833e-005, 3.506453e-005, 3.651093e-005, 
    3.728976e-005, 3.810036e-005, 4.134286e-005, 3.393601e-005, 
    2.924711e-005, 2.352508e-005, 1.756458e-005, 1.436978e-005, 
    1.311411e-005, 1.414726e-005, 1.643607e-005, 1.907455e-005, 2.1268e-005, 
    2.285746e-005, 2.355684e-005, 2.486019e-005, 2.670394e-005, 
    2.923119e-005, 3.239422e-005, 3.528705e-005, 3.759175e-005, 
    3.911764e-005, 4.037331e-005, 4.197864e-005, 4.498271e-005, 
    5.002129e-005, 6.424695e-005, 6.876102e-005, 7.395849e-005, 
    7.677186e-005, 7.948984e-005, 8.168328e-005, 8.252569e-005, 
    8.297077e-005, 8.626094e-005, 6.820471e-005, 5.951036e-005, 
    4.828878e-005, 3.597051e-005, 2.622712e-005, 1.912225e-005, 1.454461e-005,
  2.57026e-005, 2.48602e-005, 2.236474e-005, 1.805731e-005, 1.414724e-005, 
    1.228758e-005, 1.285979e-005, 1.45764e-005, 1.686522e-005, 1.791426e-005, 
    1.63248e-005, 1.289158e-005, 8.806674e-006, 6.215852e-006, 5.087344e-006, 
    4.896605e-006, 5.230393e-006, 5.580072e-006, 5.278074e-006, 
    5.055554e-006, 7.34437e-006, 9.871612e-006, 9.903397e-006, 8.266255e-006, 
    6.470171e-006, 4.880712e-006, 3.847563e-006, 3.402516e-006, 3.67272e-006, 
    4.801232e-006, 6.295326e-006, 7.980154e-006, 9.299401e-006, 
    1.003055e-005, 1.057097e-005, 1.111139e-005, 1.160412e-005, 
    1.297105e-005, 1.484661e-005, 1.767584e-005, 2.098191e-005, 
    2.347737e-005, 2.471713e-005, 2.595691e-005, 2.770532e-005, 3.00895e-005, 
    3.703543e-005, 4.588872e-005, 5.369296e-005, 5.73805e-005, 5.636321e-005, 
    5.097489e-005, 4.565029e-005, 4.417208e-005, 4.383828e-005, 
    4.633373e-005, 5.167429e-005, 5.528235e-005, 5.539367e-005, 
    5.515519e-005, 4.986222e-005, 4.142223e-005, 3.128155e-005, 
    2.309587e-005, 1.449691e-005, 1.203318e-005, 1.503725e-005, 
    2.031424e-005, 3.199675e-005, 4.134281e-005, 3.072526e-005, 
    3.657441e-005, 4.76212e-005, 6.114747e-005, 7.445124e-005, 8.821589e-005, 
    7.221007e-005, 7.214659e-005, 7.163794e-005, 7.634275e-005, 
    9.276174e-005, 0.0001016468, 0.0001125664, 0.0001235178, 0.0001357724, 
    0.0001456111, 0.0001511107, 0.000148647, 0.0001397143, 0.0001233747, 
    0.0001013449, 6.321378e-005, 4.464893e-005, 3.353863e-005, 2.735565e-005, 
    2.619534e-005,
  0.0001359791, 0.0001279682, 7.750303e-005, 6.082961e-005, 4.836827e-005, 
    4.159717e-005, 3.975341e-005, 4.09455e-005, 4.701724e-005, 5.170613e-005, 
    5.000542e-005, 4.339327e-005, 3.271212e-005, 2.093423e-005, 
    1.362272e-005, 1.030076e-005, 9.426556e-006, 9.172247e-006, 
    1.072991e-005, 1.104781e-005, 1.16677e-005, 1.263726e-005, 1.147698e-005, 
    9.331183e-006, 9.12456e-006, 1.130213e-005, 1.533935e-005, 1.993288e-005, 
    2.45423e-005, 2.738743e-005, 2.910405e-005, 2.966035e-005, 3.145644e-005, 
    3.404725e-005, 3.682882e-005, 4.057994e-005, 4.530062e-005, 
    5.087962e-005, 5.599765e-005, 6.335683e-005, 7.332275e-005, 
    8.099983e-005, 8.804114e-005, 9.179224e-005, 0.0001056204, 0.0001169214, 
    0.0001352798, 0.0001585654, 0.0001760017, 0.0001817713, 0.0001729975, 
    0.0001604726, 0.0001486471, 0.0001357407, 0.0001203388, 0.0001050482, 
    9.134714e-005, 7.947389e-005, 7.133582e-005, 6.117928e-005, 
    4.833646e-005, 3.932416e-005, 3.547774e-005, 3.361807e-005, 
    3.724202e-005, 4.086597e-005, 4.704896e-005, 6.00348e-005, 7.424457e-005, 
    8.966232e-005, 9.554328e-005, 9.395386e-005, 9.862689e-005, 0.0001068762, 
    0.0001282226, 0.0001608859, 0.0001904179, 0.0002070756, 0.0001894803, 
    0.0001876841, 0.0002120348, 0.0002122572, 0.0002205701, 0.0002247663, 
    0.0002255291, 0.0002248457, 0.0002254338, 0.0002220641, 0.0002150387, 
    0.0002048343, 0.0001942644, 0.0001820415, 0.0001661788, 0.0001542896, 
    0.0001475821, 0.000142019,
  0.0002118121, 0.0002022754, 0.000189973, 0.0001753022, 0.0001622687, 
    0.0001519055, 0.0001463741, 0.00014639, 0.0001544485, 0.0001665443, 
    0.0001834084, 0.000192516, 0.0001817077, 0.0001522869, 0.0001170486, 
    8.902652e-005, 7.556388e-005, 7.648577e-005, 8.959873e-005, 0.0001054297, 
    0.0001111994, 0.0001024733, 8.120635e-005, 5.537772e-005, 3.644728e-005, 
    2.881791e-005, 3.062992e-005, 3.206037e-005, 2.889731e-005, 
    2.886556e-005, 4.216935e-005, 7.449894e-005, 0.0001050482, 0.0001041422, 
    0.0001222144, 0.0001477252, 0.0001952818, 0.0002380222, 0.000271067, 
    0.0002856424, 0.0002917302, 0.0002992322, 0.0003163031, 0.0003470592, 
    0.0003769253, 0.0004060601, 0.0004100337, 0.000375908, 0.0003143481, 
    0.0002579227, 0.0002062811, 0.0001802617, 0.000169056, 0.0001709951, 
    0.0001571192, 0.0001463746, 0.0001365519, 0.0001139815, 0.0001012499, 
    9.541656e-005, 9.749876e-005, 0.0001304642, 0.0001879071, 0.0002496574, 
    0.0003131721, 0.0003768777, 0.0004306808, 0.000508437, 0.0005922967, 
    0.00067862, 0.0007197076, 0.000743597, 0.0007112039, 0.0006813696, 
    0.0006337177, 0.0005915812, 0.0005241089, 0.0004805101, 0.0004514388, 
    0.0004364025, 0.0004216047, 0.0004240206, 0.0004287253, 0.000423067, 
    0.00040331, 0.000383728, 0.0003708375, 0.0003589005, 0.000346439, 
    0.0003304174, 0.0003107081, 0.0002806197, 0.0002461285, 0.0002202999, 
    0.0002096187, 0.0002113989,
  0.0003993682, 0.0004110984, 0.0004085712, 0.0004083802, 0.000395458, 
    0.0003817727, 0.0003875108, 0.0004028332, 0.0004292499, 0.0004510414, 
    0.0004825921, 0.0005141587, 0.0005210571, 0.0005157482, 0.0005173218, 
    0.0005036047, 0.0004762819, 0.0004584801, 0.0004288684, 0.0003947586, 
    0.0003589324, 0.0003248225, 0.000291873, 0.0002607356, 0.0002318393, 
    0.0001874616, 0.0001553546, 0.0001264423, 0.0001013289, 6.685359e-005, 
    4.758977e-005, 0.0001315927, 0.0001936448, 0.0002958945, 0.0003153654, 
    0.0003521454, 0.0004133396, 0.0004588615, 0.0004990592, 0.000463201, 
    0.0004808281, 0.0004565094, 0.0004521541, 0.0004904123, 0.0005522424, 
    0.0005541497, 0.0003977788, 0.0001977456, -1.935824e-005, -0.0001474528, 
    -0.0001890168, -0.0001943097, -0.0001697529, -0.0001749026, 
    -0.0001345621, -0.0001080977, -7.854938e-005, -3.216905e-005, 
    8.026906e-005, 0.000197428, 0.0003305769, 0.0003920095, 0.0004324769, 
    0.0004772996, 0.0005211367, 0.0005642266, 0.0005754801, 0.0005876394, 
    0.0006304435, 0.0006701483, 0.0007179589, 0.0007450434, 0.0007942691, 
    0.0008482947, 0.0008777156, 0.0008647614, 0.0008108469, 0.0007657541, 
    0.0007202798, 0.0006488971, 0.0006557319, 0.000679065, 0.0006914627, 
    0.0006607705, 0.000611402, 0.0005769741, 0.0005503349, 0.0005161298, 
    0.0004778873, 0.0004529647, 0.0004378171, 0.0004116705, 0.0003728083, 
    0.0003446589, 0.0003446589, 0.0003671818,
  0.0005311026, 0.0005593154, 0.0006142788, 0.0006427619, 0.0006823394, 
    0.0007200253, 0.0007115059, 0.0006832927, 0.0006652209, 0.0006632658, 
    0.0006244513, 0.0006176962, 0.0006759656, 0.0007376208, 0.0008017553, 
    0.0008674476, 0.000870086, 0.000913637, 0.0009302946, 0.0008151701, 
    0.0007094714, 0.0006192856, 0.0005372697, 0.0004843246, 0.0004773152, 
    0.0004850875, 0.0004626603, 0.0004794452, 0.000493814, 0.0004729126, 
    0.0004261828, 0.0003654652, 0.0003094368, 0.0002702726, 0.0002548075, 
    0.0002902206, 0.0003544982, 0.0003717437, 0.0003791347, 0.0004318568, 
    0.0005227898, 0.0006164247, 0.0007288151, 0.0008116898, 0.000798211, 
    0.0007628612, 0.0006930206, 0.0004401854, 0.000128, 1.29235e-005, 
    -1.702178e-005, -3.358396e-005, -5.032099e-005, -9.48098e-005, 
    -0.0001403638, -0.0001854089, -0.0001686083, -5.340436e-005, 
    8.036406e-005, 0.0001917377, 0.0002798571, 0.0003377611, 0.0003814555, 
    0.0004261509, 0.0004558577, 0.0004893001, 0.0005400989, 0.0005672628, 
    0.0005667384, 0.0005907551, 0.0006209388, 0.0006318109, 0.0006468629, 
    0.0006666514, 0.0006801935, 0.0006575121, 0.0005994013, 0.0005886727, 
    0.0006016425, 0.0005943789, 0.0005864792, 0.0006051715, 0.0005000131, 
    0.0004986459, 0.0005303398, 0.0005977484, 0.0006535542, 0.0006795577, 
    0.0006629318, 0.0006389628, 0.0006312701, 0.0006130708, 0.0006056322, 
    0.0005610955, 0.0005076423, 0.0005118385,
  0.0005676916, 0.0006119262, 0.0006229572, 0.0006059818, 0.0005835546, 
    0.0005762589, 0.00059751, 0.0006155346, 0.0005989724, 0.0005941088, 
    0.0006017061, 0.0005953326, 0.0006021352, 0.0006194285, 0.0006545556, 
    0.0006973597, 0.0007657064, 0.000850965, 0.0008922589, 0.0008178407, 
    0.0006783975, 0.0006134363, 0.0006064747, 0.0005849851, 0.0005660707, 
    0.0005788498, 0.0005933931, 0.0005891179, 0.0005734935, 0.0005686933, 
    0.0005460435, 0.0004937029, 0.0004497541, 0.0004354487, 0.0004481007, 
    0.0005056551, 0.0005566929, 0.0005713317, 0.0005255709, 0.0005277647, 
    0.0006320332, 0.0008194768, 0.0009939522, 0.001018779, 0.0009418335, 
    0.000886838, 0.0008114502, 0.0006873296, 0.0005030003, 0.0003718385, 
    0.0002816999, 0.0002145297, 0.0001605204, 0.0001372187, 0.0001221024, 
    0.0001169848, 0.0001596776, 0.0002272935, 0.0003019022, 0.0003439118, 
    0.0003691525, 0.0003713616, 0.0003867797, 0.0004100334, 0.00042383, 
    0.0004331442, 0.0004630578, 0.0004962618, 0.0005163201, 0.0005226941, 
    0.0005420856, 0.0005743518, 0.0005772761, 0.0005669449, 0.0005611903, 
    0.0005673249, 0.00060126, 0.0006684, 0.0006402347, 0.000561906, 
    0.0005730637, 0.0006034225, 0.0006493423, 0.0004915567, 0.0004798584, 
    0.0005370153, 0.0006039632, 0.0006580527, 0.0006836271, 0.0006762675, 
    0.0006711814, 0.0006519808, 0.0006216858, 0.0005617633, 0.000506911, 
    0.0005140475,
  0.0005457415, 0.0005575353, 0.0006041066, 0.0006415064, 0.0006484841, 
    0.0006582912, 0.0006958656, 0.000729928, 0.0007430252, 0.0007548349, 
    0.0007658021, 0.0007638948, 0.0007570123, 0.0007343465, 0.000727671, 
    0.0007657069, 0.0008674636, 0.0009689503, 0.0009662802, 0.0009002225, 
    0.0008787648, 0.0009243502, 0.0009605102, 0.0009397673, 0.0009013023, 
    0.0009089955, 0.0009490815, 0.0009625759, 0.0009323922, 0.0008716746, 
    0.0007859077, 0.0006824974, 0.000621208, 0.0006303475, 0.0006790799, 
    0.0007201042, 0.0007170364, 0.0006583058, 0.0006086663, 0.0006559221, 
    0.0008073174, 0.0009727166, 0.001034817, 0.001014805, 0.001014996, 
    0.0009911377, 0.0009154794, 0.0008167434, 0.0006526476, 0.0005317852, 
    0.0005071168, 0.0004870896, 0.0004736586, 0.0004791263, 0.000478093, 
    0.0004601958, 0.0004760111, 0.00051837, 0.0005472666, 0.0005523046, 
    0.0005323095, 0.0004968802, 0.0004585902, 0.0004634704, 0.0004744697, 
    0.0004627071, 0.0004573348, 0.0004723547, 0.0004844349, 0.0004595281, 
    0.0004370846, 0.0004522959, 0.0004643602, 0.000460784, 0.0004828298, 
    0.0006081103, 0.0006940058, 0.0006821172, 0.0006657764, 0.0006711488, 
    0.0006244658, 0.0006003859, 0.0006896667, 0.0006313971, 0.0005817742, 
    0.0005817588, 0.0006254367, 0.0006691471, 0.0006885703, 0.0006892378, 
    0.000657957, 0.0006271536, 0.0006117362, 0.0005683277, 0.0005330418, 
    0.0005242522,
  0.0006951969, 0.0007340754, 0.0007859394, 0.000828966, 0.0008487068, 
    0.0008978057, 0.0009899619, 0.001078924, 0.00112691, 0.001161513, 
    0.001186928, 0.001198658, 0.001183352, 0.001127991, 0.001070452, 
    0.001028618, 0.001059835, 0.001175293, 0.001199771, 0.001319298, 
    0.001602889, 0.001744732, 0.001661174, 0.001479864, 0.001348718, 
    0.001281993, 0.00123264, 0.001176071, 0.001106962, 0.001015425, 
    0.0009142398, 0.0008467515, 0.0008061407, 0.000790548, 0.0007961113, 
    0.0007734299, 0.0006917636, 0.000650676, 0.000681893, 0.0007385258, 
    0.0009184675, 0.001098235, 0.001119375, 0.001109568, 0.001167822, 
    0.001061503, 0.0009574099, 0.0008762521, 0.0008356413, 0.0007804395, 
    0.0007908186, 0.0008338452, 0.0008499306, 0.0008185543, 0.0007627807, 
    0.0007415297, 0.0007476327, 0.0007563112, 0.0007479824, 0.0007326286, 
    0.0007033828, 0.0006218748, 0.000565799, 0.0005404316, 0.0005256333, 
    0.0005137445, 0.0005104863, 0.0004933672, 0.000495418, 0.0005033016, 
    0.0004979135, 0.0004917784, 0.0004960853, 0.0004891874, 0.0005254587, 
    0.0006059487, 0.0006308244, 0.0005736046, 0.0006292039, 0.0006839279, 
    0.0006538713, 0.0006360216, 0.0006821635, 0.0006480222, 0.0006330335, 
    0.0006356407, 0.0006877747, 0.0007399884, 0.0007269704, 0.0007023658, 
    0.000672325, 0.0006284718, 0.0006136103, 0.0006066328, 0.0006006565, 
    0.000643508,
  0.0009024143, 0.000957489, 0.0009836992, 0.0009719529, 0.001009877, 
    0.001179488, 0.001442146, 0.00166734, 0.001807133, 0.001930015, 
    0.002019183, 0.002004036, 0.001831342, 0.001665782, 0.001580285, 
    0.001522541, 0.001522302, 0.001584418, 0.001656945, 0.001710733, 
    0.001706457, 0.001619833, 0.001439667, 0.001257818, 0.001165756, 
    0.001110299, 0.001036866, 0.0009581088, 0.0008967714, 0.0008502328, 
    0.0008259933, 0.0008395994, 0.0008308413, 0.000774018, 0.0007316112, 
    0.0007311027, 0.0007534344, 0.0008309996, 0.0009043692, 0.0009248094, 
    0.001030318, 0.001163069, 0.001200485, 0.001219606, 0.001260439, 
    0.001295359, 0.001034006, 0.001081514, 0.001182476, 0.001291306, 
    0.001316802, 0.00128247, 0.001188422, 0.00105327, 0.0009783111, 
    0.0009238566, 0.0008383752, 0.0008014203, 0.0008072536, 0.00080417, 
    0.0007640994, 0.0007073721, 0.0007002992, 0.0006762031, 0.0006204606, 
    0.000598256, 0.0005911989, 0.0005865414, 0.0006029764, 0.0006342889, 
    0.0006426652, 0.0006384691, 0.000643889, 0.0006457805, 0.0006415844, 
    0.0006365776, 0.0006006081, 0.0005121073, 0.0005907221, 0.0007466632, 
    0.0007418157, 0.0007225038, 0.0007464569, 0.0008274079, 0.0008890787, 
    0.0008966126, 0.0009231088, 0.000949224, 0.0009236811, 0.0008856612, 
    0.0008450667, 0.0007862411, 0.0007713637, 0.000788196, 0.0008180458, 
    0.0008574808,
  0.0009430093, 0.0009566471, 0.0009601759, 0.0009619561, 0.001113336, 
    0.001405986, 0.001559878, 0.001651621, 0.001758575, 0.001805163, 
    0.001683537, 0.001549548, 0.001417177, 0.001298206, 0.001223517, 
    0.00121824, 0.001234977, 0.001235406, 0.001242622, 0.001229255, 
    0.001129039, 0.001014536, 0.0009314395, 0.0008589444, 0.0008224025, 
    0.000797749, 0.0007685344, 0.0007463293, 0.0007661972, 0.0009379862, 
    0.001061965, 0.0009845747, 0.0009411192, 0.0008732011, 0.0008193026, 
    0.0008868221, 0.0009358255, 0.0009428193, 0.0009442172, 0.0009065624, 
    0.001129882, 0.001264017, 0.00139068, 0.001405304, 0.001361436, 
    0.001372863, 0.001406702, 0.001163753, 0.001360528, 0.001370001, 
    0.001205, 0.001098395, 0.001056449, 0.0009853221, 0.0009482079, 
    0.0008796542, 0.0008107834, 0.000843748, 0.000874965, 0.0008536982, 
    0.0008648238, 0.0008688769, 0.0008544447, 0.0008250559, 0.0008249921, 
    0.0008047898, 0.0007607145, 0.0007500025, 0.000756837, 0.0007976377, 
    0.000869879, 0.0008614068, 0.0008283621, 0.0007916302, 0.0007003951, 
    0.0006165034, 0.000523726, 0.0004735794, 0.0006164401, 0.0006966754, 
    0.0007770853, 0.0008909702, 0.001129182, 0.001369748, 0.001607578, 
    0.001580636, 0.001459281, 0.001347478, 0.001230671, 0.001107265, 
    0.001015997, 0.0009664544, 0.0009573628, 0.0009322339, 0.0009154333, 
    0.0009386232,
  0.0009710314, 0.0009679324, 0.0009584432, 0.0009739087, 0.001152324, 
    0.001263205, 0.001414061, 0.001441862, 0.001570337, 0.001615033, 
    0.001245786, 0.00116857, 0.001189106, 0.00114643, 0.001128071, 
    0.001132171, 0.001132028, 0.001111445, 0.001015521, 0.0009155273, 
    0.0007935371, 0.0007392885, 0.0007542614, 0.0007574083, 0.0008595008, 
    0.0009488435, 0.0009576329, 0.001026234, 0.00113996, 0.001234866, 
    0.001067766, 0.001000469, 0.0009774528, 0.0009739716, 0.001003011, 
    0.001050632, 0.001013153, 0.001015154, 0.0009641489, 0.0008954848, 
    0.0009709042, 0.001531157, 0.001830038, 0.00177428, 0.001630005, 
    0.001582305, 0.001484347, 0.001331234, 0.001220052, 0.001040714, 
    0.0008889521, 0.0008362141, 0.0008506775, 0.0008631079, 0.0008722469, 
    0.0008871239, 0.0009151455, 0.0009973524, 0.001057943, 0.001082071, 
    0.00111812, 0.00110178, 0.001085345, 0.001051331, 0.001021401, 
    0.0009738291, 0.000936429, 0.0009078505, 0.000883786, 0.0008955952, 
    0.0009071985, 0.0008366108, 0.0007657688, 0.0007461868, 0.0006989008, 
    0.0006358959, 0.0005766242, 0.0005978425, 0.0007721428, 0.0008779843, 
    0.0009024939, 0.001154677, 0.001610407, 0.001947261, 0.001856535, 
    0.001714406, 0.001539471, 0.001333318, 0.001183034, 0.001107804, 
    0.001084026, 0.001056973, 0.001012961, 0.0009553758, 0.0009166878, 
    0.0009595556,
  0.0009798845, 0.0009921864, 0.001000309, 0.001030223, 0.001127641, 
    0.0009562969, 0.0007452327, 0.0009803935, 0.00151577, 0.001852816, 
    0.001724498, 0.001669663, 0.001683189, 0.00150927, 0.001452208, 0.001404, 
    0.001346511, 0.001416447, 0.001383004, 0.001323256, 0.001304707, 
    0.00129606, 0.001298889, 0.001293214, 0.001363007, 0.001397657, 
    0.001375008, 0.001440272, 0.001437188, 0.001218002, 0.001007272, 
    0.000713666, 0.0006144047, 0.000526635, 0.0006707194, 0.00100929, 
    0.001019224, 0.001068911, 0.001282294, 0.001252365, 0.001195717, 
    0.001650333, 0.001593797, 0.001614857, 0.001601617, 0.001567794, 
    0.001375135, 0.001159686, 0.001000342, 0.0008716276, 0.0008894131, 
    0.0009425329, 0.001034388, 0.001072042, 0.001061901, 0.001101702, 
    0.001115451, 0.001163086, 0.00119424, 0.001229923, 0.001222596, 
    0.001163738, 0.001155617, 0.001167282, 0.001101226, 0.001039475, 
    0.0009979578, 0.0008731857, 0.0008375496, 0.0008548275, 0.0007862905, 
    0.0007811571, 0.0007887064, 0.0007491121, 0.000705719, 0.0006347336, 
    0.0006483719, 0.0008533159, 0.001002407, 0.001167122, 0.001147668, 
    0.001460871, 0.001695601, 0.001967669, 0.001950806, 0.001644724, 
    0.001448155, 0.001359162, 0.001336544, 0.001288463, 0.001278593, 
    0.001207337, 0.001115148, 0.001072599, 0.001008734, 0.0009902157,
  0.0009707147, 0.0009618923, 0.001075936, 0.001264796, 0.001374531, 
    0.0009726686, 0.001033116, 0.001266527, 0.001789857, 0.002167609, 
    0.002088673, 0.001979607, 0.002003624, 0.001954606, 0.00194467, 
    0.001957084, 0.001983214, 0.001985821, 0.001925772, 0.001835903, 
    0.00175535, 0.001715582, 0.001709638, 0.001728998, 0.001711053, 
    0.001614795, 0.001500464, 0.001352185, 0.001241256, 0.001195654, 
    0.001029779, 0.0005864939, 0.0006624386, 0.0007168297, 0.0006946733, 
    0.001028666, 0.001230892, 0.001298936, 0.00149026, 0.00163784, 
    0.001464876, 0.001544811, 0.001356173, 0.001373976, 0.001389807, 
    0.00137442, 0.001344061, 0.001346637, 0.001361133, 0.001369382, 
    0.00136652, 0.001307218, 0.001294963, 0.001273696, 0.00123609, 
    0.001215729, 0.001178186, 0.001248392, 0.001288622, 0.001295918, 
    0.001299859, 0.001249982, 0.001214808, 0.001204968, 0.00115514, 
    0.001091847, 0.001060472, 0.0009564739, 0.0009161178, 0.0008911779, 
    0.0007513221, 0.0008151541, 0.000805188, 0.0007829526, 0.0007341392, 
    0.0007280996, 0.001103545, 0.0009137485, 0.00135619, 0.001472506, 
    0.001446614, 0.001738771, 0.001871936, 0.001976111, 0.002098308, 
    0.001847188, 0.001619674, 0.001561992, 0.001537483, 0.001468691, 
    0.001402076, 0.001320903, 0.001210087, 0.001143839, 0.001103531, 
    0.001043766,
  0.001173767, 0.001295138, 0.001465512, 0.001720033, 0.001146968, 
    0.001040698, 0.0015004, 0.001809201, 0.002043295, 0.002270637, 
    0.002478393, 0.002368084, 0.00231352, 0.002168338, 0.002150504, 
    0.002136787, 0.00223573, 0.002205738, 0.002093093, 0.001957291, 
    0.001845266, 0.001817706, 0.001736737, 0.001663002, 0.00158167, 
    0.001525419, 0.001488814, 0.001456611, 0.001429829, 0.001401314, 
    0.001269882, 0.0008830545, 0.001007304, 0.001329201, 0.001170462, 
    0.001286126, 0.001485189, 0.00178903, 0.001807849, 0.001751663, 
    0.001651876, 0.001655453, 0.001663447, 0.001787044, 0.001774599, 
    0.001709096, 0.001676594, 0.001636951, 0.001619278, 0.001534241, 
    0.001459807, 0.001397626, 0.001370954, 0.001334318, 0.001367903, 
    0.001409658, 0.001423407, 0.001507315, 0.001551883, 0.001632166, 
    0.001656899, 0.001626063, 0.001625157, 0.001538484, 0.001433023, 
    0.001265352, 0.001156681, 0.001083375, 0.000945854, 0.0008673826, 
    0.000800469, 0.0008818163, 0.0008433992, 0.0008401079, 0.0008182535, 
    0.00106942, 0.001814303, 0.001288813, 0.001378315, 0.001994166, 
    0.001650795, 0.001740617, 0.001909846, 0.001604526, 0.001998966, 
    0.001875036, 0.001745462, 0.001644836, 0.001586407, 0.001490213, 
    0.001363167, 0.001284457, 0.001205827, 0.001133618, 0.001119933, 
    0.001089081,
  0.001552471, 0.001643897, 0.00178617, 0.002062608, 0.001705678, 
    0.001669837, 0.002236541, 0.002422635, 0.002200843, 0.002186967, 
    0.002654123, 0.0026512, 0.001923849, 0.001991305, 0.002267377, 
    0.002332067, 0.002323627, 0.00221734, 0.002121559, 0.001999553, 
    0.001939726, 0.001911768, 0.001861813, 0.00180092, 0.001788888, 
    0.00179108, 0.001759911, 0.001749231, 0.001797232, 0.001843597, 
    0.001907921, 0.001822711, 0.001723623, 0.001447425, 0.001668327, 
    0.001664863, 0.001590189, 0.001865927, 0.002125581, 0.00206218, 
    0.002055581, 0.002181672, 0.002247189, 0.002253501, 0.002139076, 
    0.001948054, 0.001868264, 0.001801125, 0.001730856, 0.001627731, 
    0.001615286, 0.001631959, 0.00162789, 0.00165774, 0.00178701, 
    0.001913387, 0.002021105, 0.002106126, 0.002191719, 0.002274591, 
    0.00228006, 0.002209807, 0.002063465, 0.001888053, 0.001752518, 
    0.001562024, 0.001399644, 0.001315468, 0.001197276, 0.001111953, 
    0.001028936, 0.001015283, 0.0009950977, 0.001049821, 0.001146985, 
    0.001518632, 0.002188304, 0.001774057, 0.001761882, 0.002058491, 
    0.001660444, 0.002813753, 0.002512631, 0.001825828, 0.001823983, 
    0.002067139, 0.001807579, 0.001760276, 0.001693917, 0.001591381, 
    0.001573452, 0.001468215, 0.001396546, 0.001377027, 0.001403683, 
    0.001433056,
  0.001966543, 0.002002493, 0.00226051, 0.002477486, 0.002348758, 
    0.001801475, 0.002161217, 0.002068806, 0.00225954, 0.002167257, 
    0.00237341, 0.002735616, 0.002394344, 0.00205935, 0.002202176, 
    0.00235672, 0.002316172, 0.002298911, 0.002325932, 0.002314137, 
    0.002339396, 0.002267282, 0.0022494, 0.002213988, 0.002187157, 
    0.002183802, 0.00223217, 0.002242438, 0.002331701, 0.002474387, 
    0.002619934, 0.002615499, 0.002417707, 0.002627374, 0.002623592, 
    0.002162505, 0.002037605, 0.002613164, 0.00263683, 0.002538316, 
    0.002654538, 0.002858274, 0.002799145, 0.002665647, 0.002517589, 
    0.002309052, 0.002235493, 0.00214289, 0.002051003, 0.001988348, 
    0.00198509, 0.002009058, 0.002118286, 0.002314935, 0.00253536, 
    0.002673818, 0.002756787, 0.002762208, 0.002804345, 0.002782425, 
    0.002777911, 0.002736299, 0.002573013, 0.002426783, 0.002232614, 
    0.002047601, 0.001889562, 0.001767349, 0.001633342, 0.00153451, 
    0.001489704, 0.001487064, 0.001583766, 0.001633392, 0.001630624, 
    0.00194227, 0.002297609, 0.00228308, 0.001773676, 0.001770418, 
    0.001961851, 0.002431871, 0.002274673, 0.002120591, 0.001783308, 
    0.001814336, 0.001964871, 0.00195756, 0.001964029, 0.001886431, 
    0.001924451, 0.001845011, 0.001838446, 0.001832026, 0.001863275, 
    0.001921353,
  0.002414305, 0.002459477, 0.002634684, 0.002672466, 0.00235982, 
    0.001776186, 0.002080185, 0.001987108, 0.002187792, 0.002027878, 
    0.002212367, 0.0026999, 0.002525616, 0.002263625, 0.002375428, 
    0.002495306, 0.002602244, 0.002674976, 0.002738938, 0.002701251, 
    0.002729861, 0.002688328, 0.002697039, 0.002663342, 0.002657335, 
    0.002665473, 0.00271314, 0.002768502, 0.002924362, 0.003092371, 
    0.0032156, 0.003338672, 0.003294723, 0.003137365, 0.002981265, 
    0.003130833, 0.00317146, 0.003135649, 0.003002134, 0.002939543, 
    0.003167947, 0.003162209, 0.003083166, 0.002992457, 0.002861183, 
    0.002721898, 0.002682324, 0.00263208, 0.002595808, 0.002620349, 
    0.002630999, 0.002689777, 0.002821337, 0.002969775, 0.003157251, 
    0.003211185, 0.003262078, 0.00326645, 0.003233196, 0.003218079, 
    0.00317402, 0.003054731, 0.00291489, 0.002798223, 0.002636957, 
    0.002478392, 0.002352668, 0.002275817, 0.002209505, 0.002141858, 
    0.002159023, 0.002139044, 0.002073558, 0.001983023, 0.002045472, 
    0.002796873, 0.00263478, 0.001860158, 0.001023071, 0.0005913591, 
    0.001260124, 0.001002201, 0.001929666, 0.00242165, 0.001725595, 
    0.001673444, 0.002207438, 0.002285353, 0.002260686, 0.002312629, 
    0.002313629, 0.002283017, 0.002328841, 0.002318589, 0.002358373, 
    0.002408584,
  0.002890174, 0.002886915, 0.002963688, 0.003056178, 0.002699393, 
    0.002478059, 0.002335184, 0.002255298, 0.002131272, 0.002163983, 
    0.002335852, 0.002640279, 0.002520465, 0.002460448, 0.002596648, 
    0.002684036, 0.002885537, 0.002971655, 0.003107933, 0.003094312, 
    0.003124686, 0.003090419, 0.003072156, 0.003000991, 0.003034053, 
    0.00307557, 0.003086682, 0.003171798, 0.003308507, 0.003501261, 
    0.003614685, 0.003560133, 0.003518935, 0.003473653, 0.00342368, 
    0.003287112, 0.003257435, 0.003207954, 0.002836991, 0.003165612, 
    0.003343634, 0.003323875, 0.003240794, 0.003153406, 0.003041094, 
    0.002891939, 0.002777327, 0.002791297, 0.002798639, 0.002816902, 
    0.002889588, 0.002981586, 0.003127625, 0.003258217, 0.003402522, 
    0.003449744, 0.003436329, 0.003376136, 0.003264813, 0.00326273, 
    0.003219431, 0.003203377, 0.003183302, 0.003066191, 0.003003806, 
    0.002834607, 0.002727572, 0.002680206, 0.002651708, 0.002618837, 
    0.002550348, 0.002479188, 0.002399015, 0.002362029, 0.002621794, 
    0.003093372, 0.001380555, 0.0004950855, 0.0007144772, 0.0004964834, 
    0.0007234262, 0.001048184, 0.001093309, 0.002411366, 0.00233906, 
    0.002085258, 0.002288834, 0.002582263, 0.002574459, 0.002643887, 
    0.002664774, 0.00270958, 0.002717462, 0.002766688, 0.002810129, 
    0.002847258,
  0.0032722, 0.00327689, 0.003229061, 0.003192902, 0.003279909, 0.003383256, 
    0.003244226, 0.002763127, 0.002531736, 0.002215991, 0.002306811, 
    0.002471923, 0.002523201, 0.002601258, 0.002803342, 0.002896804, 
    0.003103195, 0.003198069, 0.003226124, 0.003173655, 0.003145728, 
    0.003099538, 0.003132235, 0.003203554, 0.003330471, 0.003330583, 
    0.003301065, 0.003319535, 0.003317039, 0.003445912, 0.003457008, 
    0.003388582, 0.003396705, 0.003403157, 0.003435059, 0.003349688, 
    0.003191171, 0.003002008, 0.002726667, 0.002907149, 0.00336412, 
    0.003223965, 0.003043322, 0.002948765, 0.002838219, 0.002708582, 
    0.002636611, 0.002677858, 0.002813645, 0.002938528, 0.003183164, 
    0.003390172, 0.003608661, 0.003679661, 0.003646329, 0.00363652, 
    0.003503118, 0.003382368, 0.003306344, 0.003249617, 0.003211677, 
    0.003208559, 0.003186036, 0.003111793, 0.003056876, 0.002933774, 
    0.002969394, 0.002898471, 0.002813928, 0.002794696, 0.002713902, 
    0.002643475, 0.002625307, 0.002666236, 0.00293719, 0.003281451, 
    0.001337608, 0.001565585, 0.002097753, 0.001131869, 0.0008300487, 
    0.0008328464, 0.001079863, 0.001443085, 0.00286077, 0.002524613, 
    0.002517971, 0.002713777, 0.002952892, 0.00298683, 0.003065731, 
    0.003159335, 0.003202312, 0.00323814, 0.00319338, 0.003220972,
  0.003509236, 0.00352785, 0.003408037, 0.002749617, 0.00360206, 0.003628763, 
    0.003941187, 0.003432481, 0.003116624, 0.002614594, 0.002482176, 
    0.002567499, 0.00258646, 0.002771648, 0.002947748, 0.003078543, 
    0.003224533, 0.003285397, 0.003187358, 0.003195131, 0.003221277, 
    0.00320589, 0.003248744, 0.003283694, 0.003467087, 0.00337442, 
    0.00337714, 0.003356921, 0.003297806, 0.003520619, 0.003382445, 
    0.00314304, 0.002980661, 0.003370067, 0.003548244, 0.003282867, 
    0.002937926, 0.002651151, 0.002789419, 0.003272073, 0.00336045, 
    0.003081182, 0.002942678, 0.002951609, 0.00293465, 0.002918201, 
    0.002979647, 0.003112128, 0.003404956, 0.003637841, 0.003816655, 
    0.003833186, 0.003716471, 0.003539247, 0.003342248, 0.003199056, 
    0.003126357, 0.003088877, 0.003082898, 0.003072405, 0.003106307, 
    0.003084296, 0.003077682, 0.003081784, 0.003099205, 0.003070911, 
    0.003016997, 0.002941912, 0.002963513, 0.002866523, 0.00286557, 
    0.002832366, 0.002814706, 0.002837723, 0.002833657, 0.003319485, 
    0.002156276, 0.002644078, 0.003114382, 0.002378022, 0.002058934, 
    0.00177625, 0.001423582, 0.002126901, 0.002573759, 0.002789132, 
    0.002785288, 0.002951102, 0.00321107, 0.003375059, 0.003484365, 
    0.00345224, 0.003469532, 0.003450634, 0.00340322, 0.00349099,
  0.003522955, 0.003574055, 0.003306551, 0.002802085, 0.003243733, 
    0.003796721, 0.003669614, 0.003370079, 0.00335412, 0.003251266, 
    0.00287234, 0.002559868, 0.002452502, 0.002804823, 0.003097249, 
    0.00325343, 0.003379269, 0.00336932, 0.003248997, 0.003160162, 
    0.003136607, 0.003114419, 0.003203301, 0.003188407, 0.003259219, 
    0.003207322, 0.003199853, 0.003188435, 0.0033742, 0.003472714, 
    0.003340835, 0.003055543, 0.002778834, 0.003105342, 0.003181143, 
    0.002941834, 0.002841907, 0.002835326, 0.003106073, 0.003420867, 
    0.003257468, 0.003027158, 0.002996163, 0.002965486, 0.003027173, 
    0.003138641, 0.003324369, 0.003536928, 0.003772566, 0.003929967, 
    0.004041802, 0.004067518, 0.00396066, 0.003786538, 0.003642801, 
    0.003413331, 0.003365804, 0.003271693, 0.00322862, 0.003232814, 
    0.003178375, 0.003147045, 0.003177248, 0.003143726, 0.003137589, 
    0.003099682, 0.003073867, 0.003109662, 0.003043666, 0.002910059, 
    0.002926003, 0.002796639, 0.00263612, 0.002581267, 0.00241353, 
    0.002741909, 0.002740574, 0.002848164, 0.003326768, 0.003060549, 
    0.002880431, 0.00166998, 0.001928441, 0.0031, 0.003010547, 0.002969442, 
    0.002927495, 0.003072852, 0.00322393, 0.003360908, 0.0034256, 
    0.003459791, 0.003531665, 0.003486222, 0.003463143, 0.003447106,
  0.003168572, 0.003470233, 0.00306573, 0.003013563, 0.003298618, 
    0.003372945, 0.003234532, 0.003101492, 0.003313497, 0.003412899, 
    0.003063424, 0.00299379, 0.002123786, 0.002830505, 0.003103003, 
    0.003272504, 0.003469948, 0.003506474, 0.00344272, 0.003268564, 
    0.003114577, 0.002955455, 0.002977883, 0.003092755, 0.003223279, 
    0.00322835, 0.002981838, 0.003002506, 0.003186882, 0.003258755, 
    0.003206909, 0.002979742, 0.002943553, 0.003050951, 0.00311216, 
    0.003032148, 0.003006876, 0.003058517, 0.003169477, 0.003115674, 
    0.003036391, 0.002950815, 0.002994906, 0.002942201, 0.002981795, 
    0.003013503, 0.002998324, 0.003020767, 0.003084617, 0.003114911, 
    0.003192587, 0.003259979, 0.003437061, 0.003503311, 0.003546989, 
    0.003514247, 0.003486682, 0.003408672, 0.003421515, 0.003400503, 
    0.003395941, 0.003432466, 0.003458645, 0.00342037, 0.003434677, 
    0.003321873, 0.00335053, 0.003358381, 0.003227029, 0.003320299, 
    0.003115576, 0.002918515, 0.002810579, 0.002840236, 0.002784556, 
    0.00274935, 0.002805154, 0.002811495, 0.002797669, 0.002328953, 
    0.002411764, 0.002653424, 0.002987973, 0.003020829, 0.003099842, 
    0.003177473, 0.003114909, 0.003146363, 0.003098283, 0.003058467, 
    0.003079323, 0.003126036, 0.003073268, 0.003071088, 0.002930149, 
    0.002930595,
  0.003128882, 0.003180381, 0.003226615, 0.003097884, 0.003171528, 
    0.00316833, 0.003170367, 0.003224537, 0.003455816, 0.003418749, 
    0.003024482, 0.003222688, 0.002585109, 0.002085893, 0.002976961, 
    0.003232418, 0.003400931, 0.003440622, 0.003436966, 0.003366427, 
    0.003182828, 0.003005713, 0.003032545, 0.002925575, 0.002932185, 
    0.003146764, 0.003260711, 0.003071262, 0.003208514, 0.003226744, 
    0.00320594, 0.003303578, 0.003200725, 0.002901383, 0.002988152, 
    0.003038093, 0.003052207, 0.003005017, 0.002986642, 0.002941946, 
    0.003015362, 0.003028588, 0.003085982, 0.003092293, 0.003080912, 
    0.003075143, 0.002980905, 0.002914624, 0.002939975, 0.002891846, 
    0.002926623, 0.002884155, 0.002937878, 0.002956744, 0.002995607, 
    0.003045183, 0.003006637, 0.00297728, 0.002990583, 0.002996672, 
    0.003099238, 0.003208483, 0.003361786, 0.003298955, 0.003376456, 
    0.003404429, 0.003450653, 0.003510447, 0.003530983, 0.003422534, 
    0.003154393, 0.003140246, 0.002741007, 0.002656782, 0.002733948, 
    0.002552085, 0.002575113, 0.002558598, 0.003022898, 0.002835818, 
    0.002945965, 0.002897454, 0.002980299, 0.002930276, 0.002925398, 
    0.003074426, 0.003038488, 0.003031272, 0.003016554, 0.00303906, 
    0.00307112, 0.003059471, 0.003072727, 0.002985207, 0.003099317, 
    0.003076907,
  0.00330857, 0.003290163, 0.003318757, 0.003567856, 0.003892248, 
    0.003655534, 0.002982568, 0.003238505, 0.003888164, 0.003671696, 
    0.003058705, 0.001878548, 0.002083016, 0.00187049, 0.003074983, 
    0.00300217, 0.003394304, 0.003457027, 0.003397595, 0.003363963, 
    0.002964625, 0.002964959, 0.003272919, 0.003200773, 0.003081247, 
    0.003217241, 0.003383862, 0.003056038, 0.002925921, 0.002955411, 
    0.00327063, 0.003428018, 0.003391366, 0.003152421, 0.003102321, 
    0.002975961, 0.003003141, 0.002956664, 0.002934586, 0.002905341, 
    0.002950085, 0.003027793, 0.003034087, 0.003026297, 0.003060378, 
    0.003048519, 0.003022881, 0.003023343, 0.003071073, 0.00300198, 
    0.003029177, 0.003046915, 0.003046246, 0.003056098, 0.003108313, 
    0.003143726, 0.003126752, 0.003109742, 0.003121648, 0.003144456, 
    0.003145793, 0.003137225, 0.003183575, 0.00307627, 0.003203364, 
    0.003289545, 0.003394067, 0.003598535, 0.003628401, 0.003415318, 
    0.003507331, 0.002949607, 0.002908075, 0.002086116, 0.002414785, 
    0.002540383, 0.002688171, 0.002719961, 0.002740497, 0.002808064, 
    0.002744947, 0.002661755, 0.002669718, 0.002672881, 0.002670642, 
    0.002640568, 0.002643066, 0.002699396, 0.002823977, 0.002939388, 
    0.002963005, 0.003008783, 0.003213234, 0.003124764, 0.00325672, 
    0.003264572,
  0.003863957, 0.003579871, 0.003383604, 0.003972418, 0.004122609, 
    0.003159001, 0.001865754, 0.001808852, 0.0028169, 0.003095388, 
    0.002951019, 0.002597872, 0.002257363, 0.003151179, 0.002676553, 
    0.003117088, 0.002955964, 0.003151404, 0.003222818, 0.003250254, 
    0.002877256, 0.003064383, 0.00342894, 0.003277941, 0.003153026, 
    0.003252909, 0.003050424, 0.003040843, 0.003046246, 0.003255229, 
    0.003177678, 0.003375201, 0.00339232, 0.003197944, 0.003083328, 
    0.003061553, 0.003037425, 0.003069198, 0.003040461, 0.00294406, 
    0.002885552, 0.002872186, 0.002876777, 0.002988055, 0.003018241, 
    0.002925033, 0.002929421, 0.002894549, 0.002900144, 0.002874617, 
    0.002827615, 0.002823547, 0.002847482, 0.002883118, 0.002958428, 
    0.002973782, 0.002964184, 0.002971144, 0.003030812, 0.003080007, 
    0.003083853, 0.00306613, 0.002914002, 0.00281137, 0.002843544, 
    0.002902512, 0.003299797, 0.003609931, 0.003826622, 0.003110396, 
    0.002877824, 0.002620745, 0.001313288, 0.002664743, 0.00281927, 
    0.002789833, 0.002723441, 0.002659133, 0.002717337, 0.00263297, 
    0.002569616, 0.002580822, 0.002533631, 0.002491409, 0.002501773, 
    0.002419472, 0.002446078, 0.002370756, 0.002416436, 0.002467347, 
    0.002582947, 0.002756327, 0.002379801, 0.002078915, 0.002977358, 
    0.003636425,
  0.002365558, 0.002026098, 0.001680946, 0.001941093, 0.001057118, 
    0.001645009, 0.001168856, 0.001172766, 0.001578364, 0.002046062, 
    0.003295012, 0.002343449, 0.002070189, 0.002532054, 0.003066684, 
    0.003167202, 0.003082581, 0.003015602, 0.003128437, 0.003351375, 
    0.003266066, 0.003362466, 0.003336543, 0.00321457, 0.003292708, 
    0.003143711, 0.003040779, 0.002857527, 0.002959127, 0.003284728, 
    0.003179459, 0.003283059, 0.003381098, 0.003185054, 0.00304197, 
    0.003104834, 0.003106901, 0.003180334, 0.003088128, 0.00292095, 
    0.002801105, 0.002779074, 0.002853302, 0.002891337, 0.002831701, 
    0.002772097, 0.002734935, 0.002694961, 0.002656016, 0.002631158, 
    0.002635259, 0.002706451, 0.002766054, 0.002794111, 0.002802294, 
    0.002733391, 0.002677077, 0.002596792, 0.002563097, 0.002547313, 
    0.002510708, 0.002490109, 0.002355799, 0.002197806, 0.001798123, 
    0.001735082, 0.002328876, 0.00290167, 0.003161848, 0.002786192, 
    0.002426672, 0.001777299, 0.002035934, 0.003013393, 0.002761813, 
    0.002769252, 0.002742117, 0.002637833, 0.002579611, 0.002545994, 
    0.002547937, 0.00250591, 0.002543513, 0.002453867, 0.002415977, 
    0.002350776, 0.00230829, 0.002251213, 0.002203114, 0.002109002, 
    0.00210123, 0.00243934, 0.001861143, 0.000711998, 0.0008291407, 
    0.001924897,
  0.001792242, 0.001749167, 0.001070134, 0.0008870452, 0.0009449488, 
    0.0011175, 0.0006212881, 0.000696724, 0.0008252, 0.001855279, 
    0.002973257, 0.00173289, 0.002059127, 0.002610589, 0.003362862, 
    0.004183039, 0.004043711, 0.003656996, 0.003629992, 0.003372673, 
    0.003486652, 0.003366044, 0.003253018, 0.003062489, 0.00309536, 
    0.003025202, 0.002784824, 0.002465233, 0.002411952, 0.002858942, 
    0.003045592, 0.003285952, 0.003214648, 0.00320133, 0.003168173, 
    0.003234264, 0.003153313, 0.003077623, 0.003008435, 0.002912907, 
    0.002866097, 0.002839951, 0.002847072, 0.002773797, 0.002716212, 
    0.002713636, 0.002646908, 0.002593869, 0.002595156, 0.00257168, 
    0.002534838, 0.002497612, 0.002543449, 0.002552146, 0.002492858, 
    0.002433285, 0.002391052, 0.002278836, 0.002238814, 0.002201254, 
    0.002141302, 0.002160771, 0.00220844, 0.001944399, 0.001493629, 
    0.001451254, 0.001494775, 0.002611974, 0.002702219, 0.002845018, 
    0.002863044, 0.002950624, 0.002823848, 0.002927134, 0.002901589, 
    0.002845641, 0.002701238, 0.002712887, 0.002690397, 0.002553783, 
    0.00257564, 0.002557565, 0.002577115, 0.002486262, 0.002419043, 
    0.002339315, 0.002255122, 0.002219455, 0.00215114, 0.002064339, 
    0.001904789, 0.002042293, 0.001443038, 0.001843423, 0.001938932, 
    0.001509333,
  0.001049328, 0.001706966, 0.001760134, 0.001289479, 0.001824268, 
    0.001777078, 0.0008382169, 0.0004561758, 0.001081848, 0.001322381, 
    0.001808851, 0.00143892, 0.001941332, 0.002064769, 0.003154518, 
    0.003616939, 0.003922973, 0.004015287, 0.004638387, 0.004427882, 
    0.00385323, 0.003366377, 0.003058657, 0.00270656, 0.002624718, 
    0.002721262, 0.002586508, 0.002039576, 0.002007136, 0.002529258, 
    0.002790533, 0.002974164, 0.003161449, 0.003084473, 0.003198341, 
    0.003255529, 0.003205001, 0.003174802, 0.003138879, 0.003092833, 
    0.00298246, 0.002901079, 0.002828935, 0.002755295, 0.002681989, 
    0.002566723, 0.002506053, 0.002457047, 0.002391227, 0.002376778, 
    0.002358437, 0.002362857, 0.002379339, 0.002330351, 0.002230755, 
    0.002173391, 0.002069967, 0.002006483, 0.00195907, 0.00189894, 
    0.001879836, 0.001856613, 0.001838446, 0.001636283, 0.00153408, 
    0.001637061, 0.001046085, 0.002678297, 0.003007046, 0.003245387, 
    0.003226411, 0.00324307, 0.00304113, 0.00300872, 0.002930691, 
    0.002575589, 0.002609206, 0.002639312, 0.002710011, 0.002607986, 
    0.002568644, 0.002520274, 0.002458256, 0.002445843, 0.002376016, 
    0.002280251, 0.002212794, 0.002172104, 0.002121369, 0.002028179, 
    0.001831627, 0.001799759, 0.002133575, 0.001529949, 0.001890692, 
    0.0007525929,
  0.001332315, 0.001009466, 3.536651e-005, 0.001555619, 0.00218498, 
    0.002585888, 0.002223669, 0.001578777, 0.002936618, 0.0025812, 
    0.00223446, 0.00180076, 0.002167003, 0.002815168, 0.002117396, 
    0.001958577, 0.002103472, 0.002090995, 0.003275873, 0.004320242, 
    0.004213748, 0.003094959, 0.002595664, 0.002246588, 0.002231346, 
    0.002200446, 0.002015925, 0.001587264, 0.001710876, 0.002191687, 
    0.002558235, 0.002865141, 0.003136892, 0.002679426, 0.002815565, 
    0.003038952, 0.003083659, 0.003043719, 0.003091926, 0.003130088, 
    0.002994699, 0.002827108, 0.002698643, 0.002616279, 0.002603056, 
    0.002554195, 0.002515061, 0.002420822, 0.002332593, 0.002268109, 
    0.002225081, 0.002241627, 0.002264388, 0.002280092, 0.002296321, 
    0.002238751, 0.002096685, 0.001991558, 0.001900911, 0.001841037, 
    0.001848079, 0.001751836, 0.001716043, 0.001721319, 0.001705265, 
    0.002297576, 0.002514044, 0.002575239, 0.003044209, 0.003213471, 
    0.003054749, 0.002908882, 0.002924921, 0.002949286, 0.002897151, 
    0.002806777, 0.002679795, 0.002460372, 0.00257243, 0.002577845, 
    0.00255521, 0.002472386, 0.002339095, 0.002310596, 0.00225625, 
    0.002251068, 0.002211793, 0.002162393, 0.002157354, 0.002083811, 
    0.001949342, 0.001767429, 0.00182128, 0.002252436, 0.002601115, 
    0.001657169,
  0.002899137, 0.002965863, 0.002522674, 0.002582868, 0.00269305, 
    0.002771409, 0.002657763, 0.002754434, 0.003250931, 0.002886072, 
    0.002915128, 0.002523582, 0.002457286, 0.002942692, 0.002803373, 
    0.002389145, 0.00283607, 0.002263547, 0.001813015, 0.001724196, 
    0.001955176, 0.001981115, 0.001930842, 0.001678372, 0.001712259, 
    0.001651907, 0.001423201, 0.001343315, 0.001636346, 0.002014304, 
    0.002088737, 0.00241429, 0.002733406, 0.002430296, 0.002526825, 
    0.002852568, 0.00272608, 0.002713172, 0.002765687, 0.002980238, 
    0.002960874, 0.002761668, 0.002583695, 0.002504175, 0.002478043, 
    0.002419854, 0.002379799, 0.002301089, 0.002248542, 0.002217627, 
    0.002159405, 0.002102263, 0.002078707, 0.002155001, 0.002219232, 
    0.002216832, 0.002160882, 0.002085812, 0.001953236, 0.001870697, 
    0.001849956, 0.001717363, 0.001774234, 0.001869999, 0.002572679, 
    0.002620124, 0.002752622, 0.002345386, 0.003117068, 0.00293719, 
    0.002904369, 0.003017269, 0.003207477, 0.003142865, 0.003179472, 
    0.003228379, 0.002904134, 0.00269245, 0.002655093, 0.002646035, 
    0.002607839, 0.002518894, 0.002414435, 0.002294, 0.002126853, 
    0.002045218, 0.0019979, 0.002015034, 0.002118237, 0.002097432, 
    0.002032408, 0.001852099, 0.001669789, 0.001969115, 0.002066644, 
    0.002786875,
  0.003296916, 0.002658002, 0.002814214, 0.00290262, 0.002805075, 
    0.002574969, 0.003098011, 0.002449197, 0.002666363, 0.002532897, 
    0.002529892, 0.002800434, 0.002742324, 0.002763525, 0.00237689, 
    0.002323978, 0.001587869, 0.001585119, 0.002575096, 0.002024143, 
    0.002095255, 0.001351516, 0.0006929727, 0.0008299525, 0.001408641, 
    0.001627779, 0.001898225, 0.001932287, 0.002080378, 0.002234747, 
    0.002157467, 0.002091313, 0.002222157, 0.002207548, 0.002261654, 
    0.002605836, 0.002541861, 0.002512678, 0.002537186, 0.00271144, 
    0.002782948, 0.002702489, 0.002572266, 0.002393755, 0.002301552, 
    0.002257143, 0.002185283, 0.002060272, 0.001962123, 0.001951426, 
    0.001956052, 0.00192636, 0.001884399, 0.001891932, 0.001932687, 
    0.001982293, 0.002027306, 0.00206841, 0.001999252, 0.001901517, 
    0.001827654, 0.001710447, 0.001781465, 0.002461038, 0.002749111, 
    0.002184504, 0.002047954, 0.002110991, 0.002611926, 0.003306245, 
    0.002829902, 0.002964083, 0.002948619, 0.002880717, 0.002966022, 
    0.003087918, 0.003149081, 0.003198846, 0.003002214, 0.002782964, 
    0.002668364, 0.00260687, 0.002519497, 0.002348344, 0.002056695, 
    0.00169592, 0.001429717, 0.001478146, 0.001711018, 0.00180877, 
    0.001844502, 0.0017598, 0.001668501, 0.001854086, 0.002677917, 0.003274996,
  0.002559679, 0.002310419, 0.002436688, 0.002810064, 0.001971706, 
    0.002456936, 0.001869426, 0.001974265, 0.001750072, 0.002115807, 
    0.001763933, 0.002076993, 0.002072367, 0.001942507, 0.001995787, 
    0.001716582, 0.001591063, 0.0008308745, 0.001512162, 0.002009456, 
    0.002275229, 0.002268236, 0.002306048, 0.002169244, 0.001563931, 
    0.001361053, 0.001511209, 0.001498604, 0.001787059, 0.002221269, 
    0.002270985, 0.002252643, 0.002164907, 0.00203535, 0.002069794, 
    0.002181212, 0.002040308, 0.002262372, 0.00258468, 0.002286008, 
    0.002095096, 0.001947848, 0.001826701, 0.001780844, 0.001750693, 
    0.001692438, 0.001604827, 0.001524561, 0.001469677, 0.001479039, 
    0.001502674, 0.001510003, 0.001515851, 0.001538754, 0.001594481, 
    0.001656311, 0.001727915, 0.001797725, 0.001821932, 0.00181079, 
    0.001765316, 0.001707618, 0.001814239, 0.001927757, 0.002482112, 
    0.002570073, 0.002041564, 0.002613229, 0.002796683, 0.002894863, 
    0.002911265, 0.002771044, 0.002579021, 0.002455249, 0.00281922, 
    0.002902777, 0.002935953, 0.002781583, 0.00258341, 0.002504651, 
    0.002240134, 0.001964189, 0.001812126, 0.001594274, 0.001393448, 
    0.001136304, 0.0008051563, 0.0007563606, 0.000955089, 0.001181078, 
    0.001399406, 0.001458187, 0.001410216, 0.001663226, 0.002427977, 
    0.002457144,
  0.001609978, 0.001711418, 0.001884954, 0.001999157, 0.00207178, 
    0.001886846, 0.001782339, 0.001796199, 0.001957051, 0.001812332, 
    0.001835824, 0.001724863, 0.001688864, 0.001722623, 0.002032108, 
    0.001988109, 0.002001397, 0.001828083, 0.00189662, 0.002093808, 
    0.002058347, 0.001985057, 0.002154891, 0.001796484, 0.001673905, 
    0.002203639, 0.002100626, 0.002174521, 0.002276834, 0.002263102, 
    0.002228293, 0.002167258, 0.00216996, 0.002183517, 0.002222237, 
    0.002250832, 0.002155306, 0.001931939, 0.001881345, 0.001578713, 
    0.001305676, 0.001376629, 0.001385102, 0.001377997, 0.001366363, 
    0.001302085, 0.001220975, 0.001198548, 0.001226536, 0.001261712, 
    0.001275381, 0.001279943, 0.001282232, 0.001287127, 0.001316151, 
    0.001383385, 0.00144156, 0.001499511, 0.00155875, 0.001619563, 
    0.00165574, 0.001707588, 0.00179337, 0.002027369, 0.002106873, 
    0.002206707, 0.002264135, 0.002592771, 0.002583632, 0.002616691, 
    0.002287165, 0.002215227, 0.002188365, 0.002189225, 0.002171644, 
    0.002306956, 0.00231913, 0.002317398, 0.00221448, 0.002198443, 
    0.001792193, 0.001427555, 0.0008977409, 0.0007949672, 0.0008473727, 
    0.0009082165, 0.0006799391, 0.00047288, 0.0004435237, 0.0004896177, 
    0.0008117212, 0.00111766, 0.001193254, 0.001274873, 0.001508586, 
    0.001820104,
  0.001335114, 0.001486477, 0.00170862, 0.001795087, 0.001689738, 
    0.001612506, 0.001383496, 0.001386152, 0.001307584, 0.001458917, 
    0.001528963, 0.001613682, 0.001776013, 0.001947802, 0.001916045, 
    0.001894508, 0.001994563, 0.002108098, 0.002234651, 0.002332306, 
    0.002477027, 0.002577115, 0.002353908, 0.002044757, 0.001944654, 
    0.001884524, 0.001903502, 0.00199078, 0.002048159, 0.002041214, 
    0.002027337, 0.001999124, 0.002062878, 0.00211441, 0.002185792, 
    0.002277996, 0.002283798, 0.002075068, 0.001267036, 0.001127083, 
    0.001301336, 0.001393811, 0.00136002, 0.001266242, 0.001260011, 
    0.001278735, 0.001264715, 0.001241843, 0.001219591, 0.00121123, 
    0.001223041, 0.001246533, 0.001300813, 0.001348655, 0.001356332, 
    0.001364104, 0.001357413, 0.001403857, 0.00145669, 0.001485412, 
    0.001526627, 0.001606211, 0.001682933, 0.00167815, 0.001719141, 
    0.001735799, 0.002023681, 0.002166448, 0.002034427, 0.001985249, 
    0.00181505, 0.001623648, 0.001749612, 0.001783276, 0.001844677, 
    0.001834759, 0.00178547, 0.001734002, 0.001622201, 0.001557145, 
    0.001500241, 0.001426125, 0.0008723894, 0.0008420148, 0.0008541737, 
    0.0007472686, 0.0004075384, 4.564971e-005, -0.00011444, -6.328989e-005, 
    0.0002797302, 0.0007302454, 0.0009974008, 0.001085378, 0.001190394, 
    0.001241622,
  0.001344523, 0.001224439, 0.001345684, 0.001305311, 0.001309984, 
    0.001311256, 0.00128123, 0.001180365, 0.001280373, 0.001432563, 
    0.001431704, 0.00138515, 0.001418241, 0.001599695, 0.001729775, 
    0.001712275, 0.001923864, 0.002150425, 0.00225285, 0.002179496, 
    0.002238767, 0.002431202, 0.002322483, 0.002098306, 0.002071794, 
    0.002165429, 0.002197155, 0.002201017, 0.00214127, 0.00203743, 
    0.001953618, 0.001960135, 0.001997646, 0.002009059, 0.002031295, 
    0.002121306, 0.002169625, 0.001964331, 0.001151084, 0.001028998, 
    0.001288636, 0.001509603, 0.001758337, 0.001346095, 0.001247104, 
    0.001238902, 0.00122482, 0.001203013, 0.001208211, 0.001234182, 
    0.001276446, 0.001349275, 0.001427619, 0.001501672, 0.001532269, 
    0.001508014, 0.00146521, 0.001445437, 0.001432736, 0.001445103, 
    0.001441256, 0.001674748, 0.001728932, 0.00172685, 0.001745495, 
    0.001769877, 0.001765315, 0.001687241, 0.001586311, 0.001523288, 
    0.00145108, 0.001522589, 0.001619689, 0.001609294, 0.001623551, 
    0.00119435, 0.001245339, 0.001172097, 0.001175419, 0.001222293, 
    0.001178805, 0.0007503512, 0.0006358461, 0.0005581062, 0.0005007265, 
    0.0004821462, 0.0003592013, 9.770459e-005, -0.0001151878, -8.929428e-005, 
    0.0001937868, 0.0005621761, 0.0008130409, 0.0009734165, 0.001157094, 
    0.001319171,
  0.000857655, 0.0009366842, 0.0009253984, 0.001164007, 0.001211612, 
    0.001416477, 0.001338451, 0.001185847, 0.001219781, 0.001278004, 
    0.001359686, 0.001503404, 0.001698955, 0.001540455, 0.001689053, 
    0.001737675, 0.001802048, 0.001878612, 0.00202891, 0.002128824, 
    0.002190574, 0.002335373, 0.002326362, 0.002343734, 0.002267727, 
    0.002191607, 0.002274292, 0.002357785, 0.002289279, 0.002134307, 
    0.001981752, 0.001890675, 0.001884874, 0.001956717, 0.002019454, 
    0.002088578, 0.002035777, 0.001883555, 0.001113208, 0.0009528636, 
    0.001010227, 0.001133474, 0.00165933, 0.001635409, 0.001133903, 
    0.00111076, 0.001178249, 0.00125494, 0.001355902, 0.001462395, 
    0.001561023, 0.001597452, 0.001591635, 0.00158914, 0.001647902, 
    0.001504056, 0.001463827, 0.001438459, 0.001428493, 0.001403985, 
    0.00153451, 0.001549833, 0.001566252, 0.001583259, 0.00167362, 
    0.001694108, 0.001611059, 0.001400106, 0.001398452, 0.001417336, 
    0.001391905, 0.001305786, 0.0009373836, 0.0008273134, 0.0007941101, 
    0.000807652, 0.0008249283, 0.0009069284, 0.0009797574, 0.0009510517, 
    0.0006337957, 0.0005161292, 0.0003699786, 0.0002258457, 0.0002525803, 
    0.0003730142, 0.0004377207, 0.0004120353, 0.0002870089, 0.0002713692, 
    0.0004197927, 0.0006171083, 0.0007425472, 0.0008166479, 0.000929324, 
    0.001069291,
  0.0006049485, 0.0006984412, 0.0008293162, 0.0009660251, 0.001111159, 
    0.001195685, 0.00130539, 0.001225853, 0.001226362, 0.001187914, 
    0.00119079, 0.001221562, 0.001287605, 0.001371337, 0.001452351, 
    0.001534877, 0.001592414, 0.001658265, 0.001719364, 0.00182705, 
    0.001891184, 0.001948707, 0.00203015, 0.002088325, 0.002114821, 
    0.00217282, 0.002180577, 0.002164381, 0.002143669, 0.002110498, 
    0.002031105, 0.00202694, 0.002070682, 0.002099086, 0.002089882, 
    0.002033091, 0.001948294, 0.001883793, 0.001888497, 0.00185159, 
    0.00180753, 0.001834282, 0.001802207, 0.001734098, 0.00168988, 
    0.001705218, 0.001558749, 0.001132092, 0.001171844, 0.001291387, 
    0.001392302, 0.00141085, 0.001627494, 0.001682807, 0.001699481, 
    0.001675655, 0.001593956, 0.001546876, 0.001494392, 0.001450666, 
    0.001426348, 0.001447932, 0.001467626, 0.001524926, 0.001660094, 
    0.001718426, 0.00162797, 0.00141182, 0.001259359, 0.00116102, 
    0.001023563, 0.0008489462, 0.0007544211, 0.0006537293, 0.0005964295, 
    0.000562971, 0.0006804941, 0.0008000536, 0.0006618672, 0.000597971, 
    0.0004832284, 0.0004091579, 0.0003195922, 0.0002259421, 0.0002049142, 
    0.0002261801, 0.0003709951, 0.000541083, 0.0006100652, 0.0006260071, 
    0.000628043, 0.0005713631, 0.000462994, 0.0004116707, 0.000524967, 
    0.0005883863,
  0.0003579776, 0.0004175673, 0.0005266834, 0.000850678, 0.0009576003, 
    0.001046134, 0.0008640452, 0.001078511, 0.001061695, 0.001038933, 
    0.001019923, 0.001017396, 0.001055526, 0.001138544, 0.001245276, 
    0.001333047, 0.001377249, 0.001412901, 0.001453782, 0.001525323, 
    0.001616145, 0.001713054, 0.001824173, 0.001913819, 0.001993402, 
    0.002075068, 0.002083747, 0.002071016, 0.00203441, 0.001968862, 
    0.001919905, 0.001898003, 0.001896557, 0.001920288, 0.001936738, 
    0.001862908, 0.001745351, 0.001740821, 0.001599583, 0.001620388, 
    0.001731523, 0.001732572, 0.001623933, 0.001565298, 0.001452256, 
    0.001406336, 0.00144407, 0.001406909, 0.00130353, 0.001326625, 
    0.001338577, 0.001177581, 0.001479324, 0.001543443, 0.001600695, 
    0.001627318, 0.0016078, 0.001597946, 0.001569287, 0.001527278, 
    0.001480278, 0.001473618, 0.001457231, 0.00145081, 0.00144469, 
    0.001378108, 0.001268403, 0.001172273, 0.001077763, 0.00101223, 
    0.001048787, 0.001012278, 0.001010355, 0.0009346646, 0.000487424, 
    0.0005165746, 0.0005563751, 0.000788562, 0.0008465615, 0.0008057281, 
    0.0005630348, 0.0005083573, 0.0006484515, 0.0005109799, 0.0004923197, 
    0.0005087708, 0.0004803354, 0.0004805881, 0.0005220412, 0.0006035166, 
    0.000587034, 0.0006890139, 0.0004584473, 0.0002696197, 0.0002188999, 
    0.0002489253,
  0.0004528998, 0.0004571122, 0.000453297, 0.0004308699, 0.0003853482, 
    0.0008303802, 0.000923268, 0.0009771194, 0.0009968127, 0.0009501302, 
    0.0008985838, 0.0007333285, 0.0007048929, 0.0007514004, 0.00103674, 
    0.001137384, 0.001254861, 0.001325989, 0.001397038, 0.001514802, 
    0.001632182, 0.001704725, 0.001774741, 0.001815399, 0.001803796, 
    0.001811632, 0.001838589, 0.001842483, 0.00180947, 0.001785088, 
    0.001715581, 0.001646552, 0.00154845, 0.001541282, 0.001496936, 
    0.001536084, 0.001560641, 0.00152394, 0.001470216, 0.001391474, 
    0.001220099, 0.001113479, 0.001007621, 0.0009646895, 0.0009806957, 
    0.000978407, 0.0009479052, 0.0009042588, 0.0008590231, 0.0005751783, 
    0.0006489605, 0.0007496681, 0.0008313819, 0.001215888, 0.001328548, 
    0.001422088, 0.00147036, 0.001501529, 0.001523925, 0.00141395, 
    0.001341788, 0.001313512, 0.001260822, 0.00120492, 0.001175372, 
    0.001154137, 0.001127101, 0.001100715, 0.001021322, 0.0006290758, 
    0.0009253984, 0.0008756649, 0.0008765389, 0.0006142789, 0.0008253101, 
    0.00050831, 0.0006648549, 0.0006756317, 0.0006128801, 0.0004712595, 
    0.0005033188, 0.0005132372, 0.0007333292, 0.0006959292, 0.0006895713, 
    0.0006407909, 0.0005948239, 0.0005708865, 0.0005644972, 0.0005527511, 
    0.0005306734, 0.0005129506, 0.0004208088, 0.0004182979, 0.0004251003, 
    0.0004634694,
  0.0006662216, 0.0006691138, 0.000629107, 0.0005634786, 0.0005011084, 
    0.0005561989, 0.0007286235, 0.0008559073, 0.0008686702, 0.0008083829, 
    0.0007101381, 0.0006410764, 0.0005977163, 0.0005810591, 0.0005630981, 
    0.0007052911, 0.000504304, 0.0005380961, 0.000578675, 0.001034595, 
    0.001248853, 0.001397944, 0.001516247, 0.001635154, 0.001705186, 
    0.001735704, 0.001714469, 0.001685048, 0.001662096, 0.001548846, 
    0.001483615, 0.001356633, 0.001226457, 0.001130566, 0.001011818, 
    0.0005713161, 0.0005531325, 0.0005361889, 0.0008008801, 0.0007135239, 
    0.000416948, 0.0003551973, 0.0002850548, 0.0002324118, 0.0002052959, 
    0.0002001617, 0.0002106682, 0.0002249097, 0.0002228753, 0.0002161516, 
    0.0002069327, 0.0002125276, 0.0002315058, 0.0002806678, 0.0003342484, 
    0.0003749703, 0.0003879245, 0.0003825361, 0.0003898158, 0.000398685, 
    0.0004223997, 0.0004621998, 0.0005222494, 0.000779788, 0.0008393298, 
    0.0008942932, 0.0009311368, 0.0009074542, 0.0008556535, 0.0005601896, 
    0.0007125707, 0.0006672712, 0.0005357435, 0.0006044717, 0.0006173782, 
    0.0005787865, 0.0005483641, 0.0004417752, 0.0004233215, 0.0004492614, 
    0.0004653945, 0.0007194853, 0.0005984794, 0.000606252, 0.0006015791, 
    0.0006040743, 0.0006109567, 0.0006343219, 0.0006628048, 0.0006633769, 
    0.0007397346, 0.0005195632, 0.0004758055, 0.0004479582, 0.0004867082, 
    0.0005911994,
  0.0004883618, 0.0005237907, 0.0006237989, 0.0007042256, 0.0007137624, 
    0.0007114899, 0.0007227752, 0.0006951501, 0.0006293631, 0.0005627808, 
    0.0005008234, 0.0004596885, 0.0004334943, 0.0003884167, 0.0003250293, 
    0.0002739285, 0.0002488946, 0.0002342875, 0.0002440468, 0.0002795709, 
    0.0003497456, 0.0004159308, 0.0004953556, 0.0005387163, 0.0005865113, 
    0.0008620434, 0.0008654608, 0.0009028763, 0.0008706106, 0.000807239, 
    0.0007601115, 0.0004939414, 0.0004382783, 0.0003760355, 0.0002994235, 
    0.0002374665, 0.0002021962, 0.0002002253, 0.0002158016, 0.0002263875, 
    0.0002351773, 0.0002400093, 0.0002343827, 0.0002257999, 0.0002240674, 
    0.0002265945, 0.0002340332, 0.0002431564, 0.0002569691, 0.0002696686, 
    0.0002805248, 0.000294623, 0.0003065758, 0.0003173524, 0.0003211829, 
    0.0003232176, 0.000323297, 0.0003255382, 0.000325093, 0.0003287965, 
    0.0003315464, 0.0003434671, 0.000368485, 0.0004224794, 0.0004685735, 
    0.0005777532, 0.0006184112, 0.0006398852, 0.0006749167, 0.0006641878, 
    0.0006348938, 0.000580821, 0.0005560566, 0.0005514477, 0.000514159, 
    0.0004577013, 0.0004811937, 0.0004915094, 0.0005950783, 0.0006311268, 
    0.0006471805, 0.000626152, 0.0005734138, 0.000513825, 0.0004742158, 
    0.0004764731, 0.000519245, 0.0005776258, 0.0006350211, 0.0006694169, 
    0.000655557, 0.0006444312, 0.0004595609, 0.0003811533, 0.0004009737, 
    0.0004517729,
  0.0003777039, 0.0003610624, 0.0004026904, 0.0004161848, 0.0004822584, 
    0.0004838957, 0.0004737708, 0.0003934081, 0.000354514, 0.000321819, 
    0.0002938602, 0.0002752796, 0.0002508815, 0.0002439513, 0.0002521211, 
    0.0002592099, 0.0002759469, 0.0002995823, 0.0003110738, 0.0003184332, 
    0.0003230744, 0.0003178292, 0.0003089122, 0.0003060829, 0.000301108, 
    0.0004376585, 0.0004248791, 0.0003142846, 0.0003331357, 0.0003428471, 
    0.0003482832, 0.0003487759, 0.0003395092, 0.0003293208, 0.000315286, 
    0.0003031425, 0.0003017122, 0.0003066077, 0.0003152546, 0.0003265871, 
    0.0003380789, 0.0003513033, 0.0003615872, 0.0003668324, 0.000368692, 
    0.0003666098, 0.0003616507, 0.0003573908, 0.0003551338, 0.0003566756, 
    0.0003589327, 0.0003674682, 0.0003797067, 0.0003924225, 0.0004068071, 
    0.0004210169, 0.000432747, 0.0004449859, 0.0004558577, 0.0004706397, 
    0.0004814956, 0.000490508, 0.0005014117, 0.0005125697, 0.0005228852, 
    0.0005321677, 0.0005393361, 0.000546902, 0.0005519884, 0.000554865, 
    0.0005294497, 0.0006523463, 0.0007611767, 0.0005146838, 0.0005046858, 
    0.0005048447, 0.0005043518, 0.0005062273, 0.0005096447, 0.0005163682, 
    0.0005057985, 0.0004863911, 0.0004702102, 0.0004587503, 0.0004592112, 
    0.0004677465, 0.0004898401, 0.0005210732, 0.0005600466, 0.0005869082, 
    0.000601436, 0.0005927419, 0.000531977, 0.0004894431, 0.0004490071, 
    0.0003949814,
  0.0006130552, 0.0005854461, 0.0005615568, 0.0005409415, 0.0005263344, 
    0.0005091683, 0.000493051, 0.0004804148, 0.0004746134, 0.0004688594, 
    0.0004681919, 0.0004669202, 0.0004643295, 0.0004601015, 0.0004567318, 
    0.000453823, 0.0004480379, 0.0004431899, 0.0004358625, 0.000425356, 
    0.0004140076, 0.0003992412, 0.0003876223, 0.0003782604, 0.0003718387, 
    0.0003691053, 0.0003693595, 0.0003744618, 0.0003815347, 0.0003889098, 
    0.000398383, 0.0004093184, 0.0004160576, 0.0004206831, 0.0004221771, 
    0.0004233057, 0.0004221932, 0.0004214144, 0.0004167415, 0.0004114325, 
    0.0004060282, 0.00040037, 0.0003983988, 0.0003987008, 0.0004013395, 
    0.0004036282, 0.0004079517, 0.0004142299, 0.0004195068, 0.0004278836, 
    0.0004360371, 0.0004408692, 0.0004503899, 0.0004612142, 0.0004723244, 
    0.0004839753, 0.0004944815, 0.0005041615, 0.0005124107, 0.0005218519, 
    0.0005318655, 0.0005392563, 0.0005499695, 0.0005601894, 0.0005676125, 
    0.0005743993, 0.0005790563, 0.000579867, 0.0005831735, 0.0005948716, 
    0.0006145812, 0.0006382321, 0.0006574485, 0.0006738997, 0.000702176, 
    0.0007230456, 0.0007466963, 0.0007738285, 0.0008057924, 0.0008302224, 
    0.0008557332, 0.0008726451, 0.0008922112, 0.0009024793, 0.0009074542, 
    0.0009061827, 0.0009044183, 0.0008898589, 0.0008687826, 0.0008411261, 
    0.0008020254, 0.0007486355, 0.0007136199, 0.0006898895, 0.0006663974, 
    0.0006419357,
  0.0006766813, 0.0006680661, 0.0006647443, 0.0006638383, 0.0006566381, 
    0.0006503121, 0.0006404892, 0.0006301261, 0.0006203665, 0.0006096379, 
    0.0005998625, 0.0005901351, 0.0005813295, 0.0005737636, 0.0005637184, 
    0.0005543248, 0.0005461073, 0.0005378101, 0.0005300536, 0.0005229011, 
    0.0005159234, 0.0005098518, 0.0005041137, 0.0005006487, 0.0004953716, 
    0.0004912233, 0.0004887597, 0.0004874244, 0.0004863117, 0.0004870908, 
    0.0004867411, 0.0004878535, 0.0004890617, 0.0004918112, 0.0004932578, 
    0.0004932575, 0.0004934643, 0.0004950063, 0.0004947518, 0.0004957849, 
    0.0004960075, 0.0004965321, 0.0004986462, 0.0004994567, 0.0005021745, 
    0.0005045587, 0.0005086595, 0.0005121564, 0.0005160824, 0.0005188955, 
    0.0005226305, 0.0005256189, 0.0005312455, 0.000536904, 0.0005411, 
    0.0005478712, 0.0005555165, 0.0005603165, 0.0005640679, 0.0005696625, 
    0.000575528, 0.000582871, 0.0005920581, 0.0006000213, 0.0006114019, 
    0.0006214629, 0.0006298553, 0.0006377709, 0.0006470534, 0.000657496, 
    0.0006692105, 0.000678763, 0.0006876322, 0.0006974551, 0.0007071353, 
    0.0007180071, 0.0007287199, 0.0007398142, 0.0007488742, 0.0007557247, 
    0.0007641013, 0.0007679637, 0.0007670736, 0.0007690126, 0.0007700613, 
    0.0007679157, 0.0007625592, 0.0007576479, 0.00074827, 0.0007357928, 
    0.0007281473, 0.0007190877, 0.0007107588, 0.0007028908, 0.0006951978, 
    0.0006882206,
  4.820882e-006, 4.518879e-006, 4.232779e-006, 3.946676e-006, 3.803621e-006, 
    3.596993e-006, 3.469837e-006, 3.342679e-006, 3.279101e-006, 
    3.263205e-006, 3.183733e-006, 3.104263e-006, 3.167842e-006, 
    3.088366e-006, 3.136051e-006, 3.19963e-006, 3.231419e-006, 3.231419e-006, 
    3.358575e-006, 3.374471e-006, 3.565206e-006, 3.708256e-006, 
    3.867202e-006, 3.930782e-006, 4.1692e-006, 4.359934e-006, 4.502985e-006, 
    4.677825e-006, 4.836769e-006, 5.043401e-006, 5.28182e-006, 5.552025e-006, 
    5.790442e-006, 6.044758e-006, 6.410331e-006, 6.728224e-006, 7.06201e-006, 
    7.379902e-006, 7.666005e-006, 7.999792e-006, 8.413053e-006, 
    8.746843e-006, 9.064737e-006, 9.382627e-006, 9.73231e-006, 9.907151e-006, 
    1.025683e-005, 1.047935e-005, 1.070188e-005, 1.079724e-005, 
    1.086083e-005, 1.090851e-005, 1.084493e-005, 1.094029e-005, 
    1.071777e-005, 1.079724e-005, 1.071777e-005, 1.057472e-005, 
    1.024094e-005, 1.003431e-005, 1.014557e-005, 1.006609e-005, 
    9.970729e-006, 9.811782e-006, 9.764099e-006, 9.652838e-006, 
    9.684623e-006, 9.573363e-006, 9.652835e-006, 9.716412e-006, 
    9.811782e-006, 9.986623e-006, 1.00502e-005, 9.764099e-006, 1.00661e-005, 
    1.03363e-005, 1.011378e-005, 1.024094e-005, 1.036809e-005, 1.030451e-005, 
    1.012967e-005, 9.907148e-006, 9.684623e-006, 9.382627e-006, 
    9.112424e-006, 8.746847e-006, 8.444847e-006, 8.06338e-006, 7.618331e-006, 
    7.173283e-006, 6.855393e-006, 6.410344e-006, 6.060662e-006, 
    5.742768e-006, 5.424878e-006, 5.059304e-006,
  5.742768e-006, 5.329508e-006, 4.963929e-006, 4.550669e-006, 4.04204e-006, 
    3.485729e-006, 3.088364e-006, 2.722791e-006, 2.500266e-006, 
    2.468476e-006, 2.389007e-006, 2.389006e-006, 2.452585e-006, 
    2.627426e-006, 2.770476e-006, 2.961212e-006, 3.072473e-006, 
    3.247314e-006, 3.294998e-006, 3.342682e-006, 3.358576e-006, 
    3.549311e-006, 3.75594e-006, 3.867202e-006, 4.073832e-006, 4.280461e-006, 
    4.471196e-006, 4.614247e-006, 4.916245e-006, 5.202347e-006, 5.42487e-006, 
    5.742762e-006, 6.283175e-006, 6.82359e-006, 7.713685e-006, 8.826308e-006, 
    1.006609e-005, 1.170324e-005, 1.334038e-005, 1.512056e-005, 
    1.696433e-005, 1.879219e-005, 2.031808e-005, 2.192343e-005, 
    2.303605e-005, 2.309963e-005, 2.438709e-005, 2.475266e-005, 
    2.478444e-005, 2.470498e-005, 2.480035e-005, 2.616728e-005, 
    2.599244e-005, 2.685075e-005, 2.535667e-005, 2.785211e-005, 
    2.756601e-005, 2.689843e-005, 2.638981e-005, 2.583351e-005, 
    2.538846e-005, 2.462551e-005, 2.383077e-005, 2.294068e-005, 
    2.203468e-005, 2.104924e-005, 1.976177e-005, 1.829946e-005, 
    1.686895e-005, 1.547023e-005, 1.485035e-005, 1.461193e-005, 
    1.481856e-005, 1.539076e-005, 1.599475e-005, 1.694842e-005, 
    1.766368e-005, 1.839484e-005, 1.834716e-005, 1.842662e-005, 
    1.858558e-005, 1.745707e-005, 1.710738e-005, 1.458015e-005, 
    1.343574e-005, 1.125819e-005, 9.81176e-006, 8.428942e-006, 7.443472e-006, 
    6.871276e-006, 6.601062e-006, 6.616952e-006, 6.696435e-006, 
    6.712336e-006, 6.648763e-006, 6.235503e-006,
  4.757308e-006, 3.438054e-006, 2.484376e-006, 1.975748e-006, 1.657854e-006, 
    1.419437e-006, 1.451228e-006, 1.546593e-006, 1.84859e-006, 2.198272e-006, 
    2.627425e-006, 3.215523e-006, 3.883098e-006, 4.63014e-006, 5.440762e-006, 
    6.060651e-006, 6.601065e-006, 6.855378e-006, 6.775905e-006, 
    6.108332e-006, 5.234133e-006, 4.137408e-006, 3.263209e-006, 2.75458e-006, 
    2.563847e-006, 2.595637e-006, 3.02479e-006, 3.37447e-006, 3.835413e-006, 
    4.280461e-006, 4.72551e-006, 5.138768e-006, 5.695078e-006, 6.108337e-006, 
    6.934853e-006, 8.095154e-006, 9.875355e-006, 1.218007e-005, 
    1.512057e-005, 1.845842e-005, 2.173269e-005, 2.425993e-005, 
    2.659643e-005, 2.769315e-005, 2.791567e-005, 2.802694e-005, 
    2.716863e-005, 2.605602e-005, 2.55156e-005, 2.66759e-005, 2.894883e-005, 
    3.231847e-005, 3.614909e-005, 4.009093e-005, 4.274534e-005, 4.39374e-005, 
    4.288836e-005, 4.029753e-005, 3.661001e-005, 3.269994e-005, 
    3.017271e-005, 2.910776e-005, 2.898062e-005, 2.918726e-005, 2.93303e-005, 
    2.925083e-005, 2.896473e-005, 2.829717e-005, 2.64216e-005, 2.282942e-005, 
    1.944388e-005, 1.634444e-005, 1.419867e-005, 1.345162e-005, 
    1.403972e-005, 1.602654e-005, 1.81882e-005, 2.184397e-005, 2.632623e-005, 
    2.9982e-005, 3.250921e-005, 3.362184e-005, 3.276354e-005, 3.036344e-005, 
    2.63898e-005, 2.251154e-005, 1.945977e-005, 1.861733e-005, 1.81246e-005, 
    1.718686e-005, 1.750475e-005, 1.610605e-005, 1.394436e-005, 
    1.109923e-005, 8.460716e-006, 6.362654e-006,
  7.093811e-006, 5.965296e-006, 5.170556e-006, 4.582456e-006, 4.07383e-006, 
    3.787727e-006, 3.771835e-006, 3.883095e-006, 3.994357e-006, 
    4.344036e-006, 4.518877e-006, 4.630139e-006, 4.693718e-006, 
    5.122871e-006, 5.997072e-006, 7.634215e-006, 9.477992e-006, 
    1.125819e-005, 1.262512e-005, 1.275227e-005, 1.12264e-005, 8.874002e-006, 
    6.585182e-006, 4.820877e-006, 3.978461e-006, 3.962567e-006, 
    4.216882e-006, 4.836771e-006, 5.408973e-006, 5.822232e-006, 
    5.854021e-006, 5.663287e-006, 5.313605e-006, 5.329497e-006, 
    5.552023e-006, 6.108334e-006, 7.364006e-006, 8.746836e-006, 
    1.020915e-005, 1.18145e-005, 1.361058e-005, 1.624907e-005, 1.955513e-005, 
    2.222542e-005, 2.483213e-005, 2.767729e-005, 3.975714e-005, 
    3.111051e-005, 3.298605e-005, 2.993429e-005, 3.425758e-005, 
    4.203005e-005, 5.193235e-005, 6.283601e-005, 7.372376e-005, 
    8.063792e-005, 7.98273e-005, 6.482282e-005, 5.269531e-005, 4.039289e-005, 
    3.187339e-005, 2.813812e-005, 2.731162e-005, 2.834483e-005, 
    3.049057e-005, 3.201645e-005, 3.255687e-005, 3.23979e-005, 3.146012e-005, 
    2.988658e-005, 2.855144e-005, 2.740702e-005, 2.767723e-005, 
    2.953691e-005, 3.236617e-005, 3.527486e-005, 3.891473e-005, 
    4.374667e-005, 4.911901e-005, 5.401457e-005, 6.480695e-005, 
    6.868521e-005, 7.062434e-005, 7.008392e-005, 6.793815e-005, 
    6.539503e-005, 6.680965e-005, 6.89872e-005, 7.429597e-005, 5.706631e-005, 
    5.027934e-005, 4.098099e-005, 3.09039e-005, 2.178039e-005, 1.446888e-005, 
    9.589254e-006,
  2.931442e-005, 2.492751e-005, 2.106514e-005, 1.766368e-005, 1.450066e-005, 
    1.283173e-005, 1.327678e-005, 1.532718e-005, 1.772726e-005, 
    1.895114e-005, 1.804515e-005, 1.524772e-005, 1.187808e-005, 
    9.573359e-006, 8.76273e-006, 9.525675e-006, 1.181449e-005, 1.450068e-005, 
    1.648749e-005, 1.712327e-005, 2.001609e-005, 1.96664e-005, 1.728221e-005, 
    1.413509e-005, 1.143303e-005, 1.027272e-005, 9.923046e-006, 
    1.038399e-005, 1.144892e-005, 1.275228e-005, 1.313375e-005, 
    1.264102e-005, 1.194165e-005, 1.146481e-005, 1.175092e-005, 
    1.245028e-005, 1.272047e-005, 1.2339e-005, 1.111513e-005, 1.094028e-005, 
    1.311783e-005, 1.554971e-005, 1.887169e-005, 2.139891e-005, 
    2.308375e-005, 2.418047e-005, 2.629447e-005, 2.658051e-005, 
    2.570632e-005, 2.735932e-005, 3.629207e-005, 5.399861e-005, 
    7.222968e-005, 8.982499e-005, 0.0001018571, 0.00010564, 0.0001033036, 
    9.384626e-005, 8.704345e-005, 8.189358e-005, 7.995439e-005, 
    8.032002e-005, 7.99704e-005, 8.095583e-005, 7.912796e-005, 7.545628e-005, 
    7.178466e-005, 7.138721e-005, 7.613981e-005, 8.014514e-005, 
    7.294494e-005, 8.960237e-005, 9.770866e-005, 0.0001094865, 0.0001242527, 
    0.0001404969, 0.0001211532, 0.000121328, 0.0001220115, 0.0001216459, 
    0.0001373499, 0.0001354902, 0.000131898, 0.0001223295, 0.0001122523, 
    0.0001018572, 9.801073e-005, 9.653246e-005, 9.422775e-005, 8.985674e-005, 
    8.960243e-005, 5.825837e-005, 5.142375e-005, 4.487518e-005, 3.86445e-005, 
    3.354235e-005,
  0.0001057354, 0.0001037804, 5.619209e-005, 4.233206e-005, 3.320856e-005, 
    3.134891e-005, 3.713454e-005, 4.913496e-005, 6.388512e-005, 
    7.456624e-005, 7.50272e-005, 6.591959e-005, 5.115356e-005, 3.605374e-005, 
    2.683486e-005, 2.281353e-005, 2.271817e-005, 2.535666e-005, 
    3.052241e-005, 3.360596e-005, 3.67372e-005, 3.743656e-005, 3.60378e-005, 
    3.219131e-005, 2.979126e-005, 2.848791e-005, 2.929852e-005, 
    3.204826e-005, 3.637155e-005, 3.913722e-005, 3.842196e-005, 
    3.382843e-005, 3.020446e-005, 2.872631e-005, 2.979125e-005, 
    3.227076e-005, 3.289065e-005, 3.125351e-005, 2.871035e-005, 
    2.928256e-005, 3.335155e-005, 3.611723e-005, 3.707089e-005, 
    3.535429e-005, 3.521121e-005, 3.2382e-005, 3.26522e-005, 4.43029e-005, 
    6.200955e-005, 8.456397e-005, 0.0001133649, 0.0001380492, 0.000154214, 
    0.0001617005, 0.000157377, 0.000144407, 0.000134457, 0.0001343298, 
    0.0001450588, 0.0001526723, 0.0001560102, 0.0001569003, 0.0001589984, 
    0.0001603176, 0.0001580924, 0.0001490007, 0.0001436761, 0.0001464098, 
    0.0001624156, 0.0001921701, 0.0002182849, 0.0002331463, 0.0002444157, 
    0.0002506622, 0.0002512027, 0.0002512027, 0.0002425879, 0.0002279172, 
    0.0002057124, 0.000198242, 0.0002297928, 0.000217395, 0.0002021521, 
    0.0001806785, 0.0001610168, 0.0001535782, 0.0001604923, 0.0001660555, 
    0.000159793, 0.000143501, 0.0001352359, 0.0001347272, 0.0001379697, 
    0.0001392095, 0.0001319455, 0.0001186418,
  0.0001935689, 0.000196875, 0.0001909146, 0.0001711257, 0.0001506218, 
    0.0001350451, 0.0001295932, 0.0001286237, 0.0001306105, 0.000141085, 
    0.0001569477, 0.0001707283, 0.0001770862, 0.0001681376, 0.0001497952, 
    0.0001369206, 0.0001303243, 0.0001294024, 0.0001360145, 0.0001451858, 
    0.0001476494, 0.0001388598, 0.0001274634, 0.0001145252, 0.0001052586, 
    0.0001048931, 0.0001073568, 0.0001072455, 9.802659e-005, 8.098764e-005, 
    5.612848e-005, 3.824721e-005, 3.196893e-005, 5.767029e-005, 
    7.656892e-005, 9.948888e-005, 0.000132502, 0.0001611601, 0.0001907715, 
    0.0002094635, 0.0002147405, 0.0002125788, 0.0002069364, 0.0002043298, 
    0.0002007217, 0.0002075882, 0.000220558, 0.0002181581, 0.0001906605, 
    0.000142945, 0.0001132856, 9.265461e-005, 9.422807e-005, 0.000115797, 
    0.0001426906, 0.0001555175, 0.000158744, 0.0001619229, 0.0001728107, 
    0.000183031, 0.0001940143, 0.0002054584, 0.0002271862, 0.0002556852, 
    0.0002758234, 0.0003016044, 0.0003200899, 0.0003467769, 0.0003920606, 
    0.0004254392, 0.0004749509, 0.0005450142, 0.0005516423, 0.0005826209, 
    0.0005399438, 0.0005167378, 0.0004689903, 0.0004090042, 0.0003553282, 
    0.0003169904, 0.0003067385, 0.0003194225, 0.0003278784, 0.0003146381, 
    0.0002927035, 0.0002830238, 0.0002848833, 0.0002826104, 0.0002704193, 
    0.0002556055, 0.0002487867, 0.0002467365, 0.0002342909, 0.0002138027, 
    0.0001943636, 0.0001892138,
  0.0003133188, 0.0003120949, 0.0003179917, 0.0003321698, 0.0003512432, 
    0.0003485888, 0.0003468721, 0.0003312796, 0.0003185003, 0.0003200899, 
    0.0003437252, 0.0003546289, 0.0003870695, 0.0004052847, 0.0004399349, 
    0.0004463086, 0.0004163632, 0.0004299055, 0.0004393945, 0.0004285226, 
    0.0004244377, 0.000388198, 0.0003485728, 0.0003105371, 0.0002721358, 
    0.00023321, 0.0002162507, 0.000204441, 0.0001938713, 0.000158347, 
    6.708014e-005, 9.704125e-005, 0.0001287672, 0.0001417056, 0.0001674541, 
    0.0003003962, 0.0003726215, 0.0003884365, 0.0004318762, 0.0003926007, 
    0.0003713018, 0.0003463947, 0.0003232684, 0.0003473645, 0.0003950165, 
    0.0004098143, 0.0003538812, 0.0001935209, -1.331326e-006, -0.0001568273, 
    -0.0002200399, -0.0002036847, -0.0001741524, -0.0001381829, 
    -7.972261e-005, -2.156408e-005, 2.797926e-005, 4.899176e-005, 
    8.602627e-005, 0.00015992, 0.0002390752, 0.0003360636, 0.0003850029, 
    0.0004079072, 0.0004671619, 0.000558333, 0.0006160464, 0.0006507917, 
    0.0006889228, 0.000691927, 0.0006917522, 0.000713242, 0.0007491158, 
    0.0008120902, 0.0008628415, 0.0008531618, 0.000790712, 0.0007219203, 
    0.000611993, 0.0004918145, 0.0004583562, 0.0005114763, 0.000526608, 
    0.0004927048, 0.0004461817, 0.0004194472, 0.0004093538, 0.0003991177, 
    0.000392442, 0.0004029961, 0.0004221967, 0.0004137249, 0.000384622, 
    0.0003542473, 0.0003328852, 0.0003202648,
  0.0005102844, 0.000529803, 0.0005502278, 0.0005836221, 0.0006067647, 
    0.0006338329, 0.0006137739, 0.0005677749, 0.0005625455, 0.0005684742, 
    0.0005056907, 0.0005084404, 0.0005480179, 0.0006316234, 0.0006855854, 
    0.0007177561, 0.000751993, 0.0008070358, 0.0008412568, 0.0008674987, 
    0.0008373151, 0.0007582713, 0.0006487103, 0.0005422168, 0.0004548443, 
    0.0003884051, 0.0003687432, 0.0003609706, 0.0003672489, 0.0003188497, 
    0.0002775553, 0.0002359753, 0.0002060935, 0.000210671, 0.0002336071, 
    0.0002909547, 0.0003718422, 0.0003864495, 0.0003692356, 0.0003938882, 
    0.0004861718, 0.000582668, 0.000686205, 0.0007527082, 0.0007195368, 
    0.0006641592, 0.0005776142, 0.0004145035, 8.365791e-005, -9.701634e-005, 
    -0.0001067754, -8.992711e-005, -9.116647e-005, -0.0001267227, 
    -0.0001778079, -0.0002017771, -0.0001880282, -0.0001120518, 
    1.694844e-005, 0.0001344888, 0.0002508527, 0.0003162113, 0.0003457116, 
    0.0003895808, 0.0004348801, 0.000478002, 0.0005259721, 0.0005505611, 
    0.0005629747, 0.0006118505, 0.0006500932, 0.0006286036, 0.0006254409, 
    0.000634898, 0.0006232951, 0.0005783292, 0.0005189627, 0.0005312487, 
    0.0005487329, 0.0005338397, 0.0005246534, 0.000501415, 0.000411992, 
    0.0003153528, 0.0003616693, 0.0004255818, 0.000479178, 0.0005132882, 
    0.0005211402, 0.0005326001, 0.0005508632, 0.0005541856, 0.00055684, 
    0.0005538358, 0.0005448394, 0.0005249552,
  0.0005064374, 0.0005579833, 0.0006155851, 0.0006060803, 0.0005576022, 
    0.0005537553, 0.0005724952, 0.0006051743, 0.0006239938, 0.0006043958, 
    0.0005834943, 0.0005648024, 0.0005694912, 0.000591696, 0.0006361692, 
    0.0006861414, 0.0007408031, 0.000807147, 0.0008398739, 0.0007567771, 
    0.0006283487, 0.0005731944, 0.0006019638, 0.000565883, 0.0005088057, 
    0.00050426, 0.0005281018, 0.0005528976, 0.0005538829, 0.0005377021, 
    0.0004950732, 0.0004330208, 0.0003883888, 0.0003903913, 0.0004405226, 
    0.0004907656, 0.0005455064, 0.0005831127, 0.0005828112, 0.0005582697, 
    0.0006080358, 0.0007449994, 0.0008521923, 0.0008383794, 0.00076536, 
    0.0007360661, 0.0006977282, 0.0006272201, 0.0004596598, 0.000322633, 
    0.0002347995, 0.0001728898, 0.0001396229, 0.0001214393, 9.867828e-005, 
    8.787028e-005, 0.0001079449, 0.000145488, 0.0002000541, 0.0002781758, 
    0.000354263, 0.0003972738, 0.0004248829, 0.0004307162, 0.0004195264, 
    0.0004168241, 0.0004463242, 0.000495391, 0.0005275141, 0.000568633, 
    0.0006018369, 0.0006073681, 0.0005941442, 0.0005696504, 0.0005147983, 
    0.0004644608, 0.0005153236, 0.0006378065, 0.000630511, 0.0005350481, 
    0.000545729, 0.0005621482, 0.0005752458, 0.0003826825, 0.0003451235, 
    0.0004243422, 0.0005103478, 0.0005389897, 0.0005458242, 0.0005573477, 
    0.0005753881, 0.0006214345, 0.0006056672, 0.0005593027, 0.0004978543, 
    0.0004806085,
  0.0005710809, 0.0005841302, 0.0006107856, 0.0006266325, 0.0006286509, 
    0.0006460713, 0.0006711211, 0.0006813258, 0.0006882239, 0.0006921822, 
    0.0006902586, 0.0006984121, 0.000706916, 0.0006946451, 0.0006965366, 
    0.0007329667, 0.0008165881, 0.0009131643, 0.0009500075, 0.0008869376, 
    0.0008321016, 0.0008801352, 0.0009370698, 0.0009246878, 0.0008905777, 
    0.0008825669, 0.0008925167, 0.0008908319, 0.0008854596, 0.0008678804, 
    0.0008210707, 0.0007450157, 0.0006835829, 0.0006814534, 0.0007122406, 
    0.0007223333, 0.0007197903, 0.0007020677, 0.0006724875, 0.0006923242, 
    0.0007910933, 0.0009032455, 0.0009242897, 0.000855498, 0.000869358, 
    0.0008635721, 0.0007975781, 0.0007196949, 0.000655862, 0.000529103, 
    0.0004268214, 0.000381792, 0.0003661043, 0.0003764359, 0.0003776751, 
    0.0003685676, 0.0003830795, 0.0004205275, 0.0004756176, 0.0005230312, 
    0.0005235556, 0.0005151159, 0.0005393708, 0.0005364148, 0.0004782085, 
    0.000431845, 0.00044154, 0.0004672892, 0.0004835492, 0.0004859334, 
    0.0004969332, 0.0005020979, 0.0004941509, 0.0004576091, 0.0004364853, 
    0.0005092346, 0.0006150771, 0.0006926898, 0.000628985, 0.0005895826, 
    0.0005296445, 0.0005293419, 0.000608942, 0.0005641193, 0.0005405319, 
    0.0005392763, 0.0005799027, 0.0006335629, 0.0006715986, 0.0007000652, 
    0.0006857598, 0.0006446089, 0.0006104514, 0.0005806016, 0.0005598911, 
    0.0005587148,
  0.0006478201, 0.0006916253, 0.0007444113, 0.0007781717, 0.0007824311, 
    0.0008196565, 0.0009016404, 0.0009847363, 0.001016303, 0.001024027, 
    0.001053639, 0.001088099, 0.001083696, 0.00103045, 0.0009827977, 
    0.0009594331, 0.0009694141, 0.001058551, 0.001121795, 0.001250525, 
    0.001518063, 0.00167224, 0.001623619, 0.001466867, 0.001357608, 
    0.001308239, 0.001247331, 0.00117811, 0.001131014, 0.001070456, 
    0.0009876932, 0.0009131473, 0.0008741585, 0.000853098, 0.0008278731, 
    0.0007752148, 0.0006974107, 0.0006410806, 0.0006432896, 0.0006735688, 
    0.0008338811, 0.001013267, 0.001048331, 0.0009664423, 0.001006322, 
    0.0009484175, 0.0009112242, 0.0008513969, 0.0007948447, 0.000712892, 
    0.0006844881, 0.0006781467, 0.0006814208, 0.0006903536, 0.0006825966, 
    0.0006667501, 0.0006764932, 0.0006645885, 0.0006507761, 0.0006911163, 
    0.0006970288, 0.0006391886, 0.0006144885, 0.0005925382, 0.0005434873, 
    0.0005251137, 0.0005092667, 0.0004667169, 0.0004713899, 0.0004897318, 
    0.0004742984, 0.0004567672, 0.0004467848, 0.0004409356, 0.000463347, 
    0.0005166419, 0.0005443306, 0.0005982448, 0.000574403, 0.0005879765, 
    0.0005400069, 0.0005588098, 0.0006444817, 0.0006098794, 0.0005493853, 
    0.0005445695, 0.0005906159, 0.0006450387, 0.0006828201, 0.0007067253, 
    0.0006739348, 0.0006349138, 0.00062889, 0.0006181924, 0.0005848934, 
    0.0006005499,
  0.0009235907, 0.0009869621, 0.001008038, 0.0009843074, 0.0009999797, 
    0.001141283, 0.001403861, 0.001603656, 0.001708925, 0.001820601, 
    0.001935073, 0.001940939, 0.001750363, 0.001546641, 0.00147386, 
    0.001416465, 0.001380178, 0.001422712, 0.001497766, 0.001577636, 
    0.00160124, 0.001539187, 0.00140038, 0.001220088, 0.001121255, 
    0.001066753, 0.001001426, 0.0009408044, 0.0008911015, 0.0008302894, 
    0.0008086567, 0.0008153482, 0.0007787589, 0.0007143542, 0.000635819, 
    0.0005895183, 0.0006043478, 0.0006942796, 0.000819338, 0.0008547031, 
    0.0009381021, 0.001072316, 0.00109158, 0.001081693, 0.001138437, 
    0.001218785, 0.001008276, 0.0009886785, 0.001028113, 0.001109875, 
    0.001143269, 0.001104503, 0.001015573, 0.0009547113, 0.0009164219, 
    0.0008373624, 0.0007676012, 0.0007412639, 0.0007419153, 0.0007875646, 
    0.0007825578, 0.000709109, 0.0006824536, 0.0006356924, 0.0005870545, 
    0.0005758968, 0.0005519912, 0.0005444889, 0.0005717482, 0.0005668844, 
    0.0005558217, 0.000557173, 0.0005620047, 0.0005693799, 0.0005408805, 
    0.0004895097, 0.0004836605, 0.0004720096, 0.0005396726, 0.0006530327, 
    0.0006441479, 0.0006163642, 0.0006398563, 0.0006875559, 0.0007198378, 
    0.0007254169, 0.0007709549, 0.0008538291, 0.0008967286, 0.000908236, 
    0.0008929139, 0.0008468353, 0.0008222149, 0.0008105482, 0.0008279048, 
    0.0008692625,
  0.001123624, 0.001107014, 0.001068152, 0.001053385, 0.001169607, 
    0.001401874, 0.001585901, 0.001709768, 0.00182424, 0.001865773, 
    0.001699834, 0.001538346, 0.001414289, 0.001326869, 0.001298052, 
    0.00126828, 0.001222424, 0.001191223, 0.001173008, 0.001148387, 
    0.001038809, 0.0008983808, 0.0008198787, 0.0007620696, 0.0007306621, 
    0.000726609, 0.0006897813, 0.0006753327, 0.0006903061, 0.000826681, 
    0.0009953068, 0.0009662989, 0.0008813906, 0.0007510865, 0.0006170948, 
    0.0006986507, 0.000853511, 0.0008719335, 0.0008711065, 0.0008768444, 
    0.001039541, 0.001212761, 0.00127885, 0.001244486, 0.001260316, 
    0.001299449, 0.001326819, 0.001091103, 0.001194339, 0.00119596, 
    0.001029909, 0.0009586224, 0.0009413129, 0.0008693105, 0.0008447212, 
    0.0007751347, 0.0007066294, 0.0007212525, 0.0007602735, 0.000801059, 
    0.0007623238, 0.0007101102, 0.0007460639, 0.0007806504, 0.0007966245, 
    0.0007811114, 0.0007423125, 0.0007784571, 0.0007826053, 0.0007474464, 
    0.0007532164, 0.0007415977, 0.0007194085, 0.0006913235, 0.00060918, 
    0.0005675042, 0.0005472549, 0.0005270843, 0.0006119297, 0.0006887638, 
    0.0007332214, 0.0007852442, 0.0009942101, 0.001190111, 0.001368988, 
    0.001373152, 0.001320844, 0.001336277, 0.001323561, 0.001266643, 
    0.001225794, 0.001197629, 0.001210837, 0.001181241, 0.001164664, 
    0.001161389,
  0.00111361, 0.001107618, 0.001070091, 0.001117806, 0.001307492, 
    0.001369941, 0.001515949, 0.001573012, 0.001743942, 0.001790959, 
    0.001429437, 0.00131819, 0.00139423, 0.001415338, 0.001382151, 
    0.001321561, 0.001222362, 0.001109686, 0.0009684293, 0.0008012503, 
    0.0006697392, 0.0006079553, 0.0006301757, 0.0006511733, 0.0006959643, 
    0.0007812865, 0.0008410024, 0.0009063929, 0.00105232, 0.001270219, 
    0.001111845, 0.00100106, 0.001015906, 0.001020467, 0.0009652181, 
    0.0009332383, 0.0009222077, 0.001007959, 0.001002634, 0.000986469, 
    0.0010898, 0.001486846, 0.00163732, 0.001570579, 0.001513517, 
    0.001478296, 0.001423395, 0.00129104, 0.001185945, 0.0009919694, 
    0.000810883, 0.0007848935, 0.0007736413, 0.0007144324, 0.0007084571, 
    0.0007160231, 0.0007524695, 0.0008292878, 0.0008606641, 0.0008954732, 
    0.0009226212, 0.0009304564, 0.0009414246, 0.0009295028, 0.000934653, 
    0.0009109387, 0.0009093489, 0.0009431094, 0.0009324281, 0.0009055501, 
    0.0008668778, 0.0007929206, 0.0007667905, 0.0007512299, 0.0006711055, 
    0.0006454675, 0.0006073359, 0.0006805463, 0.0008351691, 0.0009657904, 
    0.001043277, 0.001228734, 0.001524756, 0.001836195, 0.001799352, 
    0.001803404, 0.00178511, 0.001727015, 0.001554352, 0.001428308, 
    0.00137301, 0.001306267, 0.001267119, 0.001200124, 0.00115999, 0.001160547,
  0.001106632, 0.001110843, 0.001056246, 0.001119746, 0.00119952, 
    0.0008528912, 0.000833293, 0.001306284, 0.001894717, 0.002009921, 
    0.001934454, 0.001927668, 0.001975986, 0.001898549, 0.001802816, 
    0.001718607, 0.001564509, 0.001448161, 0.001304935, 0.00112113, 0.001096, 
    0.001105743, 0.001124927, 0.001179636, 0.001230292, 0.00126321, 
    0.0013533, 0.001441705, 0.001442977, 0.001351553, 0.001088705, 
    0.0009524231, 0.0007803012, 0.001151073, 0.001289976, 0.001417355, 
    0.001190874, 0.001183498, 0.00141869, 0.001506587, 0.001302151, 
    0.001560201, 0.001424588, 0.001485386, 0.00149125, 0.001475102, 
    0.001341651, 0.001162757, 0.001046902, 0.0009359894, 0.0009481171, 
    0.0009940034, 0.001010932, 0.000965219, 0.0009140382, 0.0009125443, 
    0.0009234799, 0.0009524552, 0.0009870101, 0.001029815, 0.001050223, 
    0.001092503, 0.001056248, 0.0009934166, 0.0009716088, 0.0009565251, 
    0.001003319, 0.0009918269, 0.0009724833, 0.0009434605, 0.0008666739, 
    0.0008530198, 0.0008151261, 0.0007415032, 0.000671884, 0.0006474378, 
    0.0006811824, 0.000868659, 0.001149786, 0.001267215, 0.00127033, 
    0.001538201, 0.001770439, 0.001986334, 0.002167755, 0.002017742, 
    0.001880414, 0.001715428, 0.001568991, 0.001408392, 0.001301565, 
    0.00119984, 0.001152394, 0.001120462, 0.001096905, 0.001126342,
  0.001101548, 0.001125278, 0.001177698, 0.001337551, 0.001400013, 
    0.00104644, 0.001295936, 0.00173264, 0.002095054, 0.002264695, 
    0.002289793, 0.002280764, 0.002308708, 0.002308866, 0.002223671, 
    0.002145678, 0.002064584, 0.001907005, 0.001780087, 0.001658843, 
    0.001593643, 0.001557197, 0.001568197, 0.001626863, 0.001661021, 
    0.001600558, 0.001551714, 0.001492109, 0.001388715, 0.00145215, 
    0.001330842, 0.001367192, 0.001484828, 0.001530381, 0.001416498, 
    0.001676118, 0.001615735, 0.001633744, 0.001721926, 0.002002799, 
    0.001721673, 0.001365523, 0.001171595, 0.001294889, 0.001343017, 
    0.001413845, 0.001409743, 0.001469173, 0.001492649, 0.001451991, 
    0.001451562, 0.001353826, 0.001266517, 0.001158991, 0.001073557, 
    0.001078357, 0.00101613, 0.0009849137, 0.001028717, 0.001053196, 
    0.001046743, 0.001027416, 0.0009699557, 0.0009885374, 0.00106046, 
    0.001110401, 0.001149374, 0.001118793, 0.001095444, 0.001053435, 
    0.000951821, 0.0009179488, 0.0007634545, 0.0007599723, 0.0006955191, 
    0.0007306151, 0.001086956, 0.0008495697, 0.001472191, 0.001581514, 
    0.001569643, 0.001816247, 0.001979995, 0.002132897, 0.002231444, 
    0.00203033, 0.00168413, 0.001548629, 0.00147928, 0.001292855, 0.00122187, 
    0.001203782, 0.001185025, 0.001121639, 0.001081155, 0.001094745,
  0.001274195, 0.001363189, 0.001514726, 0.001777052, 0.001266102, 
    0.00130541, 0.001908768, 0.002165069, 0.002368155, 0.002450646, 
    0.002663967, 0.002573051, 0.002691766, 0.002374177, 0.002351369, 
    0.002225435, 0.002211687, 0.002055651, 0.001843426, 0.001687198, 
    0.001590861, 0.001585663, 0.00164743, 0.001658907, 0.001648542, 
    0.001630454, 0.001564112, 0.001581133, 0.001590433, 0.001736551, 
    0.001799192, 0.001835732, 0.001690694, 0.00140073, 0.001475022, 
    0.001831933, 0.001787079, 0.002084006, 0.002094258, 0.002182871, 
    0.001758215, 0.001497003, 0.001526536, 0.001747963, 0.001763094, 
    0.0017822, 0.001763825, 0.00177856, 0.001769278, 0.001674625, 
    0.001580577, 0.001438638, 0.001356415, 0.001288419, 0.001226477, 
    0.001204861, 0.001160356, 0.001223346, 0.001268709, 0.001248603, 
    0.00126995, 0.001319222, 0.001392147, 0.001410522, 0.001420678, 
    0.001351727, 0.00128098, 0.001247316, 0.001179605, 0.001130204, 
    0.001072095, 0.001031245, 0.0009231782, 0.0008873846, 0.0007387381, 
    0.0010322, 0.001743753, 0.001177761, 0.001495286, 0.001870177, 
    0.001653471, 0.001999083, 0.002087837, 0.001875692, 0.00246228, 
    0.001958074, 0.001669555, 0.001460366, 0.00147669, 0.001381403, 
    0.001258585, 0.001188936, 0.001147753, 0.001103693, 0.001131398, 
    0.001161009,
  0.001555417, 0.001670764, 0.001890713, 0.002193345, 0.002008824, 
    0.002005978, 0.002597004, 0.002575864, 0.002392504, 0.002371588, 
    0.002824996, 0.002864, 0.002165148, 0.002145041, 0.002348126, 
    0.002227073, 0.002110232, 0.001987955, 0.001845079, 0.001732545, 
    0.001738665, 0.001783598, 0.001870303, 0.001921548, 0.001934184, 
    0.001890696, 0.001833699, 0.001854902, 0.00196308, 0.002158599, 
    0.002344788, 0.002096817, 0.001886229, 0.001579512, 0.002262024, 
    0.002216963, 0.002128955, 0.00244289, 0.002504704, 0.002193457, 
    0.001957151, 0.002000226, 0.002189243, 0.0022574, 0.002176845, 
    0.002048911, 0.001989704, 0.001900074, 0.001894908, 0.001893605, 
    0.001872735, 0.001766322, 0.001692872, 0.001670747, 0.001678043, 
    0.001669873, 0.001732943, 0.001853693, 0.0019136, 0.001970868, 
    0.002055061, 0.002118433, 0.002093859, 0.001945421, 0.001807981, 
    0.001723978, 0.001568926, 0.001502408, 0.001364919, 0.001313739, 
    0.001192844, 0.001148658, 0.001082093, 0.00106453, 0.001139599, 
    0.001445537, 0.002095577, 0.001857126, 0.002009937, 0.001905988, 
    0.001454215, 0.002907726, 0.003057263, 0.00273287, 0.002577851, 
    0.002341148, 0.001721609, 0.001631598, 0.001540125, 0.001411856, 
    0.0014082, 0.001345973, 0.001330713, 0.001296923, 0.00134216, 0.001395485,
  0.001997603, 0.002001164, 0.002205615, 0.002358807, 0.002287012, 
    0.001906956, 0.002445958, 0.002156963, 0.002332964, 0.002475188, 
    0.002366326, 0.002847359, 0.002617697, 0.002224816, 0.002262566, 
    0.002279462, 0.002194807, 0.002135282, 0.002079349, 0.002059002, 
    0.00215752, 0.002219062, 0.00229553, 0.002296373, 0.002269591, 
    0.002245367, 0.002279127, 0.002333407, 0.002545186, 0.002704356, 
    0.002828222, 0.002778423, 0.00269674, 0.003315598, 0.003234805, 
    0.002628603, 0.002427886, 0.002651808, 0.002862013, 0.002511013, 
    0.002520391, 0.002678224, 0.00272257, 0.002660948, 0.00255536, 
    0.002376926, 0.002303239, 0.002195857, 0.002265092, 0.002335109, 
    0.002293242, 0.002247561, 0.002263343, 0.002350606, 0.00243995, 
    0.002558632, 0.002727451, 0.002728308, 0.002802392, 0.002801646, 
    0.002806731, 0.002803362, 0.00264882, 0.002459404, 0.00227997, 
    0.002199687, 0.002019522, 0.001933993, 0.001791704, 0.001690425, 
    0.001595661, 0.001648557, 0.001659859, 0.001667695, 0.00166609, 
    0.001840326, 0.002281226, 0.00246681, 0.002081956, 0.001896624, 
    0.001718065, 0.002713813, 0.002940628, 0.002483754, 0.002460103, 
    0.002015707, 0.001852883, 0.001850181, 0.001826053, 0.00171948, 
    0.001754464, 0.001686896, 0.00172792, 0.001728762, 0.001809173, 0.00187558,
  0.002341704, 0.00238125, 0.002550242, 0.002676381, 0.002485614, 
    0.001840724, 0.002662443, 0.002080558, 0.002152099, 0.002085771, 
    0.002119832, 0.002641857, 0.002537367, 0.002305449, 0.002443064, 
    0.002408637, 0.002507692, 0.002519852, 0.002506848, 0.002536874, 
    0.00260433, 0.002623452, 0.002677526, 0.002647452, 0.002692578, 
    0.002744298, 0.002811581, 0.002916358, 0.003083568, 0.003123637, 
    0.003127929, 0.003244739, 0.003395325, 0.003360737, 0.003305981, 
    0.003543302, 0.003261556, 0.003135448, 0.002945142, 0.002942869, 
    0.003124703, 0.003151167, 0.003115818, 0.003026586, 0.002919264, 
    0.00280376, 0.002761589, 0.002764054, 0.002792316, 0.002762465, 
    0.002744598, 0.002760636, 0.00288827, 0.003098095, 0.003279643, 
    0.003324067, 0.003406579, 0.003384579, 0.003374724, 0.003293216, 
    0.003185198, 0.003075192, 0.00285885, 0.002747048, 0.002599547, 
    0.002520582, 0.002394761, 0.002324013, 0.00224184, 0.002189261, 
    0.002227343, 0.002174732, 0.002062199, 0.002000703, 0.002083656, 
    0.002811389, 0.003036044, 0.002178357, 0.001314248, 0.0008986536, 
    0.001172788, 0.001150295, 0.002002053, 0.002487552, 0.00214935, 
    0.001816086, 0.002131864, 0.002127064, 0.002136824, 0.002136092, 
    0.002146981, 0.002142292, 0.002200275, 0.002239661, 0.002348619, 
    0.00233719,
  0.002718231, 0.002727292, 0.002762307, 0.002937863, 0.00234722, 
    0.002851015, 0.002934397, 0.002727053, 0.002215042, 0.002363545, 
    0.002242093, 0.002578931, 0.0025432, 0.002514176, 0.002600975, 
    0.002682641, 0.002820892, 0.002840808, 0.002946205, 0.002928674, 
    0.002987104, 0.002957365, 0.002958873, 0.002962068, 0.003020244, 
    0.003067624, 0.003125148, 0.003224153, 0.003224362, 0.00330512, 
    0.003428403, 0.003370354, 0.003510224, 0.003510384, 0.003519172, 
    0.003442483, 0.003343858, 0.003408054, 0.003199931, 0.003268817, 
    0.003394974, 0.003370656, 0.003310667, 0.00323269, 0.003110984, 
    0.003007878, 0.002929438, 0.002897188, 0.002883263, 0.002903117, 
    0.003053891, 0.003140979, 0.003304295, 0.003499702, 0.003632311, 
    0.003624316, 0.003578508, 0.003471473, 0.003353029, 0.003313052, 
    0.003249792, 0.00316792, 0.003098445, 0.002987692, 0.002873074, 
    0.002789199, 0.002701781, 0.002654828, 0.002592823, 0.002579487, 
    0.00258656, 0.002446228, 0.002426581, 0.002408065, 0.002634069, 
    0.003283728, 0.002177086, 0.001464563, 0.001940224, 0.001981264, 
    0.001173279, 0.001311865, 0.001324881, 0.002639505, 0.00252934, 
    0.002184667, 0.002188926, 0.002444081, 0.002557377, 0.002592616, 
    0.002597623, 0.002625343, 0.002647199, 0.002709202, 0.002744997, 
    0.002681753,
  0.003022613, 0.003040317, 0.003051843, 0.003012422, 0.00248927, 
    0.003270821, 0.003254467, 0.003251733, 0.00299424, 0.002305545, 
    0.002442795, 0.002499316, 0.002594966, 0.002693625, 0.00281927, 
    0.00297267, 0.003120538, 0.003153695, 0.00323757, 0.003126148, 
    0.003091801, 0.003092214, 0.003188932, 0.003301673, 0.003359511, 
    0.003289163, 0.00330911, 0.00330792, 0.003270393, 0.003354235, 
    0.003416495, 0.003371846, 0.003407052, 0.003411457, 0.003404448, 
    0.003309509, 0.003185371, 0.002926895, 0.002800009, 0.003044293, 
    0.003533861, 0.003349356, 0.003140643, 0.003028763, 0.002841843, 
    0.00274797, 0.002673708, 0.002711823, 0.002989534, 0.003238332, 
    0.003501913, 0.003674526, 0.003819248, 0.003838081, 0.003754651, 
    0.003638303, 0.003457105, 0.003332015, 0.003267135, 0.003251303, 
    0.003204303, 0.003143298, 0.003147941, 0.003036058, 0.002994208, 
    0.002898254, 0.002888177, 0.002864907, 0.002812183, 0.002789311, 
    0.00275172, 0.002716165, 0.002773736, 0.002721679, 0.002978027, 
    0.003370416, 0.001765654, 0.002532312, 0.003957547, 0.004198668, 
    0.00237216, 0.00123012, 0.001522595, 0.001802465, 0.002835326, 
    0.002555947, 0.00265683, 0.002768792, 0.00303237, 0.003042623, 
    0.003058614, 0.003043545, 0.003086478, 0.003083393, 0.003012503, 
    0.002993828,
  0.003299782, 0.003333636, 0.003253225, 0.002732902, 0.003147146, 
    0.002568091, 0.003104245, 0.003013601, 0.002914498, 0.002726782, 
    0.002718756, 0.00269749, 0.002718912, 0.002905771, 0.003003793, 
    0.003124112, 0.003236774, 0.003186293, 0.003141979, 0.00316358, 
    0.003069421, 0.00305526, 0.003195608, 0.003272552, 0.003432818, 
    0.003333159, 0.003330346, 0.00309827, 0.003237046, 0.003559452, 
    0.003432709, 0.003385136, 0.003249792, 0.003482871, 0.00353599, 
    0.003106186, 0.00280139, 0.002673598, 0.002814012, 0.003397262, 
    0.003493296, 0.003119633, 0.00298235, 0.00292176, 0.002905564, 
    0.003024915, 0.003184242, 0.00339642, 0.00379299, 0.003931606, 
    0.003889231, 0.003730427, 0.00355999, 0.003395183, 0.003277658, 
    0.003233548, 0.003204398, 0.003172005, 0.003144046, 0.003099445, 
    0.003117964, 0.003071742, 0.00307144, 0.003009627, 0.003026379, 
    0.003011581, 0.00307516, 0.00299014, 0.003015604, 0.002952915, 
    0.002943996, 0.002946477, 0.002863459, 0.002829174, 0.002810609, 
    0.003149007, 0.002247021, 0.002910491, 0.003746608, 0.004665252, 
    0.003282632, 0.001786603, 0.001649941, 0.002003357, 0.002470769, 
    0.002950944, 0.003076686, 0.003230147, 0.003367029, 0.003343999, 
    0.003407419, 0.003318934, 0.003316997, 0.00326103, 0.003203478, 
    0.003308967,
  0.003351945, 0.00346154, 0.003200853, 0.002831877, 0.002974737, 
    0.003336385, 0.003356287, 0.003013775, 0.003354426, 0.003419737, 
    0.002964359, 0.002533982, 0.00257216, 0.002921347, 0.003151469, 
    0.003348291, 0.003456231, 0.00335112, 0.003181444, 0.003109459, 
    0.00304763, 0.003021833, 0.003129406, 0.003079737, 0.003169954, 
    0.003154712, 0.003049854, 0.002852729, 0.003373833, 0.003528552, 
    0.00347149, 0.003233262, 0.002899237, 0.003124606, 0.003100511, 
    0.002830828, 0.002785908, 0.002867846, 0.003189266, 0.003415033, 
    0.003259266, 0.002983829, 0.003030591, 0.003029637, 0.003126863, 
    0.003361482, 0.00363053, 0.003904171, 0.004142653, 0.004201958, 
    0.004111532, 0.003931163, 0.003789796, 0.003588682, 0.003473271, 
    0.003341058, 0.003299732, 0.003203094, 0.003201218, 0.003190888, 
    0.003203047, 0.003170399, 0.003187884, 0.003140088, 0.00313993, 
    0.003149958, 0.003190838, 0.003188536, 0.003215667, 0.003074842, 
    0.003022643, 0.002933554, 0.002706692, 0.002698027, 0.002412956, 
    0.002738973, 0.003068818, 0.003077097, 0.003366904, 0.003472953, 
    0.003265751, 0.001356607, 0.001527537, 0.003074061, 0.00302935, 
    0.003107583, 0.003201965, 0.003279833, 0.003369685, 0.003374454, 
    0.003355602, 0.003283236, 0.00333246, 0.003329713, 0.003296984, 
    0.003243895,
  0.003089607, 0.003492964, 0.003141312, 0.003081566, 0.003193511, 
    0.003368018, 0.003439162, 0.003223313, 0.003495537, 0.003737677, 
    0.003271711, 0.003091912, 0.002468353, 0.002947813, 0.003193397, 
    0.003340136, 0.00356115, 0.003678773, 0.003581353, 0.003379349, 
    0.003249712, 0.003023358, 0.003006, 0.003037028, 0.003102545, 
    0.003073284, 0.002783256, 0.003011104, 0.003232975, 0.003193827, 
    0.003203634, 0.003055243, 0.002825312, 0.002945459, 0.003027093, 
    0.002929119, 0.002961513, 0.003104405, 0.00324237, 0.003208783, 
    0.003115276, 0.002985228, 0.002842097, 0.002814535, 0.002834355, 
    0.0028324, 0.00288978, 0.00292737, 0.003080228, 0.003235757, 0.003425999, 
    0.003497619, 0.003617354, 0.003569147, 0.003555637, 0.003501054, 
    0.003483936, 0.003438715, 0.003533335, 0.003506346, 0.003497986, 
    0.003463462, 0.003406417, 0.003379969, 0.00342565, 0.00342975, 
    0.003367048, 0.003375407, 0.00332124, 0.003326721, 0.003174707, 
    0.00302037, 0.002898648, 0.002933379, 0.002788421, 0.002991378, 
    0.002976343, 0.002867592, 0.002886681, 0.002234002, 0.002397032, 
    0.002701622, 0.003135892, 0.003164789, 0.003180778, 0.003336625, 
    0.003279753, 0.003179125, 0.003015984, 0.003049012, 0.003077019, 
    0.003133254, 0.003155267, 0.003153296, 0.003044799, 0.002981825,
  0.003144601, 0.003151532, 0.003259234, 0.003151771, 0.002993984, 
    0.003214667, 0.003432754, 0.003564857, 0.003824873, 0.003607627, 
    0.003091675, 0.003207848, 0.002858452, 0.00230629, 0.00301379, 
    0.003219465, 0.003466355, 0.003488973, 0.003442196, 0.003365982, 
    0.003212089, 0.003040254, 0.002971113, 0.002890639, 0.002904579, 
    0.003070723, 0.003114052, 0.00312157, 0.003031719, 0.003072791, 
    0.003139835, 0.003321873, 0.003255052, 0.002889367, 0.003051618, 
    0.003079498, 0.003112225, 0.003082486, 0.003067115, 0.003006224, 
    0.002964532, 0.002968807, 0.002828697, 0.002865858, 0.0028516, 
    0.002756361, 0.002756346, 0.002696184, 0.002764577, 0.002710871, 
    0.00275032, 0.0027408, 0.00286462, 0.002907805, 0.002958413, 0.002981922, 
    0.003075397, 0.003152678, 0.003276734, 0.003221231, 0.003280327, 
    0.003285889, 0.003352487, 0.003375933, 0.003380667, 0.003437795, 
    0.003455436, 0.003463097, 0.00352186, 0.003667263, 0.003423281, 
    0.003300829, 0.003139865, 0.00296369, 0.002914291, 0.002918486, 
    0.002695294, 0.0024866, 0.003128309, 0.002837596, 0.002998468, 
    0.00302347, 0.00311685, 0.003061106, 0.003103402, 0.003277417, 
    0.003210086, 0.00315382, 0.003005017, 0.003140248, 0.003107727, 
    0.003154457, 0.003206225, 0.003082296, 0.003163755, 0.003182545,
  0.003145745, 0.003140341, 0.003185388, 0.002842924, 0.002116065, 
    0.001957151, 0.002174972, 0.002699667, 0.003184147, 0.002776962, 
    0.002880975, 0.002154022, 0.002995973, 0.002641618, 0.003355509, 
    0.003111733, 0.00323269, 0.003317963, 0.003279928, 0.003368476, 
    0.003030909, 0.003010087, 0.003260076, 0.003121538, 0.003003618, 
    0.003062697, 0.003185928, 0.002923222, 0.002607094, 0.002924096, 
    0.00319211, 0.003395688, 0.003426461, 0.003104452, 0.003282456, 
    0.003185373, 0.003160767, 0.003068959, 0.002947971, 0.002981888, 
    0.00290186, 0.002913987, 0.002872169, 0.002858482, 0.00289838, 0.0029453, 
    0.003025852, 0.003007321, 0.003000963, 0.002927942, 0.002976961, 
    0.003012709, 0.003055036, 0.003071535, 0.00309056, 0.003096966, 
    0.00314565, 0.003124209, 0.003223946, 0.003222469, 0.003316978, 
    0.003447456, 0.003500244, 0.003470935, 0.003429146, 0.00352639, 
    0.003589284, 0.003689278, 0.003734943, 0.003644869, 0.003629815, 
    0.00340753, 0.002815519, 0.002390958, 0.002426932, 0.002510933, 
    0.00256728, 0.002733488, 0.002760049, 0.002858087, 0.002802121, 
    0.002676301, 0.002771428, 0.00272241, 0.002772652, 0.002765005, 
    0.002807094, 0.002914799, 0.002951769, 0.003081962, 0.003067385, 
    0.003098587, 0.003292389, 0.003203586, 0.003236253, 0.003205812,
  0.002436452, 0.001939603, 0.00164069, 0.001701186, 0.0009065513, 
    0.00112534, 0.001292679, 0.001148006, 0.001129633, 0.001614369, 
    0.002677684, 0.003512531, 0.002822673, 0.003172958, 0.003072108, 
    0.003414858, 0.003091974, 0.003293216, 0.003264796, 0.003355857, 
    0.003119888, 0.003085444, 0.003362929, 0.003291484, 0.003233772, 
    0.003244197, 0.003119774, 0.003027443, 0.002869023, 0.003293836, 
    0.003443355, 0.003609041, 0.003612714, 0.003529649, 0.003527932, 
    0.003388107, 0.003189312, 0.003095154, 0.002915926, 0.002852872, 
    0.002809402, 0.002710029, 0.002702653, 0.002747493, 0.002797719, 
    0.002829699, 0.002874855, 0.002837075, 0.002811054, 0.002911, 
    0.003039714, 0.003111668, 0.003155109, 0.003103817, 0.003139755, 
    0.003151134, 0.003197948, 0.003182702, 0.003224187, 0.003277894, 
    0.003413206, 0.003554875, 0.003471332, 0.003355825, 0.003269771, 
    0.003335496, 0.003571704, 0.003637033, 0.003607595, 0.00295455, 
    0.003050236, 0.002753263, 0.002054458, 0.002617586, 0.002756711, 
    0.002719136, 0.002654398, 0.002635991, 0.002745949, 0.002705261, 
    0.002647564, 0.002651744, 0.002623688, 0.002625899, 0.002651647, 
    0.002566611, 0.002612658, 0.002564784, 0.002634609, 0.002625151, 
    0.002763148, 0.002734236, 0.002551829, 0.002237372, 0.002351734, 
    0.002410863,
  0.00141424, 0.001490868, 0.001235235, 0.001565381, 0.0006139958, 
    0.001320541, 0.001070186, 0.001085763, 0.001010613, 0.001383342, 
    0.003417956, 0.002697902, 0.0018508, 0.002217981, 0.003372737, 
    0.004734663, 0.003315372, 0.003056277, 0.003311891, 0.003395038, 
    0.003294693, 0.003300877, 0.003309285, 0.003353473, 0.003364868, 
    0.003097475, 0.00289806, 0.002759685, 0.002906073, 0.003354777, 
    0.003536593, 0.003639624, 0.003726948, 0.003751999, 0.003654325, 
    0.003543206, 0.003246279, 0.002967108, 0.002721138, 0.002641793, 
    0.002685027, 0.002649836, 0.002732789, 0.002845926, 0.002881294, 
    0.002869975, 0.002819987, 0.002818732, 0.002811708, 0.002850903, 
    0.002903068, 0.002929404, 0.002924049, 0.002837328, 0.00283221, 
    0.002794618, 0.00282409, 0.002836963, 0.002814695, 0.002860917, 
    0.002919821, 0.002957761, 0.002849139, 0.002576372, 0.002215007, 
    0.002251025, 0.002852205, 0.003270391, 0.002883121, 0.002555598, 0.00277, 
    0.00225856, 0.001745561, 0.002877543, 0.002901668, 0.002768727, 
    0.002768138, 0.002696311, 0.002691463, 0.002656607, 0.00262698, 
    0.002618492, 0.002652092, 0.002633305, 0.002565548, 0.002493974, 
    0.002457274, 0.002409972, 0.002451567, 0.002288266, 0.00235609, 
    0.002373461, 0.001409155, 0.0009822571, 0.0007938431, 0.0009540441,
  0.00141664, 0.00153089, 0.0009507379, 0.0009165339, 0.0009411541, 
    0.001017957, 0.0004575776, 0.001045614, 0.001143461, 0.001612254, 
    0.003105026, 0.002076392, 0.001923995, 0.002101473, 0.002976787, 
    0.004912112, 0.003884908, 0.003522431, 0.003818087, 0.003658997, 
    0.003665959, 0.003730984, 0.003484206, 0.003252702, 0.003153075, 
    0.003118502, 0.002842431, 0.002490683, 0.002411037, 0.003017399, 
    0.003323131, 0.003357908, 0.003527679, 0.003693411, 0.003588507, 
    0.003472826, 0.003155459, 0.002814408, 0.002704814, 0.002723761, 
    0.002832402, 0.002849344, 0.00287403, 0.002867607, 0.002854845, 
    0.002878178, 0.002840761, 0.002833497, 0.002785048, 0.002753738, 
    0.002757316, 0.002686042, 0.00261749, 0.002553277, 0.002520995, 
    0.002483802, 0.002456463, 0.002428695, 0.002389929, 0.002412214, 
    0.002441824, 0.002488983, 0.002465952, 0.002061673, 0.001655154, 
    0.001634171, 0.002046335, 0.003074443, 0.002552148, 0.00254277, 
    0.002840493, 0.00283682, 0.002562989, 0.002940342, 0.003015904, 
    0.002835961, 0.002723714, 0.002799816, 0.002795827, 0.002723381, 
    0.002720978, 0.002681626, 0.002643747, 0.002604444, 0.002589883, 
    0.002505356, 0.002424246, 0.002391677, 0.002334647, 0.002225786, 
    0.002120928, 0.002071115, 0.001313247, 0.001425573, 0.001534863, 
    0.001063781,
  0.000596941, 0.001313054, 0.001409885, 0.001097954, 0.001700406, 
    0.00169869, 0.0009828131, 0.000774595, 0.001138405, 0.001387028, 
    0.00174615, 0.001205751, 0.001644759, 0.001652452, 0.002492513, 
    0.003100655, 0.00297191, 0.003323847, 0.004402722, 0.004360618, 
    0.003883859, 0.003563869, 0.003052605, 0.002642716, 0.00263647, 
    0.002733109, 0.002525318, 0.00220579, 0.002087328, 0.0024986, 
    0.002908155, 0.003072823, 0.003233676, 0.003480598, 0.003585724, 
    0.003508843, 0.003330171, 0.003092483, 0.002902035, 0.002856003, 
    0.002945714, 0.002942408, 0.002947779, 0.002999105, 0.002931884, 
    0.002880752, 0.002860805, 0.002816839, 0.002699126, 0.002580617, 
    0.00252524, 0.002462121, 0.00245125, 0.002423737, 0.002348793, 
    0.002265744, 0.002183745, 0.002113173, 0.002047544, 0.002054251, 
    0.002065298, 0.002065234, 0.002063359, 0.001856046, 0.001698054, 
    0.00165447, 0.00173798, 0.002825106, 0.002538749, 0.002856974, 
    0.002951132, 0.003077177, 0.002863126, 0.002953645, 0.002492925, 
    0.002670102, 0.00280457, 0.002942709, 0.002934635, 0.00290898, 
    0.002847327, 0.002720948, 0.002613898, 0.002592282, 0.002617905, 
    0.002467781, 0.002374066, 0.002350907, 0.0022488, 0.002238103, 
    0.002081764, 0.002047227, 0.002261913, 0.001674579, 0.00143236, 
    0.0002890793,
  0.0009103497, 0.0005953675, -8.244067e-006, 0.001518603, 0.001814291, 
    0.002141226, 0.001622222, 0.001138772, 0.00254792, 0.002074788, 
    0.001656569, 0.001302453, 0.00178301, 0.002148173, 0.00138563, 
    0.001245392, 0.001332415, 0.001699786, 0.002670835, 0.003563901, 
    0.003463481, 0.002431492, 0.002074946, 0.002028868, 0.002137061, 
    0.002119261, 0.00207946, 0.002069606, 0.002196938, 0.00222318, 
    0.002388911, 0.002669212, 0.00286977, 0.002961719, 0.003102593, 
    0.003247136, 0.003258375, 0.003108634, 0.002945762, 0.002871899, 
    0.002943091, 0.002899809, 0.002871787, 0.002873456, 0.002845149, 
    0.002830289, 0.002832735, 0.00273759, 0.002610481, 0.002457863, 
    0.002360475, 0.002289475, 0.002224736, 0.002267064, 0.002305385, 
    0.002282593, 0.002198081, 0.00209909, 0.001991611, 0.001958979, 
    0.001923963, 0.001882701, 0.001926824, 0.001993756, 0.002018186, 
    0.002579695, 0.002534776, 0.002528926, 0.002718915, 0.003130219, 
    0.003024725, 0.002508645, 0.002484406, 0.002523475, 0.002429982, 
    0.002469081, 0.002491031, 0.00254827, 0.002686091, 0.00276299, 
    0.002765516, 0.002699666, 0.002587466, 0.002448754, 0.002464442, 
    0.002447466, 0.002367359, 0.002308214, 0.002250214, 0.00221469, 
    0.002059703, 0.001948203, 0.002026976, 0.002436785, 0.002576421, 
    0.001337771,
  0.002637138, 0.002317895, 0.001992119, 0.00246166, 0.002343739, 0.00225357, 
    0.002095131, 0.001978435, 0.00227819, 0.002335061, 0.001920753, 
    0.00186323, 0.001887946, 0.002039421, 0.001763316, 0.001402414, 
    0.001559214, 0.00137115, 0.001356415, 0.001514328, 0.001385137, 
    0.001509194, 0.001595072, 0.00145342, 0.001533147, 0.001582738, 
    0.001592545, 0.001976844, 0.002197939, 0.002022479, 0.001833079, 
    0.002066603, 0.002284867, 0.002433496, 0.002518786, 0.002732632, 
    0.002607811, 0.002583969, 0.002629556, 0.002639107, 0.002582474, 
    0.002551878, 0.00255768, 0.002638695, 0.002734253, 0.002796051, 
    0.002781746, 0.002709122, 0.00260395, 0.002415248, 0.00226754, 
    0.002184953, 0.002110598, 0.00206595, 0.00211368, 0.002194108, 
    0.002149921, 0.002072324, 0.002000337, 0.001923995, 0.001848242, 
    0.001792516, 0.001901091, 0.002043602, 0.002563244, 0.002288236, 
    0.002398942, 0.002288443, 0.002798229, 0.003176471, 0.002911764, 
    0.002442031, 0.002273104, 0.002397701, 0.002330611, 0.002202215, 
    0.002266999, 0.002275662, 0.002326382, 0.002402151, 0.00243097, 
    0.002404964, 0.002421463, 0.002338286, 0.002319912, 0.002253997, 
    0.002071593, 0.002096165, 0.002156707, 0.002109597, 0.002056143, 
    0.001907544, 0.001761806, 0.00201798, 0.002211845, 0.002661917,
  0.002853526, 0.002662361, 0.002647119, 0.002686537, 0.002473392, 
    0.002109834, 0.0017702, 0.001165905, 0.001338534, 0.001225444, 
    0.001421948, 0.001769547, 0.002182774, 0.002231223, 0.001784329, 
    0.001178126, 0.0005092991, 0.0006147912, 0.001427289, 0.001364458, 
    0.001299831, 0.0008367109, 0.0004148372, 0.0006343727, 0.001115739, 
    0.001224856, 0.001349883, 0.001726521, 0.00193555, 0.001927651, 
    0.001794676, 0.001727474, 0.001803405, 0.001851643, 0.001938078, 
    0.002271483, 0.00219781, 0.001825036, 0.002063232, 0.002087423, 
    0.002118227, 0.002157279, 0.002179373, 0.002260944, 0.002329689, 
    0.002390008, 0.002363877, 0.002297295, 0.002201148, 0.00205751, 
    0.001944167, 0.001910564, 0.001877631, 0.001795233, 0.001771201, 
    0.001817359, 0.001872623, 0.001922628, 0.001906908, 0.001862181, 
    0.00179463, 0.001747169, 0.001851804, 0.002242714, 0.002214023, 
    0.001914935, 0.001916382, 0.002000829, 0.002467003, 0.002990379, 
    0.002878655, 0.002512078, 0.002336126, 0.002124649, 0.00209971, 
    0.002127334, 0.002187289, 0.002623309, 0.002563704, 0.002452538, 
    0.002323266, 0.002305512, 0.0023706, 0.002320549, 0.002130927, 
    0.001851612, 0.001588508, 0.001543702, 0.001688518, 0.001761473, 
    0.001851849, 0.001835288, 0.001734913, 0.001611063, 0.001724456, 
    0.002188037,
  0.002054665, 0.002256446, 0.002272452, 0.002139621, 0.002099504, 
    0.001694001, 0.00122759, 0.001049602, 0.001233678, 0.001353873, 
    0.001015811, 0.001396804, 0.001597615, 0.001562935, 0.001058901, 
    0.0006630151, 0.0005575544, 0.0001500018, 0.0006553703, 0.0009717187, 
    0.001149405, 0.00112774, 0.001189109, 0.001234186, 0.0009865814, 
    0.0008403824, 0.0008588203, 0.0009273582, 0.001279931, 0.001582627, 
    0.001631726, 0.001635905, 0.001573599, 0.001437128, 0.001444026, 
    0.001539251, 0.00161742, 0.001677885, 0.001484382, 0.001733944, 
    0.001669538, 0.001624286, 0.001578367, 0.001568035, 0.001580005, 
    0.00161963, 0.001648033, 0.001622538, 0.001603225, 0.001622713, 
    0.001609092, 0.001589225, 0.001553064, 0.001459923, 0.001398379, 
    0.00140229, 0.001468172, 0.00155637, 0.00161952, 0.001661959, 
    0.001675088, 0.001638275, 0.001717097, 0.001676882, 0.001800017, 
    0.00192986, 0.00173779, 0.001963524, 0.002222638, 0.002504275, 
    0.002562847, 0.002374194, 0.002377166, 0.002284326, 0.00242156, 
    0.001980645, 0.002167008, 0.002270673, 0.002479988, 0.002449741, 
    0.0022437, 0.002018394, 0.001924505, 0.001761521, 0.001604356, 
    0.001426114, 0.001127169, 0.0009492608, 0.001056216, 0.001322577, 
    0.001555337, 0.001643408, 0.001622825, 0.001559342, 0.001405865, 
    0.001318475,
  0.001432631, 0.001466867, 0.001459444, 0.001489405, 0.001565731, 
    0.001283475, 0.001083188, 0.001177061, 0.001285573, 0.001245122, 
    0.001200458, 0.001234139, 0.001216162, 0.0009800005, 0.001270252, 
    0.001012584, 0.0009809854, 0.0007516108, 0.0008653528, 0.001031849, 
    0.001006036, 0.0008898941, 0.0009985175, 0.0008652089, 0.0007956075, 
    0.001078626, 0.001111559, 0.001163694, 0.001344733, 0.001411824, 
    0.001367812, 0.001331032, 0.001363806, 0.001281346, 0.001194354, 
    0.001221677, 0.001296048, 0.001515282, 0.001559183, 0.001468393, 
    0.001244247, 0.001249446, 0.001246409, 0.001241943, 0.001258759, 
    0.001274527, 0.001285811, 0.001287353, 0.001320812, 0.00136565, 
    0.001373359, 0.00135516, 0.001347737, 0.001328186, 0.001309749, 
    0.00129422, 0.001330064, 0.001384884, 0.001388254, 0.001428085, 
    0.001488183, 0.001543783, 0.001617819, 0.001661988, 0.001609393, 
    0.001749981, 0.001749917, 0.0019256, 0.002001147, 0.00202793, 
    0.001483429, 0.00184875, 0.0019098, 0.002011415, 0.001924233, 
    0.001909245, 0.001916095, 0.00199959, 0.002021539, 0.002061245, 
    0.001848035, 0.001544257, 0.001028542, 0.0008928184, 0.0009769327, 
    0.001093074, 0.0009193793, 0.000682964, 0.0006760657, 0.0007735314, 
    0.001028989, 0.001266723, 0.00132083, 0.001345243, 0.001433458, 0.00148634,
  0.001146876, 0.001126278, 0.001281425, 0.001304599, 0.001319969, 
    0.001276911, 0.001133366, 0.000936544, 0.0007560616, 0.0007336661, 
    0.0007662182, 0.0007485435, 0.0008907202, 0.001108921, 0.001047091, 
    0.0009560948, 0.0009856108, 0.001178539, 0.001164075, 0.00113494, 
    0.001228496, 0.001177109, 0.001063574, 0.00105213, 0.0009659012, 
    0.0008728714, 0.0009916979, 0.001116439, 0.001197009, 0.001237921, 
    0.001249604, 0.001168526, 0.001125197, 0.001089164, 0.001074652, 
    0.001120938, 0.001154634, 0.00106839, 0.0009892983, 0.001067071, 
    0.001217831, 0.001296509, 0.001277992, 0.001257392, 0.001282951, 
    0.001305521, 0.001302787, 0.001293759, 0.001285064, 0.001271316, 
    0.001262224, 0.001278866, 0.001305727, 0.001310226, 0.001314072, 
    0.001295126, 0.001296445, 0.001338613, 0.001360294, 0.001379495, 
    0.001409918, 0.001462227, 0.001405466, 0.001346831, 0.001317744, 
    0.001379001, 0.001427273, 0.001497782, 0.001333019, 0.001320287, 
    0.001421742, 0.001502789, 0.00157452, 0.001617182, 0.001649352, 
    0.001635492, 0.001586426, 0.00155327, 0.00150778, 0.001490216, 
    0.001514328, 0.001476197, 0.0009387378, 0.0009096507, 0.0009596394, 
    0.0008979524, 0.0006482485, 0.00031556, 0.0001560096, 0.0002097022, 
    0.000468052, 0.0008027134, 0.0009863125, 0.001058266, 0.001174234, 
    0.001249494,
  0.001109477, 0.001159164, 0.001095696, 0.001103978, 0.001110844, 
    0.001164743, 0.001118489, 0.001003906, 0.0009268327, 0.000941488, 
    0.0009239563, 0.0008795308, 0.0008459613, 0.0009430931, 0.0009830045, 
    0.001004144, 0.001030704, 0.001020881, 0.001036251, 0.001008483, 
    0.001018354, 0.001055849, 0.001062032, 0.0009759157, 0.001022518, 
    0.001103357, 0.001145208, 0.001208341, 0.001232501, 0.001193591, 
    0.001131602, 0.001108157, 0.001076734, 0.001015572, 0.0009849593, 
    0.001033342, 0.001078832, 0.001051065, 0.0008911653, 0.0009651864, 
    0.001184007, 0.001307587, 0.001213348, 0.001201857, 0.001211409, 
    0.001272953, 0.001265403, 0.001236252, 0.001218307, 0.001196882, 
    0.001181686, 0.001221264, 0.001287338, 0.001330921, 0.001344685, 
    0.001319588, 0.001313976, 0.001343033, 0.001368496, 0.001394753, 
    0.001361073, 0.001320636, 0.001264863, 0.001207372, 0.001208358, 
    0.001232581, 0.001282204, 0.001282379, 0.001283952, 0.001322512, 
    0.001289038, 0.001329649, 0.001405164, 0.001408248, 0.001402509, 
    0.001313039, 0.001360278, 0.001330093, 0.001260031, 0.001179699, 
    0.001119682, 0.000816429, 0.0007466841, 0.0006756033, 0.0006309235, 
    0.0006343252, 0.0005470002, 0.0003593969, 0.0001853672, 0.0001976374, 
    0.0004163785, 0.0006978558, 0.0008716937, 0.0009663152, 0.001045136, 
    0.001086541,
  0.0008436246, 0.0009822734, 0.0009164689, 0.0008865083, 0.0008386499, 
    0.001043626, 0.001023996, 0.0009229705, 0.0008604731, 0.0008340403, 
    0.0009244327, 0.0009839102, 0.001075082, 0.001156318, 0.001238128, 
    0.001295507, 0.001233201, 0.001266214, 0.001236507, 0.001207118, 
    0.001190254, 0.001183006, 0.001159673, 0.001177125, 0.001177951, 
    0.001200235, 0.001211552, 0.001248952, 0.001214969, 0.001153314, 
    0.001084635, 0.001042418, 0.001000171, 0.0009456049, 0.0008974285, 
    0.0008928343, 0.0009210319, 0.0009513106, 0.0008936292, 0.0009330478, 
    0.0009994553, 0.0009796824, 0.001001584, 0.000991269, 0.0009844508, 
    0.001086287, 0.00117331, 0.001171053, 0.001177872, 0.001206403, 
    0.001241403, 0.001261795, 0.001253212, 0.001261716, 0.001067102, 
    0.001179636, 0.001190317, 0.001229481, 0.001259983, 0.001250828, 
    0.001168605, 0.001138835, 0.001118378, 0.001118442, 0.001160451, 
    0.001235283, 0.001289499, 0.001239606, 0.00125709, 0.001302056, 
    0.00130142, 0.001251114, 0.0009510096, 0.0008982231, 0.0009442382, 
    0.001057503, 0.00112658, 0.001115104, 0.00103835, 0.0009154365, 
    0.0006683241, 0.0006226911, 0.0005146242, 0.0003824923, 0.0004198276, 
    0.0005052448, 0.0005753404, 0.0006132964, 0.0005872138, 0.0005899156, 
    0.0006595021, 0.0007612277, 0.0008344692, 0.0008622529, 0.0008987784, 
    0.0009114631,
  0.0006850287, 0.0007760408, 0.0006963299, 0.0006688642, 0.0006893994, 
    0.0008195122, 0.0008384269, 0.0008519855, 0.0008246466, 0.0008131387, 
    0.000860441, 0.0009505791, 0.001035202, 0.001121843, 0.001208738, 
    0.001256994, 0.001245137, 0.001214921, 0.001184547, 0.00117455, 
    0.001139899, 0.00108136, 0.001053719, 0.001109143, 0.001155873, 
    0.001162851, 0.001087734, 0.001069932, 0.001077021, 0.001058377, 
    0.001005019, 0.0009545854, 0.0009002581, 0.0008639381, 0.0008289549, 
    0.0008312433, 0.0008169862, 0.0008228829, 0.0007440618, 0.0007362731, 
    0.0007522637, 0.0008275241, 0.0008549104, 0.0008296068, 0.0008184961, 
    0.0008584391, 0.0008395249, 0.0007840362, 0.0008601863, 0.0009814943, 
    0.001063129, 0.001081392, 0.0009472733, 0.0009066625, 0.0008644308, 
    0.0008293833, 0.0008331183, 0.0008588037, 0.0008721715, 0.0008845376, 
    0.0009153094, 0.0009665689, 0.001021914, 0.001072396, 0.001165331, 
    0.001270346, 0.001256391, 0.00115972, 0.001104057, 0.001084077, 
    0.001046614, 0.000836934, 0.000741503, 0.0006889391, 0.0007075993, 
    0.0007318386, 0.0008143478, 0.0007989777, 0.000655751, 0.0005621954, 
    0.0004954229, 0.0004309067, 0.0003337115, 0.0002580849, 0.0003032254, 
    0.0002617417, 0.0003833021, 0.0005332194, 0.0006518727, 0.0007426944, 
    0.0007520085, 0.0006926265, 0.0005981014, 0.0005391799, 0.000629541, 
    0.0006766361,
  0.0003993874, 0.0004024552, 0.0004424299, 0.0005412307, 0.0005782964, 
    0.0006087665, 0.0006027585, 0.0006327992, 0.0006843926, 0.000775055, 
    0.0008677999, 0.0009318707, 0.0009833854, 0.001051049, 0.001121795, 
    0.001165902, 0.001153538, 0.001116869, 0.001094633, 0.001101388, 
    0.001109748, 0.001079516, 0.001033693, 0.0009931936, 0.0009822736, 
    0.001036824, 0.001055643, 0.001046043, 0.001001713, 0.0009335249, 
    0.0008980641, 0.0008495222, 0.0007856579, 0.0007364326, 0.0007056922, 
    0.0007250835, 0.0007877238, 0.0008254736, 0.0007634845, 0.0007437437, 
    0.0007048494, 0.0007410732, 0.0007848309, 0.000801139, 0.0007519452, 
    0.0007215864, 0.0006694999, 0.0006463577, 0.0006897019, 0.0006861577, 
    0.0007562852, 0.0008427976, 0.0007893769, 0.0007834486, 0.0007643588, 
    0.0007517068, 0.0007605767, 0.000782765, 0.0007894726, 0.0008067656, 
    0.0008608871, 0.0009135297, 0.0009420915, 0.0009435061, 0.0009270874, 
    0.0009005754, 0.0008766062, 0.000861634, 0.0008604103, 0.0008670699, 
    0.0008447694, 0.0008004394, 0.000769302, 0.000739913, 0.0005829858, 
    0.000550529, 0.0005061356, 0.0005753245, 0.0005786943, 0.0005500047, 
    0.0004352296, 0.000386799, 0.0004020578, 0.0003205666, 0.0002870765, 
    0.0002654123, 0.000235403, 0.0002656826, 0.0003352845, 0.0004374073, 
    0.0004386944, 0.0004640147, 0.0003511156, 0.000240108, 0.0002527442, 
    0.0003022398,
  0.000448327, 0.0004140739, 0.0003848919, 0.0003532134, 0.0002919715, 
    0.0004649847, 0.0004945165, 0.0005419781, 0.0005970369, 0.0006552748, 
    0.0006841077, 0.0006830096, 0.0006928337, 0.0007243836, 0.0008624445, 
    0.0008937567, 0.0009068062, 0.0009123695, 0.0009064882, 0.0009004807, 
    0.0008967451, 0.0008686436, 0.0008368704, 0.000810819, 0.0008283979, 
    0.0009117967, 0.0009512948, 0.0008934864, 0.0008271264, 0.0007718133, 
    0.0007631509, 0.0007668065, 0.0007783461, 0.0007776944, 0.0007861026, 
    0.0007981346, 0.0007439184, 0.0007557916, 0.0007137982, 0.0006973473, 
    0.0006766208, 0.0006578334, 0.0006318775, 0.0006238029, 0.0006121206, 
    0.0005984032, 0.0005802517, 0.0005950336, 0.0006491069, 0.000710937, 
    0.0006950905, 0.0007039276, 0.0007107148, 0.0007491633, 0.0007638182, 
    0.0007908233, 0.0008333893, 0.0008469634, 0.0008829327, 0.0008302263, 
    0.0008165732, 0.0008070997, 0.000806432, 0.0008032054, 0.0007907278, 
    0.000777456, 0.0007668065, 0.0007553147, 0.0007276104, 0.0006281105, 
    0.0006321955, 0.0006565778, 0.000652604, 0.0004872528, 0.0005959398, 
    0.0005670118, 0.0006284441, 0.0006299382, 0.000649441, 0.0005082178, 
    0.000496265, 0.0004417624, 0.0004804337, 0.0003413092, 0.0002912889, 
    0.0002436687, 0.000224643, 0.0002333533, 0.0002750605, 0.0003408957, 
    0.0004074303, 0.0004424779, 0.0004095766, 0.0004263287, 0.0004558605, 
    0.000486108,
  0.000587245, 0.0005602245, 0.0005194074, 0.0004580542, 0.0003949846, 
    0.0004197326, 0.0005281973, 0.0006314004, 0.0006892886, 0.000700749, 
    0.0006793551, 0.0006590579, 0.0006431467, 0.0006351522, 0.0006035534, 
    0.0007721472, 0.0006862211, 0.0007096496, 0.0007131782, 0.0007743565, 
    0.0007271972, 0.0006871431, 0.0006691662, 0.0006582784, 0.0006764142, 
    0.00069091, 0.0007121135, 0.000724829, 0.0006926903, 0.0006702153, 
    0.0006923722, 0.0007206805, 0.0007359711, 0.0007357963, 0.0007133849, 
    0.0005642779, 0.0005426931, 0.000541501, 0.0006326246, 0.0006456738, 
    0.0006394589, 0.0006345317, 0.0006176995, 0.0006434962, 0.0006834075, 
    0.0007238113, 0.0007652487, 0.0008014245, 0.0008464858, 0.0008499825, 
    0.0008597258, 0.0008343423, 0.0007840996, 0.0007450308, 0.0007339839, 
    0.0007372424, 0.0007516749, 0.0007674263, 0.0007686976, 0.0007455235, 
    0.0007290249, 0.0007343816, 0.0007556644, 0.0008196242, 0.0008244561, 
    0.0008173669, 0.0007915699, 0.0007580484, 0.000702481, 0.0005537875, 
    0.0006232148, 0.0006426061, 0.000523397, 0.0007590181, 0.0008432274, 
    0.0008015202, 0.0007689204, 0.0007904891, 0.0006392049, 0.0005007314, 
    0.0004320983, 0.0004781135, 0.0003266068, 0.0002768884, 0.000249645, 
    0.0002388686, 0.0002296972, 0.000240601, 0.0002761571, 0.0003475241, 
    0.0005521984, 0.0005554087, 0.0005670593, 0.0005456975, 0.0005543279, 
    0.0005905838,
  0.0005452998, 0.000504896, 0.0005353182, 0.0005743713, 0.0005665985, 
    0.0005733701, 0.0006109132, 0.0006341189, 0.0006203223, 0.000605572, 
    0.0006116121, 0.0006335783, 0.0006629832, 0.0007019567, 0.000735224, 
    0.0007832574, 0.0008055891, 0.0008053347, 0.000785403, 0.0007519608, 
    0.0006893366, 0.0006225633, 0.0005616555, 0.0005105543, 0.0005042122, 
    0.0006123271, 0.0006495202, 0.0007041341, 0.0007368927, 0.0007764066, 
    0.0008045081, 0.0008319742, 0.0008342152, 0.0007923171, 0.0007727826, 
    0.0007599716, 0.0007427419, 0.0007483209, 0.000764597, 0.0007754213, 
    0.0007886617, 0.0007934142, 0.00079645, 0.0008049853, 0.0008208004, 
    0.0008428938, 0.0008723625, 0.000902149, 0.0009258478, 0.0009455569, 
    0.0009474166, 0.0009456207, 0.0009414243, 0.0009298371, 0.0009257364, 
    0.0009208885, 0.0009198237, 0.0009252914, 0.0009298848, 0.0009380706, 
    0.0009511042, 0.0009703684, 0.0009967053, 0.001026524, 0.001099782, 
    0.0009657906, 0.0009556659, 0.0009247191, 0.0008911975, 0.0008620149, 
    0.0008313863, 0.0008283027, 0.0008343108, 0.0008911815, 0.0009295354, 
    0.0009855158, 0.0009876456, 0.0008353437, 0.0005761037, 0.0005053094, 
    0.0004264088, 0.0003374945, 0.0002509325, 0.0001824906, 0.0001417527, 
    0.000127813, 0.0001427063, 0.000181934, 0.0002440342, 0.0003212343, 
    0.0004149011, 0.0006695797, 0.0008312906, 0.0007221268, 0.000621117, 
    0.0005677587,
  0.0008228028, 0.0008095468, 0.0007800306, 0.0007443633, 0.0006429721, 
    0.000650967, 0.0006684511, 0.0008421307, 0.0008530505, 0.0008584384, 
    0.0008740313, 0.0008819944, 0.0009030865, 0.0009058204, 0.0009026416, 
    0.0008887018, 0.0008458022, 0.0008047943, 0.0007722739, 0.0007399444, 
    0.0007139409, 0.00069207, 0.000669007, 0.0006490275, 0.0006360733, 
    0.000631353, 0.0006587235, 0.0007433463, 0.0007850059, 0.0008284139, 
    0.0008442131, 0.0008497604, 0.0008442927, 0.0008268561, 0.0008087046, 
    0.0007955121, 0.0007900603, 0.0007936208, 0.0008024423, 0.000814538, 
    0.0008281278, 0.0008391587, 0.000846645, 0.0008513815, 0.0008545287, 
    0.0008548307, 0.0008554187, 0.0008557687, 0.000856039, 0.0008568971, 
    0.0008586455, 0.0008587569, 0.0008539095, 0.0008438482, 0.0008345974, 
    0.0008243297, 0.0008151585, 0.0008096114, 0.0008073701, 0.0008098497, 
    0.0008182739, 0.0008318636, 0.0008504601, 0.0008711072, 0.0008877489, 
    0.0008949967, 0.0008940273, 0.0008935982, 0.0008887028, 0.0008741114, 
    0.0008556737, 0.0007973879, 0.0006557514, 0.0005658518, 0.0005146395, 
    0.0004708022, 0.0004312883, 0.0003931253, 0.0003538338, 0.0003117609, 
    0.0002685277, 0.0002267409, 0.0001908509, 0.0001647839, 0.0001548497, 
    0.0001610487, 0.0001859872, 0.0002308417, 0.000297901, 0.00038397, 
    0.0004844875, 0.0005838287, 0.000904581, 0.0009128142, 0.0008841399, 
    0.000857787,
  0.0008962203, 0.0008698034, 0.0008476622, 0.0008272696, 0.0008085617, 
    0.0007900286, 0.0007731804, 0.0007729259, 0.0007795222, 0.0007844813, 
    0.0007913319, 0.0007988977, 0.0008056051, 0.0008098013, 0.0008132823, 
    0.0008145698, 0.0008118679, 0.0008111526, 0.00080942, 0.0008071789, 
    0.0008048582, 0.0008068451, 0.0008097698, 0.0008114387, 0.0008144906, 
    0.0008232007, 0.0008230575, 0.0008272219, 0.0008303372, 0.0008252031, 
    0.0008105009, 0.0007913002, 0.0007717342, 0.000754409, 0.0007353673, 
    0.0007190439, 0.000706042, 0.0006949476, 0.0006867143, 0.0006834398, 
    0.0006841869, 0.0006870639, 0.0006907992, 0.000695202, 0.0007011307, 
    0.0007067574, 0.0007124636, 0.000720522, 0.0007275951, 0.0007335874, 
    0.0007355901, 0.0007349384, 0.0007345729, 0.0007309488, 0.0007285487, 
    0.0007258148, 0.0007267845, 0.0007311077, 0.0007378311, 0.0007488301, 
    0.0007623723, 0.0007782987, 0.0007976423, 0.0008202128, 0.000841257, 
    0.0008605055, 0.0008785616, 0.0008955686, 0.0009089997, 0.0009208095, 
    0.0009281208, 0.0009336045, 0.0009402484, 0.0009400417, 0.0009418061, 
    0.0009430777, 0.0009408365, 0.0009365927, 0.0009332548, 0.0009288202, 
    0.0009224465, 0.000912433, 0.0009049466, 0.0009025942, 0.0009082686, 
    0.0009192675, 0.0009438246, 0.0009691606, 0.000990666, 0.0009922237, 
    0.0009940516, 0.0009888064, 0.000984372, 0.0009741678, 0.0009481162, 
    0.0009251327,
  0.0008092931, 0.0007933987, 0.000784132, 0.0007758035, 0.0007686826, 
    0.0007628174, 0.0007567616, 0.0007517707, 0.0007493231, 0.0007491164, 
    0.0007477972, 0.0007487984, 0.0007502449, 0.0007535351, 0.0007554266, 
    0.000758621, 0.0007642478, 0.0007693182, 0.0007734825, 0.0007763753, 
    0.0007778854, 0.0007781873, 0.0007793, 0.0007780284, 0.0007748336, 
    0.0007707486, 0.0007659488, 0.0007602904, 0.0007537734, 0.0007453969, 
    0.0007360668, 0.0007261966, 0.0007119867, 0.0007003041, 0.0006897022, 
    0.0006780833, 0.0006676406, 0.0006572616, 0.00064604, 0.0006365827, 
    0.0006290327, 0.0006206563, 0.0006149502, 0.0006097686, 0.0006066054, 
    0.0006046824, 0.000602012, 0.0005991034, 0.000599453, 0.0006022505, 
    0.0006067645, 0.000611501, 0.0006170642, 0.0006241532, 0.000632307, 
    0.0006428611, 0.0006550681, 0.0006655426, 0.000679482, 0.0006930243, 
    0.0007062007, 0.0007225563, 0.0007383872, 0.0007554581, 0.0007726083, 
    0.0007907758, 0.0008095632, 0.0008278895, 0.0008451034, 0.0008613159, 
    0.0008773694, 0.0008905936, 0.0009032458, 0.0009165815, 0.0009297421, 
    0.0009397875, 0.0009486248, 0.000955046, 0.0009580184, 0.0009592264, 
    0.0009601483, 0.0009587494, 0.0009559839, 0.0009516765, 0.0009466221, 
    0.0009441266, 0.0009401372, 0.0009341926, 0.0009271038, 0.0009171059, 
    0.0009054235, 0.0008919131, 0.0008781803, 0.0008629693, 0.0008445634, 
    0.0008268885,
  1.629082e-005, 1.554377e-005, 1.490798e-005, 1.411326e-005, 1.347749e-005, 
    1.284169e-005, 1.217413e-005, 1.160192e-005, 1.099793e-005, 
    1.040984e-005, 9.917097e-006, 9.456158e-006, 9.090585e-006, 
    8.740899e-006, 8.470692e-006, 8.184594e-006, 8.07333e-006, 7.803123e-006, 
    7.691862e-006, 7.628281e-006, 7.501127e-006, 7.564704e-006, 
    7.612391e-006, 7.580598e-006, 7.644179e-006, 7.803123e-006, 
    7.962066e-006, 8.200484e-006, 8.518378e-006, 8.772691e-006, 
    9.011106e-006, 9.185947e-006, 9.567415e-006, 9.901203e-006, 
    1.036215e-005, 1.082309e-005, 1.126813e-005, 1.172908e-005, 1.22536e-005, 
    1.28258e-005, 1.339801e-005, 1.39702e-005, 1.457419e-005, 1.520997e-005, 
    1.584576e-005, 1.633849e-005, 1.695837e-005, 1.7467e-005, 1.802331e-005, 
    1.850015e-005, 1.905646e-005, 1.929488e-005, 1.959688e-005, 
    1.986708e-005, 2.01214e-005, 2.043929e-005, 2.072538e-005, 2.109096e-005, 
    2.093201e-005, 2.137706e-005, 2.18698e-005, 2.210822e-005, 2.2442e-005, 
    2.266453e-005, 2.280757e-005, 2.295063e-005, 2.291884e-005, 
    2.288706e-005, 2.279169e-005, 2.283938e-005, 2.291884e-005, 
    2.290294e-005, 2.293474e-005, 2.261684e-005, 2.299831e-005, 2.30301e-005, 
    2.3046e-005, 2.272811e-005, 2.307779e-005, 2.306189e-005, 2.306189e-005, 
    2.309368e-005, 2.299831e-005, 2.285525e-005, 2.266452e-005, 
    2.239432e-005, 2.21559e-005, 2.167906e-005, 2.121812e-005, 2.078897e-005, 
    2.026444e-005, 1.967636e-005, 1.907235e-005, 1.842068e-005, 
    1.772132e-005, 1.699016e-005,
  1.830942e-005, 1.60365e-005, 1.425631e-005, 1.287347e-005, 1.179266e-005, 
    1.088666e-005, 1.017141e-005, 9.599207e-006, 9.154159e-006, 
    8.820378e-006, 8.407114e-006, 8.025647e-006, 7.580602e-006, 7.13555e-006, 
    6.769973e-006, 6.452083e-006, 6.150087e-006, 5.863985e-006, 
    5.689144e-006, 5.530195e-006, 5.546091e-006, 5.657352e-006, 
    6.054717e-006, 6.372606e-006, 6.595132e-006, 6.897129e-006, 
    7.167338e-006, 7.45344e-006, 7.834911e-006, 8.39122e-006, 9.058793e-006, 
    9.774049e-006, 1.07913e-005, 1.203108e-005, 1.371591e-005, 1.595703e-005, 
    1.862731e-005, 2.179032e-005, 2.53825e-005, 2.932436e-005, 3.325031e-005, 
    3.727165e-005, 4.070488e-005, 4.437653e-005, 4.690376e-005, 
    4.780975e-005, 5.076613e-005, 5.200591e-005, 5.299138e-005, 
    5.318211e-005, 5.389737e-005, 5.553453e-005, 5.53279e-005, 5.747365e-005, 
    5.458084e-005, 6.057313e-005, 6.043007e-005, 5.992145e-005, 
    6.019167e-005, 5.977838e-005, 5.926975e-005, 5.869754e-005, 5.70604e-005, 
    5.502588e-005, 5.30073e-005, 5.087742e-005, 4.849321e-005, 4.588649e-005, 
    4.342284e-005, 4.119761e-005, 3.960815e-005, 3.811406e-005, 
    3.668355e-005, 3.580934e-005, 3.585701e-005, 3.631799e-005, 
    3.661997e-005, 3.720805e-005, 3.65087e-005, 3.782795e-005, 3.79074e-005, 
    3.633385e-005, 3.811403e-005, 3.6461e-005, 3.774845e-005, 3.789153e-005, 
    3.890878e-005, 3.906772e-005, 3.870216e-005, 3.762131e-005, 
    3.577756e-005, 3.315497e-005, 3.018267e-005, 2.694016e-005, 
    2.380893e-005, 2.090022e-005,
  1.125223e-005, 8.391216e-006, 6.769973e-006, 6.070615e-006, 5.927563e-006, 
    6.181876e-006, 6.309034e-006, 6.51566e-006, 6.769973e-006, 7.04018e-006, 
    7.564704e-006, 8.025647e-006, 8.534273e-006, 9.090581e-006, 
    9.646898e-006, 1.033036e-005, 1.091845e-005, 1.134761e-005, 
    1.134761e-005, 1.091845e-005, 1.025089e-005, 9.265423e-006, 
    8.454801e-006, 7.834911e-006, 7.246814e-006, 6.960709e-006, 
    6.992495e-006, 7.405757e-006, 8.105115e-006, 8.899849e-006, 
    9.774049e-006, 1.061646e-005, 1.13794e-005, 1.246023e-005, 1.392253e-005, 
    1.586167e-005, 1.888163e-005, 2.269632e-005, 2.792563e-005, 
    3.398147e-005, 4.060951e-005, 4.672892e-005, 5.20059e-005, 5.528018e-005, 
    5.601133e-005, 5.7871e-005, 5.926973e-005, 6.141551e-005, 6.370433e-005, 
    6.592958e-005, 6.879057e-005, 7.249402e-005, 7.742137e-005, 
    8.242816e-005, 8.668788e-005, 8.97237e-005, 9.126548e-005, 9.008928e-005, 
    8.695805e-005, 8.315925e-005, 7.951941e-005, 7.673787e-005, 
    7.430598e-005, 7.155628e-005, 6.867935e-005, 6.61839e-005, 6.327516e-005, 
    6.043006e-005, 5.793461e-005, 5.524841e-005, 5.159267e-005, 
    4.811175e-005, 4.59501e-005, 4.5362e-005, 4.502821e-005, 4.572755e-005, 
    4.633155e-005, 4.925614e-005, 5.229199e-005, 5.491459e-005, 
    5.755312e-005, 6.14473e-005, 6.538912e-005, 6.887008e-005, 6.92833e-005, 
    6.850448e-005, 6.834551e-005, 6.847267e-005, 6.635868e-005, 
    6.116118e-005, 5.590005e-005, 4.742826e-005, 3.863855e-005, 
    2.981711e-005, 2.18857e-005, 1.562323e-005,
  2.102739e-005, 1.86273e-005, 1.754649e-005, 1.708555e-005, 1.671997e-005, 
    1.656104e-005, 1.648156e-005, 1.60683e-005, 1.51782e-005, 1.42881e-005, 
    1.347748e-005, 1.306422e-005, 1.325496e-005, 1.441526e-005, 
    1.671998e-005, 2.001014e-005, 2.436525e-005, 2.827531e-005, 
    3.091381e-005, 3.100916e-005, 2.838656e-005, 2.382482e-005, 
    1.912004e-005, 1.51464e-005, 1.268276e-005, 1.155424e-005, 1.153834e-005, 
    1.244434e-005, 1.397021e-005, 1.559146e-005, 1.702197e-005, 
    1.822996e-005, 1.937437e-005, 1.98353e-005, 1.975583e-005, 1.966046e-005, 
    2.01373e-005, 2.161549e-005, 2.446062e-005, 2.921309e-005, 3.539609e-005, 
    4.21195e-005, 4.947867e-005, 5.628157e-005, 6.222611e-005, 6.798e-005, 
    9.120192e-005, 9.186947e-005, 9.589081e-005, 9.887901e-005, 0.0001004366, 
    0.0001031387, 0.000106874, 0.000112898, 0.0001232137, 0.0001366445, 
    0.0001577843, 0.0001198122, 0.000113645, 0.0001057931, 9.8577e-005, 
    9.714649e-005, 9.738488e-005, 9.662195e-005, 9.732132e-005, 
    9.760741e-005, 9.668554e-005, 9.566828e-005, 9.261654e-005, 
    9.129726e-005, 9.368142e-005, 9.660603e-005, 9.916507e-005, 0.0001000869, 
    9.922867e-005, 9.662195e-005, 9.506429e-005, 9.533454e-005, 
    9.452386e-005, 9.248935e-005, 0.0001118808, 0.0001063336, 0.0001079549, 
    0.0001100052, 0.000117126, 0.0001227208, 0.0001247713, 0.0001241037, 
    0.0001257886, 9.584322e-005, 8.330229e-005, 7.061844e-005, 5.54391e-005, 
    4.261221e-005, 3.274171e-005, 2.549377e-005,
  4.38838e-005, 4.067307e-005, 3.854319e-005, 3.687428e-005, 3.555504e-005, 
    3.483974e-005, 3.553914e-005, 3.773256e-005, 4.229434e-005, 
    4.552095e-005, 4.506001e-005, 4.053005e-005, 3.371124e-005, 
    2.717859e-005, 2.357052e-005, 2.396788e-005, 2.80051e-005, 3.439472e-005, 
    4.21513e-005, 4.666534e-005, 5.003499e-005, 4.842963e-005, 4.191288e-005, 
    3.466495e-005, 2.989655e-005, 2.792563e-005, 2.775079e-005, 
    2.867267e-005, 3.007139e-005, 3.158138e-005, 3.275758e-005, 
    3.339336e-005, 3.44265e-005, 3.603187e-005, 3.809814e-005, 4.005319e-005, 
    4.110223e-005, 4.105455e-005, 4.135654e-005, 4.316853e-005, 
    4.548916e-005, 4.82707e-005, 5.102044e-005, 5.448544e-005, 5.828428e-005, 
    6.470563e-005, 7.872464e-005, 9.52392e-005, 0.0001092741, 0.0001162518, 
    0.0001143445, 0.0001025983, 9.21397e-005, 9.34907e-005, 0.0001088131, 
    0.0001348007, 0.0001617896, 0.000175761, 0.0001761901, 0.0001675117, 
    0.000157228, 0.0001518714, 0.0001601843, 0.0001763967, 0.0001964875, 
    0.0002127953, 0.0002254474, 0.0002397844, 0.0002567439, 0.0002750703, 
    0.0002586829, 0.0002842733, 0.0002875793, 0.0002840984, 0.0002784717, 
    0.0002656924, 0.0002352544, 0.0002144961, 0.0001970757, 0.000184662, 
    0.0001968372, 0.0001841533, 0.0001805452, 0.000178765, 0.0001848209, 
    0.0001934834, 0.000201987, 0.0002066123, 0.0002023049, 0.0001840738, 
    0.0001617101, 0.0001058567, 8.053673e-005, 6.314804e-005, 5.310262e-005, 
    4.855674e-005,
  0.0001898594, 0.0001766669, 0.0001293648, 0.0001104343, 9.611339e-005, 
    8.942166e-005, 9.029586e-005, 9.733721e-005, 0.0001072237, 0.0001177935, 
    0.0001203843, 0.0001131683, 9.794123e-005, 7.818424e-005, 6.146322e-005, 
    5.068666e-005, 4.782564e-005, 5.179932e-005, 6.311623e-005, 
    7.359067e-005, 8.247577e-005, 8.274597e-005, 7.699215e-005, 
    6.982373e-005, 6.564346e-005, 6.400634e-005, 6.664483e-005, 
    7.206475e-005, 7.842269e-005, 8.280959e-005, 8.406522e-005, 
    8.133138e-005, 7.711933e-005, 7.398811e-005, 7.209665e-005, 
    7.436957e-005, 7.664249e-005, 7.866111e-005, 7.769151e-005, 
    7.371785e-005, 6.966476e-005, 6.793224e-005, 6.920382e-005, 
    7.241455e-005, 8.600444e-005, 9.201257e-005, 9.544578e-005, 0.0001037426, 
    0.000107144, 0.0001059201, 9.660586e-005, 8.649682e-005, 7.735763e-005, 
    7.382897e-005, 8.323847e-005, 0.0001079069, 0.0001414445, 0.0001740283, 
    0.0002018438, 0.0002170232, 0.0002269573, 0.0002409921, 0.0002552972, 
    0.0002712554, 0.0002880718, 0.0003038555, 0.0003272999, 0.0003562439, 
    0.0003872383, 0.0004128604, 0.0004307894, 0.0004522948, 0.0004739433, 
    0.0004819541, 0.0004742771, 0.0004529465, 0.000425433, 0.0003976173, 
    0.0003522385, 0.0003351042, 0.000359232, 0.0003417957, 0.0003257898, 
    0.0003029017, 0.0002821431, 0.0002727176, 0.0002749428, 0.0002745454, 
    0.000269777, 0.0002658035, 0.0002637375, 0.0002588101, 0.0002486376, 
    0.0002333469, 0.0002203929, 0.000207264,
  0.000304618, 0.0002926018, 0.000278726, 0.0002593029, 0.0002569822, 
    0.0002619731, 0.0002698251, 0.0002735762, 0.0002744821, 0.0002747683, 
    0.0002766121, 0.0002719073, 0.0002687919, 0.0002649295, 0.0002514826, 
    0.0002356835, 0.0002162126, 0.0002122071, 0.0002228725, 0.0002363987, 
    0.0002403723, 0.0002342371, 0.0002195504, 0.0002019393, 0.0001869348, 
    0.0001797187, 0.0001793531, 0.0001742668, 0.0001624255, 0.0001472142, 
    0.0001426205, 0.000152364, 0.000166828, 0.0001947072, 0.0002024479, 
    0.0002112694, 0.0002337284, 0.0002421206, 0.0002442823, 0.0002422796, 
    0.0002407538, 0.0002331086, 0.0002222209, 0.0002042757, 0.0001809743, 
    0.0001633313, 0.0001535562, 0.0001440354, 0.0001027415, 5.262578e-005, 
    6.309245e-006, -1.204922e-005, -6.708549e-006, -3.879191e-006, 
    3.538025e-005, 6.753509e-005, 0.0001003257, 0.0001324962, 0.0001645397, 
    0.0001943737, 0.0002322505, 0.0002706675, 0.0003043481, 0.0003344365, 
    0.0003613617, 0.000379863, 0.0004077265, 0.0004486551, 0.0004787913, 
    0.0005364566, 0.000568818, 0.0006290583, 0.0006668876, 0.0006922234, 
    0.0006790627, 0.000663057, 0.0006386586, 0.0006097306, 0.0005717744, 
    0.0005303371, 0.0005004237, 0.0004956552, 0.0004930008, 0.0004832257, 
    0.0004728623, 0.0004637548, 0.0004483371, 0.0004248926, 0.0003913391, 
    0.0003678151, 0.0003621246, 0.0003589778, 0.0003461507, 0.0003289049, 
    0.0003177311, 0.0003131535,
  0.0004296132, 0.0004143227, 0.0003905445, 0.0003776539, 0.000385045, 
    0.0003969499, 0.000396346, 0.0003882556, 0.0003841706, 0.0003966956, 
    0.0004094908, 0.0004225562, 0.0004414389, 0.0004441724, 0.0004532803, 
    0.0004257986, 0.0004158008, 0.0004283894, 0.0004295338, 0.0004428852, 
    0.0004419793, 0.0004303921, 0.0004083781, 0.0003635078, 0.0003037439, 
    0.0002474295, 0.0002081542, 0.0001791941, 0.0001483907, 0.0001166809, 
    8.493965e-005, 7.149298e-005, 0.0001322259, 0.000171867, 0.0002154661, 
    0.0003044757, 0.000362427, 0.0003598365, 0.0003420981, 0.000323819, 
    0.000298626, 0.0002848455, 0.0002724794, 0.0002684421, 0.0002758333, 
    0.000271383, 0.0002596527, 0.0002082651, 6.616767e-005, -7.16697e-005, 
    -0.0001561334, -0.0001745392, -0.0001538289, -0.0001089904, 
    -4.987838e-005, -1.298706e-005, -7.789349e-006, -3.481982e-006, 
    3.801892e-005, 0.0001030595, 0.0001633794, 0.000228531, 0.0002754994, 
    0.0003237394, 0.0003839959, 0.0004533122, 0.0005025694, 0.0005812, 
    0.0006729274, 0.0007597278, 0.0008097319, 0.0008305062, 0.0008522184, 
    0.0008614529, 0.000878365, 0.0008764097, 0.0008504221, 0.0007587583, 
    0.0006527414, 0.0005492517, 0.000491634, 0.0005206892, 0.0005566746, 
    0.0005630646, 0.0005373468, 0.0005231372, 0.0005143951, 0.0005012979, 
    0.0004779327, 0.0004725443, 0.0004877239, 0.0005001534, 0.0004872152, 
    0.0004559348, 0.0004364798, 0.000433889,
  0.0004918086, 0.0004858801, 0.0004743407, 0.000469334, 0.000487247, 
    0.0004830193, 0.0004636913, 0.0004530577, 0.0004420909, 0.0004439666, 
    0.0004276426, 0.0004369887, 0.0004517864, 0.0004521839, 0.0004953535, 
    0.0005629053, 0.0006007503, 0.0006119718, 0.0006265475, 0.0006666973, 
    0.0006714335, 0.0006498965, 0.0006104778, 0.0005514135, 0.0004517387, 
    0.0003536851, 0.0002898842, 0.0002298346, 0.0002073916, 0.0001917987, 
    0.000190543, 0.0001804659, 0.0001743785, 0.0001448623, 0.0001369941, 
    0.0001773499, 0.0002828899, 0.0003508874, 0.0003556404, 0.0003487421, 
    0.0004024652, 0.0004847511, 0.0005803092, 0.0006395478, 0.0006288358, 
    0.0005969196, 0.0005129487, 0.0003840907, 0.0001970916, -2.225349e-005, 
    -9.040954e-005, -7.874309e-005, -7.966487e-005, -0.0001178277, 
    -0.0001947414, -0.0002344302, -0.000252407, -0.0002355271, -0.0001194177, 
    3.067474e-005, 0.0001565602, 0.0002525954, 0.0003178264, 0.0004021314, 
    0.0004853872, 0.0005683887, 0.0006393576, 0.0006925727, 0.0007416389, 
    0.0007944726, 0.0008327309, 0.0008422835, 0.0008594657, 0.0008729766, 
    0.0008625663, 0.0008049323, 0.0007210411, 0.0006929236, 0.0006710207, 
    0.0006373082, 0.0005965855, 0.0005379505, 0.0004150702, 0.0003379812, 
    0.0003255834, 0.0003465482, 0.0004097291, 0.0004784416, 0.0005134414, 
    0.0005237572, 0.0005260461, 0.0005347081, 0.0005513977, 0.0005464226, 
    0.0005250762, 0.0005009801,
  0.0003676882, 0.0004109533, 0.0004863252, 0.0005312115, 0.0005221039, 
    0.0005213569, 0.0005413361, 0.0005880026, 0.0006202529, 0.0006105255, 
    0.0005831867, 0.0005691675, 0.000580119, 0.0005987475, 0.0006298216, 
    0.0006689539, 0.0007171622, 0.0007582179, 0.0007435631, 0.000608936, 
    0.0005029829, 0.0004529308, 0.0004244477, 0.0004538684, 0.0004506577, 
    0.0004369728, 0.0004649314, 0.0004876601, 0.0004969744, 0.0005050004, 
    0.000488979, 0.0004327442, 0.0003715027, 0.000344832, 0.0003610607, 
    0.0003951546, 0.0004565869, 0.0005305288, 0.0005781963, 0.0005748109, 
    0.0006050579, 0.0006824648, 0.0007575187, 0.0007450571, 0.0006832751, 
    0.0006820988, 0.0006789356, 0.0006415993, 0.0005158731, 0.0003301292, 
    0.0002434882, 0.0002102363, 0.0001857588, 0.0001289831, 5.213358e-005, 
    1.921551e-005, 2.763979e-005, 5.253032e-005, 0.000110514, 0.0001862831, 
    0.0002580476, 0.0002985308, 0.0003379015, 0.0003879224, 0.0004340159, 
    0.0004846877, 0.0005412092, 0.0005935188, 0.0006377529, 0.0006784904, 
    0.0007191175, 0.0007431661, 0.0007586153, 0.000745296, 0.000692843, 
    0.0006191563, 0.0006579072, 0.0008592596, 0.0008937195, 0.0006678565, 
    0.0006325869, 0.0005821227, 0.000527651, 0.0003812772, 0.0002911242, 
    0.0003278248, 0.0003920549, 0.0004081875, 0.0004306147, 0.0004405805, 
    0.0004363209, 0.0004396269, 0.0004313935, 0.0004244635, 0.0004091254, 
    0.0003766844,
  0.0006065194, 0.0006313622, 0.0006673317, 0.0006794918, 0.0006822259, 
    0.0006878048, 0.0007122504, 0.0007315304, 0.000750286, 0.0007827266, 
    0.0008034848, 0.000822813, 0.0008400106, 0.0008442863, 0.0008365775, 
    0.000835561, 0.0008819725, 0.0009617477, 0.0009875444, 0.0009109175, 
    0.0008188719, 0.0008188076, 0.000827756, 0.0008215262, 0.0007967311, 
    0.0007925346, 0.0008055842, 0.000820525, 0.0008371505, 0.0008468935, 
    0.0008126083, 0.0007287175, 0.0006387546, 0.0005996693, 0.0006003529, 
    0.0006060908, 0.0006174557, 0.0006230664, 0.0006151348, 0.00064357, 
    0.000733613, 0.0008216687, 0.0008478472, 0.0008292347, 0.0008828803, 
    0.0009209784, 0.0008913665, 0.0007931064, 0.0007101689, 0.0006250055, 
    0.0005347719, 0.0004628967, 0.0004296131, 0.0004011621, 0.0003474383, 
    0.0003104517, 0.0003202748, 0.0003447682, 0.0003770501, 0.0004258305, 
    0.0004391978, 0.0004332694, 0.0004590186, 0.0004791091, 0.0004741498, 
    0.0004985165, 0.0005369494, 0.0005562296, 0.0005753026, 0.0005946308, 
    0.0006036749, 0.0006134021, 0.0005952031, 0.0005665449, 0.0005309097, 
    0.000573046, 0.0006834972, 0.0007630652, 0.0007008864, 0.0006367038, 
    0.0005836952, 0.0005554184, 0.0005448963, 0.0004789499, 0.0004451899, 
    0.0004943362, 0.0005656392, 0.0006253705, 0.0006547596, 0.0006771549, 
    0.0006745965, 0.0006607999, 0.0006370216, 0.0006048027, 0.0005919922, 
    0.0005884792,
  0.0007262062, 0.0007750983, 0.0008148025, 0.0008587027, 0.0008895062, 
    0.0009336299, 0.001011625, 0.001086997, 0.001124174, 0.00114204, 
    0.001181157, 0.00121506, 0.001210594, 0.001165533, 0.001104784, 
    0.001054334, 0.001053921, 0.001094515, 0.001124843, 0.001220973, 
    0.00143787, 0.00159691, 0.001571766, 0.001426235, 0.001326544, 
    0.001257609, 0.001169331, 0.001091225, 0.00103712, 0.0009782938, 
    0.0008897781, 0.0007988294, 0.0007503671, 0.000728528, 0.0007132371, 
    0.0007020789, 0.0006746291, 0.0006325403, 0.0006114482, 0.0006783647, 
    0.0008509164, 0.0009728917, 0.001010625, 0.0009910273, 0.001098108, 
    0.001079703, 0.001028824, 0.0009857179, 0.0009367941, 0.0008911765, 
    0.0008272328, 0.0007833955, 0.0007564705, 0.0007150653, 0.0006472589, 
    0.000614468, 0.0006425856, 0.0006411234, 0.0006057424, 0.0005955854, 
    0.0005901973, 0.00055933, 0.0005666255, 0.0005471073, 0.0005356153, 
    0.0005619209, 0.0005509853, 0.0005338667, 0.0005549113, 0.0005386039, 
    0.0005124728, 0.0005246797, 0.000550922, 0.0005560238, 0.0005419571, 
    0.0005373321, 0.0005902443, 0.000670623, 0.0006393902, 0.0006162315, 
    0.0005699145, 0.0005536862, 0.0005917381, 0.000601545, 0.0005553076, 
    0.000535646, 0.0005589956, 0.0006107315, 0.0006598942, 0.0006910632, 
    0.0006935904, 0.0006977073, 0.0007023169, 0.000678062, 0.0006605936, 
    0.0006816066,
  0.0009598099, 0.00100414, 0.001034784, 0.001052984, 0.00108916, 
    0.001221069, 0.001468405, 0.001678166, 0.001795261, 0.001884222, 
    0.001965126, 0.001980703, 0.001841752, 0.001679882, 0.001606672, 
    0.001541329, 0.001514038, 0.001502371, 0.001542219, 0.001646901, 
    0.001700258, 0.001653703, 0.001513228, 0.001326021, 0.001227475, 
    0.001168649, 0.001086951, 0.001022292, 0.0009492082, 0.000867717, 
    0.0008118795, 0.0008001332, 0.0007860027, 0.0007400997, 0.0006564301, 
    0.0006071571, 0.0006264853, 0.0006745649, 0.0007686927, 0.0008345284, 
    0.000977166, 0.001110284, 0.001191156, 0.001221959, 0.001309602, 
    0.001410882, 0.001317311, 0.001249504, 0.001284933, 0.001313909, 
    0.001316388, 0.001269197, 0.00117483, 0.001046911, 0.0009475066, 
    0.0008749957, 0.000833733, 0.0007768464, 0.0006960556, 0.0006789532, 
    0.000669146, 0.0006546662, 0.00065473, 0.0006206995, 0.0006236238, 
    0.0006253566, 0.0005962057, 0.0005931226, 0.0006095096, 0.0006110831, 
    0.0006369278, 0.0006637736, 0.0006609447, 0.0006258176, 0.0005571051, 
    0.0004972145, 0.000538588, 0.0006255778, 0.0005510794, 0.0006822911, 
    0.0006459397, 0.0006023725, 0.0006178059, 0.0006869952, 0.0006811302, 
    0.0006440324, 0.0006680647, 0.0007140636, 0.0007677241, 0.0008166786, 
    0.0008039, 0.000792122, 0.0008035344, 0.0008081277, 0.0008711657, 
    0.0009394647,
  0.001052729, 0.001034116, 0.0009876718, 0.0009920909, 0.001141501, 
    0.001406781, 0.001617143, 0.001789059, 0.002031771, 0.00213456, 
    0.001970067, 0.001758033, 0.001566855, 0.001436376, 0.001387835, 
    0.001329073, 0.001307694, 0.001281865, 0.001250742, 0.001248708, 
    0.00117041, 0.001091415, 0.00102957, 0.0009409906, 0.0008826256, 
    0.0008397251, 0.000819461, 0.0008213036, 0.0008395985, 0.0009486512, 
    0.001054573, 0.001030094, 0.000934632, 0.0007697269, 0.000669335, 
    0.0007020943, 0.0008135, 0.0008615339, 0.00092756, 0.001113287, 
    0.001251314, 0.001469769, 0.001545379, 0.001495391, 0.001492959, 
    0.001496917, 0.001484741, 0.001390328, 0.001431686, 0.001342423, 
    0.001166373, 0.001119978, 0.001097121, 0.0009815348, 0.0009368714, 
    0.0008957386, 0.000830777, 0.0007880675, 0.0007388275, 0.0007263031, 
    0.0007192767, 0.0007250467, 0.0007389854, 0.0007504462, 0.0007849373, 
    0.0007785796, 0.0007514786, 0.0007732711, 0.0008025803, 0.0007968261, 
    0.0008151368, 0.0007809158, 0.000720453, 0.0006877738, 0.0006049471, 
    0.0005628583, 0.0005978579, 0.0007043839, 0.0007599196, 0.0007893411, 
    0.0007084692, 0.0007390664, 0.0008723736, 0.0009365389, 0.0009344104, 
    0.0009247465, 0.0009688525, 0.0009803451, 0.000969267, 0.0009720312, 
    0.0009620502, 0.000988483, 0.001049391, 0.001063474, 0.001092529, 
    0.001090828,
  0.0009730645, 0.0009545777, 0.0009245854, 0.001039996, 0.001256098, 
    0.001412153, 0.001594685, 0.001729979, 0.002053227, 0.001988078, 
    0.001504961, 0.001330503, 0.001361416, 0.001339846, 0.001297409, 
    0.001190597, 0.001143612, 0.001113619, 0.001008591, 0.0009076437, 
    0.0008216696, 0.0007888945, 0.0007987954, 0.0007975558, 0.000805567, 
    0.0008262768, 0.0008820677, 0.0009699967, 0.001082516, 0.001274966, 
    0.001166773, 0.001129866, 0.001136461, 0.001057021, 0.001007191, 
    0.001026853, 0.001000179, 0.00126233, 0.001317216, 0.001430067, 
    0.001549751, 0.001879515, 0.001910112, 0.001755714, 0.001658932, 
    0.001613123, 0.001574405, 0.001477369, 0.001331918, 0.00108633, 
    0.0008778414, 0.0008828323, 0.0009447252, 0.0009257793, 0.0009196419, 
    0.0009110905, 0.0009044791, 0.0009031594, 0.0008622939, 0.0008432688, 
    0.0008707503, 0.0008877581, 0.0009034611, 0.0009691054, 0.001019587, 
    0.001014294, 0.001008684, 0.0009936467, 0.0009461064, 0.0009195777, 
    0.0008994248, 0.0007997816, 0.0007372517, 0.0007228833, 0.000638024, 
    0.0006601643, 0.0006975643, 0.001086569, 0.0009737019, 0.0009173383, 
    0.0008010054, 0.0009488566, 0.001269102, 0.00153551, 0.001413614, 
    0.001288618, 0.001278923, 0.001274027, 0.001237486, 0.001189216, 
    0.001119502, 0.001114703, 0.001132536, 0.001110681, 0.001069877, 
    0.001010798,
  0.001025645, 0.0009812834, 0.0009364597, 0.001068641, 0.001175738, 
    0.001143997, 0.001207702, 0.001698508, 0.002192592, 0.002109922, 
    0.001912736, 0.001954254, 0.001986456, 0.001878547, 0.001730188, 
    0.001620324, 0.001519918, 0.00143431, 0.001329261, 0.001302383, 
    0.001360478, 0.001357665, 0.001344361, 0.001326784, 0.00128975, 
    0.001258183, 0.001318248, 0.001415174, 0.001431307, 0.001367392, 
    0.0012643, 0.001695506, 0.001285013, 0.001240556, 0.001205476, 
    0.001241176, 0.001407622, 0.001534447, 0.001607785, 0.001583686, 
    0.001390839, 0.001493677, 0.001319345, 0.001398514, 0.001533554, 
    0.001586404, 0.001523906, 0.001330787, 0.001161272, 0.001071991, 
    0.001044351, 0.001067318, 0.001117053, 0.001126414, 0.001092876, 
    0.001086169, 0.001062171, 0.001004647, 0.0009279726, 0.0009252867, 
    0.0009456156, 0.0009904699, 0.001022686, 0.001096136, 0.001096437, 
    0.001072293, 0.001088745, 0.001023466, 0.0009811381, 0.0009759245, 
    0.0008958494, 0.0008888403, 0.0008234978, 0.0007196749, 0.0007175421, 
    0.0007741749, 0.0008198721, 0.001012388, 0.001321125, 0.001355172, 
    0.001269561, 0.001550068, 0.001626076, 0.001779302, 0.001757178, 
    0.001606193, 0.001531808, 0.001447996, 0.001450252, 0.001395448, 
    0.001285951, 0.001204696, 0.001161908, 0.001138844, 0.001061978, 
    0.001011022,
  0.001043143, 0.0010296, 0.001084438, 0.001228585, 0.001377231, 0.001332602, 
    0.001670184, 0.002167987, 0.002292856, 0.002264212, 0.002449446, 
    0.002523722, 0.002498832, 0.002324977, 0.002175122, 0.002076244, 
    0.002018499, 0.001888117, 0.00185628, 0.001888736, 0.001912531, 
    0.001862685, 0.001765219, 0.001724892, 0.001644816, 0.001572686, 
    0.001543918, 0.0015213, 0.001481054, 0.001582574, 0.001590967, 
    0.002025602, 0.00177423, 0.001125923, 0.0009136342, 0.001098489, 
    0.001203315, 0.001332283, 0.001663127, 0.001744842, 0.001476476, 
    0.001261012, 0.001126687, 0.001270882, 0.001392699, 0.001493135, 
    0.001519664, 0.001596069, 0.001585308, 0.00149533, 0.001476192, 
    0.001450825, 0.001389774, 0.001289765, 0.00116647, 0.001079671, 
    0.001015234, 0.0009222664, 0.0009264313, 0.0009921705, 0.001021576, 
    0.001073185, 0.001069784, 0.001122857, 0.001192966, 0.001169221, 
    0.001157268, 0.001131153, 0.001119249, 0.001093102, 0.001002708, 
    0.0009869263, 0.0008510724, 0.0008313339, 0.0007918831, 0.000810083, 
    0.001122838, 0.0008711806, 0.001704376, 0.001843276, 0.001812616, 
    0.002191273, 0.002320528, 0.002317492, 0.002258792, 0.002108954, 
    0.001982035, 0.001836425, 0.001731793, 0.001550913, 0.001461585, 
    0.001422072, 0.001388979, 0.001301797, 0.001176929, 0.001058036,
  0.001245595, 0.001286347, 0.001407639, 0.001689211, 0.001326688, 
    0.001538817, 0.002302933, 0.002766815, 0.002802465, 0.002655631, 
    0.002849068, 0.002800781, 0.003035574, 0.002356161, 0.002192256, 
    0.002110622, 0.002096619, 0.002067151, 0.002075161, 0.00204668, 
    0.001959166, 0.001898654, 0.001832231, 0.001798391, 0.00174586, 
    0.00175271, 0.001740997, 0.001757018, 0.001749563, 0.001885828, 
    0.001937388, 0.002050875, 0.001687384, 0.001063234, 0.0009256031, 
    0.00129787, 0.001292754, 0.00156447, 0.002030673, 0.002055675, 
    0.001679453, 0.001492104, 0.001517328, 0.001668549, 0.001680549, 
    0.001791525, 0.001840607, 0.001882887, 0.001840751, 0.001692263, 
    0.001619562, 0.001508299, 0.00134457, 0.001164595, 0.001052697, 
    0.0009955568, 0.001029746, 0.001089302, 0.001149193, 0.001207222, 
    0.001252697, 0.001324683, 0.001382191, 0.001463046, 0.001526942, 
    0.001456783, 0.001342393, 0.001293692, 0.001228396, 0.001186625, 
    0.001145824, 0.001096122, 0.001008733, 0.0009675343, 0.0008508507, 
    0.001165944, 0.001896541, 0.001149892, 0.001613522, 0.002218135, 
    0.002350328, 0.002854568, 0.003064313, 0.002844602, 0.002911805, 
    0.002418738, 0.002261843, 0.001968032, 0.001833946, 0.001710939, 
    0.001576121, 0.001461443, 0.001338594, 0.001246436, 0.001225201, 
    0.001168728,
  0.001582162, 0.00161101, 0.001787551, 0.002095795, 0.001953488, 
    0.002455219, 0.003412483, 0.003378168, 0.003185365, 0.002608679, 
    0.002905337, 0.003100917, 0.002802847, 0.002143651, 0.002138183, 
    0.002138739, 0.002125135, 0.0021931, 0.002210727, 0.002203082, 
    0.002152885, 0.002137182, 0.002116376, 0.002099656, 0.00208446, 
    0.002085652, 0.002044357, 0.002086971, 0.002150947, 0.002317172, 
    0.002485529, 0.002330921, 0.001972975, 0.0009961913, 0.001511747, 
    0.001755793, 0.001830165, 0.002195293, 0.00253744, 0.002051844, 
    0.001830448, 0.001845119, 0.001942584, 0.002027811, 0.002086638, 
    0.002166523, 0.002191477, 0.002140822, 0.002078769, 0.00197339, 
    0.0018922, 0.001678959, 0.001502019, 0.001430064, 0.001461186, 
    0.00154236, 0.001648202, 0.001797579, 0.001944237, 0.002009961, 
    0.00204307, 0.002047855, 0.00205852, 0.002050269, 0.001912862, 
    0.001790888, 0.001659153, 0.001600629, 0.001499208, 0.001453527, 
    0.001347559, 0.001294485, 0.0012609, 0.001212804, 0.001235422, 
    0.001470662, 0.002138295, 0.001901214, 0.002138104, 0.002499133, 
    0.002571518, 0.003485455, 0.003614948, 0.003420924, 0.003380901, 
    0.002937568, 0.002135418, 0.001950325, 0.001772831, 0.001622786, 
    0.001556808, 0.00148956, 0.001448123, 0.001425124, 0.001456722, 
    0.001469055,
  0.001981177, 0.001973198, 0.002131444, 0.002283492, 0.002369055, 
    0.00269874, 0.003604298, 0.003192057, 0.003144962, 0.002761537, 
    0.002423587, 0.003061373, 0.002932991, 0.002146657, 0.002221694, 
    0.002349708, 0.002369672, 0.002520687, 0.002575475, 0.002646476, 
    0.002644075, 0.002633442, 0.00255583, 0.002529858, 0.002508511, 
    0.00252776, 0.002543114, 0.002606946, 0.002702059, 0.002825353, 
    0.002963828, 0.003069481, 0.003027645, 0.003129845, 0.003157487, 
    0.002528031, 0.002343527, 0.002387219, 0.002452435, 0.002150469, 
    0.00223201, 0.002389635, 0.002455773, 0.002536947, 0.002610588, 
    0.002593819, 0.002611795, 0.002609663, 0.002527297, 0.002370162, 
    0.002302516, 0.002237841, 0.00227467, 0.002382293, 0.002487324, 
    0.002599029, 0.002696924, 0.002790272, 0.002926379, 0.002932912, 
    0.002854316, 0.002744084, 0.002607279, 0.002508861, 0.00232275, 
    0.002239098, 0.00211458, 0.002048506, 0.001941537, 0.001873236, 
    0.001794212, 0.001803382, 0.001753187, 0.001697684, 0.001716503, 
    0.001840465, 0.002185645, 0.002513298, 0.002412572, 0.002823128, 
    0.002980135, 0.003362939, 0.003549494, 0.002844491, 0.003350289, 
    0.002638195, 0.002204941, 0.002083682, 0.001958623, 0.00187969, 
    0.001873285, 0.001805844, 0.001851063, 0.001878991, 0.001898161, 
    0.00194041,
  0.002309511, 0.00236627, 0.002447222, 0.002797237, 0.002792642, 
    0.002643249, 0.003382363, 0.002935155, 0.002945565, 0.002710437, 
    0.002445442, 0.002717109, 0.002593135, 0.002347818, 0.002560185, 
    0.002645046, 0.002801877, 0.002931101, 0.003002752, 0.003043903, 
    0.003023002, 0.002999574, 0.002955182, 0.002949953, 0.002948046, 
    0.002931308, 0.002968693, 0.003084213, 0.003191531, 0.003241219, 
    0.003210304, 0.003355771, 0.003441984, 0.003285088, 0.003050787, 
    0.003265585, 0.002907719, 0.002717687, 0.002346959, 0.002635511, 
    0.00282694, 0.002912741, 0.002961142, 0.003003119, 0.002965305, 
    0.002957501, 0.003007522, 0.002992865, 0.002949093, 0.002882827, 
    0.002892651, 0.002975127, 0.003110742, 0.003248896, 0.003404854, 
    0.003429601, 0.003477016, 0.003504608, 0.003420336, 0.003299886, 
    0.003145168, 0.002995552, 0.002839422, 0.002756545, 0.002637066, 
    0.002553175, 0.002436494, 0.002377763, 0.002315409, 0.002322925, 
    0.002335737, 0.002248984, 0.00214133, 0.002103835, 0.002159927, 
    0.002492872, 0.002719895, 0.002321448, 0.002433809, 0.002899152, 
    0.002958518, 0.002813718, 0.003101697, 0.002754019, 0.002882781, 
    0.002264116, 0.002465564, 0.002383087, 0.002317443, 0.002294189, 
    0.002235156, 0.002238128, 0.002281028, 0.00231396, 0.002335768, 
    0.002380702,
  0.002630835, 0.002705031, 0.002671272, 0.002835844, 0.002070282, 
    0.00309405, 0.003489111, 0.003435847, 0.002880015, 0.002672003, 
    0.002388921, 0.002667423, 0.002622394, 0.002785506, 0.002932705, 
    0.003022686, 0.003172681, 0.003230475, 0.003262168, 0.003210956, 
    0.003238581, 0.003187798, 0.003174128, 0.003155977, 0.003176829, 
    0.003202882, 0.003179166, 0.003227709, 0.003191041, 0.003282005, 
    0.003368599, 0.003367819, 0.003380248, 0.003352355, 0.003330261, 
    0.003228441, 0.003139287, 0.003122423, 0.002865264, 0.003008347, 
    0.003177641, 0.003228918, 0.003283452, 0.003209526, 0.003041567, 
    0.003009014, 0.002951525, 0.002906224, 0.002899757, 0.003026914, 
    0.003186017, 0.003335951, 0.003473217, 0.003578534, 0.003706979, 
    0.003707726, 0.003662584, 0.003600294, 0.003485439, 0.003396954, 
    0.003280908, 0.003173176, 0.003112076, 0.00298832, 0.002878571, 
    0.002782106, 0.002706304, 0.002669602, 0.002637448, 0.00269373, 
    0.002641468, 0.00254758, 0.002569468, 0.002595646, 0.002734961, 
    0.003041409, 0.002257363, 0.00224053, 0.003002069, 0.003176877, 
    0.003139922, 0.002938857, 0.002454917, 0.003236625, 0.002581085, 
    0.002638894, 0.002417753, 0.002713792, 0.002788289, 0.002755325, 
    0.002672179, 0.002694955, 0.002692508, 0.002725344, 0.002696243, 
    0.002657951,
  0.002975225, 0.003005344, 0.003033843, 0.003020285, 0.002398252, 
    0.003312713, 0.003276205, 0.003198192, 0.003120388, 0.002522435, 
    0.002595422, 0.002733307, 0.00287299, 0.003024513, 0.003188482, 
    0.003261102, 0.003280081, 0.003300047, 0.003384316, 0.003296295, 
    0.003329735, 0.003288521, 0.003332071, 0.003362304, 0.003409209, 
    0.003372381, 0.003365373, 0.003346378, 0.003175752, 0.003231158, 
    0.003332516, 0.003329894, 0.003351558, 0.003323855, 0.003334854, 
    0.003317911, 0.00314226, 0.002882002, 0.002865804, 0.002964115, 
    0.00334827, 0.003286805, 0.00325322, 0.003144642, 0.003011988, 
    0.003026197, 0.003091509, 0.003331292, 0.003545839, 0.00377135, 
    0.004040478, 0.00412011, 0.004133111, 0.004053861, 0.003932362, 
    0.003843576, 0.003739022, 0.003632147, 0.003582554, 0.003477953, 
    0.003387162, 0.003300108, 0.003228886, 0.003123997, 0.003107624, 
    0.003038181, 0.002977991, 0.002942959, 0.00292816, 0.002967721, 
    0.002944722, 0.002964463, 0.003010906, 0.002981216, 0.003116243, 
    0.003239185, 0.002425732, 0.003544916, 0.003692752, 0.002984013, 
    0.003166975, 0.002844093, 0.002384997, 0.002774334, 0.003108565, 
    0.002888678, 0.00305592, 0.00306889, 0.003148505, 0.003079889, 
    0.003040232, 0.003000338, 0.002992216, 0.003001515, 0.00295588, 
    0.002995282,
  0.003231604, 0.003326382, 0.003328703, 0.003022302, 0.003279509, 
    0.003034478, 0.003462106, 0.002927602, 0.002702234, 0.002539458, 
    0.002903874, 0.002835685, 0.002973078, 0.003193233, 0.003278937, 
    0.003247546, 0.003235672, 0.003173096, 0.003189085, 0.003138825, 
    0.003230633, 0.003250264, 0.003300315, 0.003377913, 0.003505642, 
    0.003351623, 0.003423577, 0.003215104, 0.003268924, 0.003434321, 
    0.003202278, 0.00316405, 0.003092462, 0.003322424, 0.003490971, 
    0.003291588, 0.002917511, 0.002774188, 0.002928795, 0.003253775, 
    0.003305783, 0.00313366, 0.003045669, 0.003067937, 0.003175639, 
    0.003406428, 0.003739864, 0.00408759, 0.00434087, 0.004301276, 
    0.004168365, 0.004010739, 0.003904467, 0.00383825, 0.003726846, 
    0.003660373, 0.003633291, 0.003565788, 0.003542345, 0.003472693, 
    0.00343984, 0.00336884, 0.003347905, 0.00333856, 0.00337998, 0.003323887, 
    0.003294704, 0.003261596, 0.00326851, 0.00321272, 0.003218649, 
    0.003183331, 0.003093304, 0.003047829, 0.002987526, 0.003161889, 
    0.002770295, 0.003571747, 0.003368344, 0.002690092, 0.00256074, 
    0.002064831, 0.001978795, 0.002446856, 0.002800065, 0.003309295, 
    0.003284927, 0.003385255, 0.003340894, 0.003299393, 0.003289664, 
    0.003212595, 0.003212072, 0.003225865, 0.003165051, 0.003243046,
  0.003414454, 0.003539911, 0.003312141, 0.003015978, 0.003245147, 
    0.003603663, 0.003716165, 0.003170425, 0.003043586, 0.003275472, 
    0.00289367, 0.003127636, 0.003192294, 0.003221208, 0.003440266, 
    0.003490748, 0.003521202, 0.003313523, 0.003213387, 0.003030043, 
    0.00303982, 0.003058845, 0.003032111, 0.003034463, 0.003117925, 
    0.003067762, 0.003182346, 0.00304462, 0.003325334, 0.003277047, 
    0.003105892, 0.002959297, 0.002904156, 0.003074676, 0.003115524, 
    0.002983904, 0.00281035, 0.002897657, 0.003161652, 0.003310377, 
    0.003219746, 0.003142497, 0.00312751, 0.003236895, 0.003365245, 
    0.003624817, 0.003953408, 0.004252639, 0.004565347, 0.00456012, 
    0.004405465, 0.004287178, 0.004193081, 0.004056534, 0.004000235, 
    0.003920762, 0.003872506, 0.003817797, 0.003753964, 0.00371162, 
    0.003637377, 0.003580252, 0.003593763, 0.003534365, 0.003546523, 
    0.003518755, 0.003519772, 0.003460914, 0.003410878, 0.003281942, 
    0.003243651, 0.003103144, 0.00291441, 0.002872162, 0.002619075, 
    0.002852756, 0.003016597, 0.00298387, 0.00314663, 0.00241939, 
    0.002676723, 0.001526435, 0.001861698, 0.003127953, 0.003096245, 
    0.003134424, 0.003167341, 0.003285248, 0.003239535, 0.00328299, 
    0.003274836, 0.003267588, 0.003317624, 0.003348414, 0.003340544, 
    0.003311314,
  0.003198272, 0.003437549, 0.003158933, 0.003167627, 0.003226707, 
    0.003568616, 0.003674649, 0.003202215, 0.003114684, 0.003204582, 
    0.002894844, 0.002881175, 0.003186733, 0.003213007, 0.003306752, 
    0.003478684, 0.003631845, 0.003713161, 0.003766187, 0.003486235, 
    0.003262503, 0.003070369, 0.002995552, 0.002899025, 0.002880936, 
    0.002945628, 0.00278018, 0.00286188, 0.003162477, 0.003108896, 
    0.003187781, 0.002964653, 0.002865281, 0.00300126, 0.003094813, 
    0.002986016, 0.002955562, 0.003101427, 0.003202356, 0.003243491, 
    0.003196444, 0.003201546, 0.003115747, 0.003005043, 0.002982026, 
    0.003094606, 0.003184428, 0.003318259, 0.003632067, 0.003837997, 
    0.004018001, 0.004106058, 0.004225807, 0.004230529, 0.00421481, 
    0.004112162, 0.003988869, 0.003925528, 0.003860027, 0.003764754, 
    0.003712524, 0.003705848, 0.003659088, 0.003549129, 0.003522219, 
    0.003420765, 0.003384667, 0.00342105, 0.003404871, 0.003386004, 
    0.003259307, 0.003075281, 0.002949825, 0.00297934, 0.002888408, 
    0.00303106, 0.002964669, 0.002967229, 0.003042696, 0.001786388, 
    0.002378874, 0.002663182, 0.00301604, 0.003204422, 0.003210336, 
    0.003191691, 0.003202628, 0.003251281, 0.003055174, 0.003097326, 
    0.003035035, 0.003054442, 0.003103429, 0.00313131, 0.003032699, 
    0.003044238,
  0.003415709, 0.003387496, 0.003289554, 0.002794835, 0.002538679, 
    0.003197651, 0.003395349, 0.002830488, 0.002447698, 0.002310324, 
    0.002866202, 0.003557633, 0.003666779, 0.003438279, 0.003253235, 
    0.003375353, 0.003636707, 0.003699794, 0.003659263, 0.003458085, 
    0.003277125, 0.003151622, 0.003174638, 0.003026199, 0.002993422, 
    0.003024956, 0.002907291, 0.002934471, 0.002957534, 0.002931688, 
    0.003110899, 0.00327277, 0.003269637, 0.002964828, 0.003103143, 
    0.003117671, 0.003165863, 0.00315569, 0.003178466, 0.003161063, 
    0.003066044, 0.003015596, 0.00301992, 0.00298476, 0.002968991, 
    0.002997968, 0.002869477, 0.002816644, 0.002966275, 0.003028184, 
    0.003080286, 0.003047654, 0.00309553, 0.003150016, 0.003187973, 
    0.003192056, 0.003102031, 0.003083322, 0.003157645, 0.003184952, 
    0.00326344, 0.003290588, 0.003311109, 0.003238454, 0.003249707, 
    0.00321717, 0.003292145, 0.003494835, 0.003486264, 0.003568584, 
    0.003527496, 0.003436659, 0.003367374, 0.003252884, 0.003051549, 
    0.003165321, 0.003024116, 0.00285336, 0.003170392, 0.002792133, 
    0.002939587, 0.002895847, 0.002962952, 0.002873847, 0.002889743, 
    0.002970392, 0.002978895, 0.00310985, 0.003096452, 0.003137507, 
    0.0030248, 0.003053391, 0.003126143, 0.003098948, 0.003183791, 0.003344629,
  0.002712296, 0.002572518, 0.002200746, 0.001785406, 0.002009551, 
    0.002406692, 0.002581628, 0.002300469, 0.001480707, 0.002276069, 
    0.003534508, 0.00373279, 0.004057851, 0.004050284, 0.003670435, 
    0.003604839, 0.003596954, 0.003634021, 0.003465634, 0.003378691, 
    0.003108261, 0.003161794, 0.00314315, 0.003046401, 0.003018185, 
    0.002903538, 0.002739824, 0.002746312, 0.002748328, 0.002718259, 
    0.002960442, 0.003278874, 0.003325015, 0.003017375, 0.003137603, 
    0.003212513, 0.003199767, 0.003089236, 0.003058782, 0.003045382, 
    0.00294175, 0.003021143, 0.003089774, 0.00312786, 0.003151668, 
    0.003128622, 0.00311392, 0.003159838, 0.003258115, 0.003251806, 
    0.003259435, 0.003254825, 0.003246846, 0.003269909, 0.003276108, 
    0.003257971, 0.003232382, 0.003203597, 0.003254283, 0.003246576, 
    0.003236864, 0.003198987, 0.003193678, 0.003175909, 0.00328752, 
    0.003476681, 0.003584128, 0.003774466, 0.00380131, 0.00386834, 
    0.00389323, 0.003682913, 0.00308647, 0.002844762, 0.002747597, 
    0.002820266, 0.002818709, 0.002842013, 0.002766211, 0.002818996, 
    0.002866838, 0.002718065, 0.002713392, 0.002659112, 0.002741683, 
    0.002789972, 0.00281623, 0.002913872, 0.00296111, 0.002952112, 
    0.00305476, 0.003181472, 0.003448438, 0.003118465, 0.002990037, 
    0.002711151,
  0.00126365, 0.00130693, 0.001447011, 0.001420816, 0.001065158, 0.001399532, 
    0.001469501, 0.001323986, 0.001107566, 0.001547782, 0.003401293, 
    0.003617618, 0.002806154, 0.003046607, 0.003646038, 0.003705403, 
    0.003384111, 0.003461011, 0.003486726, 0.003567979, 0.003422862, 
    0.003258273, 0.003046796, 0.003011432, 0.002922596, 0.002807854, 
    0.002741304, 0.002668521, 0.002622873, 0.002722707, 0.003076123, 
    0.003378343, 0.003421353, 0.003182489, 0.00314709, 0.003145978, 
    0.003068127, 0.002989687, 0.002981756, 0.002984045, 0.003037563, 
    0.003179993, 0.003115239, 0.003037959, 0.003067032, 0.003072578, 
    0.003122963, 0.003176179, 0.003198668, 0.003198527, 0.003176417, 
    0.003164193, 0.003206061, 0.003235037, 0.003216583, 0.003158838, 
    0.003181249, 0.003213387, 0.003221795, 0.003172651, 0.003184348, 
    0.003154801, 0.003052058, 0.002999956, 0.003100568, 0.003363688, 
    0.003595876, 0.003621513, 0.003543582, 0.003086644, 0.003094655, 
    0.002885133, 0.002647826, 0.00303432, 0.003117036, 0.002979627, 
    0.002807805, 0.002801385, 0.002881335, 0.002762778, 0.002740858, 
    0.002690712, 0.002568353, 0.002543796, 0.002545942, 0.002450954, 
    0.002539329, 0.002500281, 0.002564158, 0.002559882, 0.002785442, 
    0.002906622, 0.00231107, 0.001547241, 0.001230159, 0.001213598,
  0.001010465, 0.001129324, 0.001078955, 0.001312668, 0.0005437841, 
    0.001064618, 0.001034513, 0.001145235, 0.0009395909, 0.001403554, 
    0.003288537, 0.00260547, 0.001954778, 0.002139362, 0.003001483, 
    0.003853447, 0.003311951, 0.00332031, 0.00360317, 0.003616823, 
    0.003574035, 0.003458292, 0.003140304, 0.003103619, 0.0030258, 
    0.002782185, 0.002441896, 0.002185708, 0.002497546, 0.002629279, 
    0.002865694, 0.003117956, 0.003341196, 0.003194092, 0.003022335, 
    0.003010001, 0.002938824, 0.002908912, 0.002940303, 0.003051136, 
    0.003063709, 0.003060132, 0.00301221, 0.003013449, 0.003048895, 
    0.003065648, 0.003045732, 0.003077712, 0.003141323, 0.003115842, 
    0.003077408, 0.003009841, 0.002973666, 0.002864121, 0.002813431, 
    0.002746819, 0.002724677, 0.002765257, 0.002740985, 0.002713695, 
    0.002740381, 0.002696417, 0.002519241, 0.002372408, 0.002366379, 
    0.002576252, 0.003130244, 0.003256159, 0.002590256, 0.002291648, 
    0.0026635, 0.002706319, 0.002581069, 0.003146615, 0.003163416, 
    0.003030552, 0.002919957, 0.002810238, 0.002758723, 0.002735121, 
    0.00271681, 0.002591878, 0.002562743, 0.002525326, 0.002412716, 
    0.002337743, 0.002332687, 0.002232265, 0.002271254, 0.002191446, 
    0.002310878, 0.002433647, 0.001232097, 0.0005111047, 0.0004476379, 
    0.0006450329,
  0.001269071, 0.001087235, 0.0006033732, 0.000627453, 0.0007280654, 
    0.0008432064, 0.0003983646, 0.000759155, 0.0009538482, 0.001487097, 
    0.002907034, 0.002022186, 0.00186038, 0.002008787, 0.002380068, 
    0.003228648, 0.003194856, 0.003274901, 0.003662012, 0.003624946, 
    0.003481402, 0.003604791, 0.003089966, 0.002686467, 0.002678202, 
    0.002769819, 0.002377603, 0.002148294, 0.002148532, 0.002289883, 
    0.00254518, 0.002495922, 0.002927223, 0.003059784, 0.002958439, 
    0.002947934, 0.002928318, 0.002828961, 0.002766861, 0.00291813, 
    0.003001878, 0.003017869, 0.003048133, 0.003000211, 0.002956802, 
    0.00300671, 0.003026085, 0.003025005, 0.003018487, 0.002985142, 
    0.002950553, 0.00285716, 0.002772713, 0.00262982, 0.002524516, 
    0.002382516, 0.002272652, 0.002324087, 0.002295619, 0.00225288, 
    0.002238526, 0.002194674, 0.002133288, 0.001942172, 0.001828779, 
    0.001955653, 0.002544655, 0.002937854, 0.00231533, 0.002144495, 
    0.002778195, 0.003052646, 0.002837401, 0.002953559, 0.002961379, 
    0.00289122, 0.002835939, 0.00295685, 0.002950571, 0.002888424, 
    0.002869954, 0.00274162, 0.002673622, 0.002574904, 0.002490202, 
    0.00235338, 0.00225787, 0.002233361, 0.002195626, 0.002094029, 
    0.002091564, 0.002070917, 0.001246149, 0.00103194, 0.001082882, 
    0.0009065457,
  0.0006555542, 0.001256323, 0.001183924, 0.0009088186, 0.001447663, 
    0.001451985, 0.0007916759, 0.0006894898, 0.001161051, 0.001171652, 
    0.00132327, 0.00115563, 0.001689577, 0.001782115, 0.002339634, 
    0.002503713, 0.002210729, 0.002164538, 0.003085916, 0.003225023, 
    0.002935853, 0.002830583, 0.002369833, 0.001877516, 0.001887177, 
    0.00210622, 0.00204787, 0.00195662, 0.001797213, 0.001767318, 
    0.001885396, 0.001865082, 0.002188188, 0.002665743, 0.002695721, 
    0.002738805, 0.002804199, 0.0027743, 0.002676867, 0.002678996, 
    0.002750266, 0.002913853, 0.003018696, 0.00303551, 0.00294248, 
    0.002908371, 0.00293857, 0.002953287, 0.002918577, 0.002889633, 
    0.002912058, 0.002845922, 0.002736629, 0.002525025, 0.002327505, 
    0.00213963, 0.001991017, 0.001972642, 0.001901943, 0.001865481, 
    0.001813632, 0.001756475, 0.001703943, 0.001571733, 0.001553423, 
    0.001812328, 0.002133098, 0.002542082, 0.00213669, 0.002518002, 
    0.003114572, 0.003040692, 0.00286461, 0.0027695, 0.002490423, 
    0.002543321, 0.002523929, 0.002651069, 0.002799176, 0.002848973, 
    0.002884943, 0.002816133, 0.002686534, 0.002622539, 0.002531113, 
    0.002306014, 0.002252609, 0.002261193, 0.002130935, 0.002071426, 
    0.001992382, 0.002048284, 0.002004112, 0.001186146, 0.0007886887, 
    0.0002217598,
  0.0006451607, 0.0005879868, 0.0003027422, 0.001418145, 0.001732045, 
    0.001987344, 0.001380666, 0.001081545, 0.002249812, 0.001782878, 
    0.001343901, 0.001225645, 0.001717425, 0.001746114, 0.001403824, 
    0.001421116, 0.001387118, 0.001430559, 0.00216643, 0.002594027, 
    0.002175697, 0.001445324, 0.001514179, 0.001293324, 0.001388915, 
    0.001531966, 0.001649236, 0.00194446, 0.001883029, 0.001671027, 
    0.001612518, 0.001598819, 0.001853973, 0.002144414, 0.002323101, 
    0.002533815, 0.002580148, 0.002533418, 0.002519304, 0.002408646, 
    0.002358895, 0.002460083, 0.002547296, 0.00259215, 0.002641266, 
    0.002707209, 0.002771804, 0.002828722, 0.002840326, 0.002839436, 
    0.002874753, 0.00283241, 0.002751237, 0.002640294, 0.002469618, 
    0.00224118, 0.001965171, 0.001829383, 0.001730138, 0.001664875, 
    0.001657454, 0.001598375, 0.001495807, 0.00144771, 0.001659966, 
    0.002114519, 0.002010822, 0.001892202, 0.002004081, 0.002533801, 
    0.002282286, 0.002326678, 0.002196344, 0.002051783, 0.002254311, 
    0.002431534, 0.002424447, 0.002283508, 0.002336007, 0.002435159, 
    0.002519175, 0.002486225, 0.002402956, 0.002374106, 0.002336976, 
    0.002206372, 0.002164934, 0.002115089, 0.00208279, 0.002079088, 
    0.001942203, 0.001894965, 0.001908428, 0.001927707, 0.001434913, 
    0.0006053452,
  0.001312889, 0.001373893, 0.001503911, 0.002433552, 0.00232717, 
    0.002008229, 0.001631753, 0.001588233, 0.002042944, 0.002150534, 
    0.001476495, 0.001305357, 0.001346444, 0.001368443, 0.001327641, 
    0.001260041, 0.001396925, 0.001275062, 0.001285727, 0.00143423, 
    0.001103575, 0.001025628, 0.001120408, 0.0009933624, 0.001032526, 
    0.000949637, 0.001118261, 0.001773913, 0.001975472, 0.001679563, 
    0.001420737, 0.001459074, 0.001591363, 0.001799787, 0.001771496, 
    0.002057504, 0.001745985, 0.001785517, 0.002159228, 0.002171785, 
    0.002019514, 0.00197067, 0.001946351, 0.001950867, 0.00202492, 
    0.002145574, 0.00226817, 0.002356401, 0.002428609, 0.002483859, 
    0.002531511, 0.002511007, 0.002470729, 0.002412492, 0.002287704, 
    0.002091662, 0.001839224, 0.001681169, 0.001564678, 0.001484029, 
    0.001502212, 0.001463508, 0.00147171, 0.001543999, 0.00150396, 
    0.001428175, 0.001542394, 0.00160826, 0.001750422, 0.001394049, 
    0.001701816, 0.001922637, 0.001597482, 0.002020882, 0.002110685, 
    0.002118411, 0.002311435, 0.002243263, 0.002184881, 0.002195277, 
    0.00223719, 0.002165999, 0.002091135, 0.002038286, 0.002004098, 
    0.00193648, 0.001830338, 0.001856277, 0.001963614, 0.00198488, 
    0.001923209, 0.001787329, 0.001666737, 0.001861253, 0.001971131, 
    0.001444785,
  0.001679135, 0.002276722, 0.002346039, 0.002382597, 0.00222915, 
    0.001770608, 0.0009094374, 0.0006047729, 0.0007919311, 0.0007546423, 
    0.0008220188, 0.001015741, 0.001236486, 0.001525384, 0.001578615, 
    0.00106689, 0.0007726182, 0.0007198006, 0.001039297, 0.0009098677, 
    0.0009306737, 0.0009246334, 0.0007685969, 0.0008400907, 0.0009444223, 
    0.0009608581, 0.0008514868, 0.001110252, 0.001390663, 0.001361305, 
    0.001127004, 0.001050122, 0.001108359, 0.001103559, 0.001166295, 
    0.001646424, 0.001683648, 0.001439731, 0.00175549, 0.001814109, 
    0.001755252, 0.001680341, 0.001682962, 0.001723589, 0.001705422, 
    0.001687811, 0.001744745, 0.001797006, 0.001802172, 0.001789631, 
    0.001793844, 0.001834677, 0.001881899, 0.0019042, 0.00189808, 
    0.001818578, 0.001710971, 0.001605097, 0.001459519, 0.001355203, 
    0.001332395, 0.001291513, 0.001356456, 0.001304038, 0.001123253, 
    0.001137796, 0.001263109, 0.001244512, 0.00122059, 0.001104721, 
    0.001296648, 0.001658692, 0.001506281, 0.001804127, 0.00190075, 
    0.001854815, 0.001917011, 0.002407456, 0.002403783, 0.002273844, 
    0.002133177, 0.002063892, 0.002050477, 0.001951279, 0.001798421, 
    0.001637266, 0.001442273, 0.00138936, 0.001534001, 0.001654434, 
    0.001773643, 0.001736498, 0.001604271, 0.00159785, 0.0013923, 0.001249695,
  0.001479038, 0.002138916, 0.002175268, 0.001647823, 0.001958577, 
    0.001339436, 0.0006390414, 0.0002903612, 0.000618536, 0.0006192834, 
    0.0005969987, 0.0007952522, 0.0008712769, 0.001170538, 0.000636498, 
    0.000267616, 0.0002803637, 0.0004342545, 0.0006151826, 0.0006732454, 
    0.0007131721, 0.0007593937, 0.0008830535, 0.0009289884, 0.0008427771, 
    0.000792089, 0.0008405678, 0.0008878857, 0.0009529416, 0.0009632092, 
    0.0008998376, 0.0008117505, 0.0007967786, 0.000757406, 0.0007251091, 
    0.000829394, 0.001274253, 0.001418734, 0.001228427, 0.001433405, 
    0.001403555, 0.00138882, 0.001355855, 0.001368364, 0.001386977, 
    0.001383576, 0.001391346, 0.001383543, 0.001371654, 0.001385577, 
    0.001409992, 0.001446674, 0.001464349, 0.001458007, 0.001432957, 
    0.001382365, 0.001336494, 0.001306756, 0.001261804, 0.001211896, 
    0.001189262, 0.001161288, 0.001239775, 0.001025948, 0.0008738665, 
    0.0008801925, 0.0009315321, 0.0009806789, 0.001053269, 0.001248837, 
    0.001186115, 0.001374244, 0.001623043, 0.001721446, 0.001952503, 
    0.00174098, 0.001771944, 0.001827162, 0.002096526, 0.002115184, 
    0.002023663, 0.001859981, 0.001749992, 0.001522953, 0.00134266, 
    0.001223087, 0.001002248, 0.0008351961, 0.0009603184, 0.001217699, 
    0.001463811, 0.001597452, 0.001591062, 0.001526642, 0.001117802, 
    0.0008435096,
  0.001258437, 0.001368269, 0.001397293, 0.001345953, 0.001272313, 
    0.00098931, 0.0007741451, 0.000640566, 0.00050249, 0.0003870162, 
    0.0004231599, 0.0006293762, 0.0006827503, 0.0005257279, 0.000843239, 
    0.0005154605, 0.0004415491, 0.0004566498, 0.000486627, 0.0005786885, 
    0.0006979126, 0.0006634702, 0.0005990972, 0.0006885678, 0.0006045967, 
    0.0005062411, 0.0005554189, 0.0006273894, 0.0006397397, 0.0006883449, 
    0.0007081656, 0.0006807791, 0.0006961173, 0.0007358538, 0.000671179, 
    0.0006289945, 0.0007034447, 0.001093736, 0.001126034, 0.001069434, 
    0.001005156, 0.001058132, 0.001085773, 0.001085598, 0.001092577, 
    0.00111502, 0.001123699, 0.001116753, 0.0011302, 0.001164326, 
    0.001190504, 0.001205731, 0.00120198, 0.00121781, 0.001250745, 
    0.001242066, 0.001196209, 0.001165088, 0.001136063, 0.001075838, 
    0.001053507, 0.001107534, 0.001230908, 0.001026933, 0.000861072, 
    0.0008097477, 0.0008334788, 0.0009276383, 0.001089063, 0.001117785, 
    0.0009015873, 0.001248072, 0.001386991, 0.001592938, 0.001573005, 
    0.001564979, 0.001515753, 0.001497601, 0.001481421, 0.001502657, 
    0.00156986, 0.001385881, 0.001012866, 0.0008681617, 0.000878382, 
    0.0009844294, 0.000849165, 0.0005777841, 0.0005360916, 0.0007105041, 
    0.0009481572, 0.00121579, 0.001355757, 0.001422086, 0.001486728, 
    0.00119772,
  0.001248486, 0.0012544, 0.001287779, 0.0012767, 0.001223771, 0.001134475, 
    0.001000849, 0.0008203024, 0.0006953389, 0.0006988831, 0.0007216763, 
    0.0006263573, 0.0005088961, 0.0005938038, 0.0006204117, 0.0005686912, 
    0.0005501416, 0.0005792442, 0.0005386977, 0.0005268089, 0.0005990341, 
    0.0006362901, 0.0006012425, 0.0005850464, 0.0004908075, 0.0003839324, 
    0.0003552267, 0.0004804283, 0.0005322923, 0.0006170264, 0.0006839423, 
    0.0006379278, 0.0006145625, 0.0006410589, 0.0006519943, 0.0006163747, 
    0.0005794992, 0.0005840603, 0.000721788, 0.0007844437, 0.0008702585, 
    0.0008959761, 0.0008947519, 0.0008930359, 0.0009017298, 0.0009481423, 
    0.001000959, 0.001033893, 0.001054937, 0.001068083, 0.001094547, 
    0.001129278, 0.001168314, 0.001191299, 0.001203188, 0.001186737, 
    0.001148606, 0.001123047, 0.00110399, 0.001062806, 0.00103124, 
    0.001084262, 0.0009844624, 0.0009211213, 0.0008125138, 0.0007716967, 
    0.0008577504, 0.000919072, 0.0008289334, 0.0007668012, 0.0009306744, 
    0.0009997995, 0.001074918, 0.001158062, 0.00127743, 0.00135463, 
    0.001334968, 0.001281244, 0.001212262, 0.001158205, 0.001264635, 
    0.00112845, 0.0008774269, 0.0008588145, 0.0008631228, 0.0008012615, 
    0.0005892124, 0.0002627685, 7.573655e-005, 0.0001621395, 0.0004438404, 
    0.0007699467, 0.0009959843, 0.001097042, 0.001222736, 0.001291082,
  0.001112891, 0.001121361, 0.001086887, 0.001090082, 0.001113588, 
    0.001133473, 0.001075267, 0.0009258259, 0.0008288692, 0.000790881, 
    0.0007141102, 0.0005428628, 0.0004385626, 0.0004197587, 0.0004366382, 
    0.0004528994, 0.0004795066, 0.0005556415, 0.0004792048, 0.0004094117, 
    0.0004353835, 0.0004891858, 0.0005284296, 0.0005532254, 0.0005420833, 
    0.0005089114, 0.0005052874, 0.0005358527, 0.0005613954, 0.000600623, 
    0.0005904823, 0.0006408521, 0.0006350507, 0.0006011636, 0.000548966, 
    0.0005420516, 0.0005409233, 0.000520753, 0.0006112726, 0.0006666975, 
    0.0007696776, 0.0008136262, 0.0005678162, 0.0007305453, 0.0007385407, 
    0.0008082697, 0.0008688597, 0.0009326451, 0.000991852, 0.001038868, 
    0.001080385, 0.001135904, 0.00118459, 0.001201247, 0.001166883, 
    0.001144918, 0.00115827, 0.001170827, 0.001151451, 0.001113893, 
    0.001031954, 0.0008604843, 0.0008044234, 0.0007672464, 0.0007331681, 
    0.0007191175, 0.000758965, 0.0007681842, 0.0007951735, 0.0008372301, 
    0.0008915574, 0.0009549775, 0.001028902, 0.001089858, 0.001133838, 
    0.001136207, 0.001142358, 0.00109504, 0.001044351, 0.001006142, 
    0.0009691231, 0.0007820604, 0.0007363632, 0.0006816857, 0.0006689224, 
    0.0006801751, 0.0005746833, 0.0003744126, 0.0002151649, 0.0002132105, 
    0.000377432, 0.0006090635, 0.0007806774, 0.0008967235, 0.0009872601, 
    0.001065922,
  0.0008303807, 0.0009541344, 0.0009009046, 0.0008835308, 0.000875758, 
    0.001001756, 0.0009721601, 0.0008809082, 0.0008131177, 0.0007476169, 
    0.0006729281, 0.0005915319, 0.00053075, 0.0004942878, 0.0004579532, 
    0.0004324587, 0.0004220954, 0.0004140688, 0.0003748569, 0.0003694049, 
    0.0003905445, 0.0004157852, 0.0004437277, 0.0004755009, 0.0005174151, 
    0.000535042, 0.0005547353, 0.0006131323, 0.0006564765, 0.0005960455, 
    0.0005727757, 0.0006046126, 0.0006438245, 0.0006329844, 0.0005845695, 
    0.0005593129, 0.0005592178, 0.0005385708, 0.0005715201, 0.0005811993, 
    0.0006518513, 0.0006855, 0.0005553553, 0.0005528757, 0.0006691772, 
    0.0007938221, 0.0009287982, 0.0009850976, 0.001062472, 0.001118262, 
    0.00114355, 0.00113182, 0.001101763, 0.001084501, 0.0009171003, 
    0.000999847, 0.00100212, 0.001029841, 0.001025852, 0.0009770398, 
    0.0007715211, 0.0007573119, 0.0007908016, 0.0007070852, 0.000681622, 
    0.0006546965, 0.0006330796, 0.0006470829, 0.0007110429, 0.0007791829, 
    0.0008180612, 0.0008649658, 0.0008468782, 0.0008749161, 0.0009334241, 
    0.001020479, 0.00108803, 0.001007873, 0.0009349172, 0.0008981372, 
    0.0006681429, 0.0006654258, 0.0005994793, 0.0005271272, 0.0005705985, 
    0.000593836, 0.0006165174, 0.0006046924, 0.0005446104, 0.0005478221, 
    0.0006043911, 0.0006741849, 0.0007340279, 0.0007470455, 0.0007952694, 
    0.0008363728,
  0.000735824, 0.0008347197, 0.0007474571, 0.0007012202, 0.00070157, 
    0.0007632719, 0.0007893406, 0.0007612053, 0.000694497, 0.0006399781, 
    0.0006032134, 0.0005523034, 0.0004947337, 0.0004401039, 0.0004083943, 
    0.0003802611, 0.0003717572, 0.0003735691, 0.0003823747, 0.0004099994, 
    0.0004437594, 0.0004497042, 0.0004576673, 0.0005097538, 0.0005670218, 
    0.0005955528, 0.0005985885, 0.0006284545, 0.0006457161, 0.0006357182, 
    0.0006312041, 0.0006714651, 0.0007185608, 0.0007258721, 0.0006954501, 
    0.000628947, 0.0005500464, 0.0004949716, 0.0004517704, 0.0004312347, 
    0.0004670608, 0.0005314179, 0.0005504121, 0.000580278, 0.0006154525, 
    0.0006817174, 0.0007519238, 0.0008092553, 0.000931866, 0.001032796, 
    0.001049359, 0.0009921701, 0.0008016413, 0.0007297024, 0.000675645, 
    0.0006497686, 0.0006702573, 0.0006959268, 0.0007316263, 0.0007146979, 
    0.0006559517, 0.000588893, 0.0005348672, 0.0004966885, 0.0005128847, 
    0.0005634136, 0.00060679, 0.0006411863, 0.000666522, 0.0006926528, 
    0.0007534337, 0.0007616188, 0.0007788008, 0.0007867799, 0.0008182193, 
    0.0008357351, 0.0009766412, 0.0009585056, 0.0007407179, 0.0006346852, 
    0.0005689447, 0.0005289384, 0.0004516754, 0.000369055, 0.0004374175, 
    0.0003935639, 0.0005626041, 0.0006563175, 0.0006988519, 0.000731817, 
    0.0007421812, 0.0007176716, 0.0006486573, 0.0005812328, 0.0006365143, 
    0.000698376,
  0.0005246801, 0.0005500475, 0.0005435306, 0.0006225412, 0.0006468128, 
    0.0006872173, 0.0006564762, 0.000685802, 0.0006712268, 0.0006704316, 
    0.000678506, 0.0006856592, 0.000673071, 0.0006408207, 0.000606742, 
    0.0005706619, 0.0005244405, 0.0004990408, 0.0004700173, 0.0004644387, 
    0.0004852447, 0.0004989137, 0.0005417496, 0.0005777985, 0.0005907365, 
    0.000595171, 0.000600162, 0.0006149758, 0.0006472578, 0.0007000593, 
    0.0007179409, 0.0007275888, 0.0007167009, 0.0006419329, 0.000560187, 
    0.0004978643, 0.0004388477, 0.0003912436, 0.0003463574, 0.0003362644, 
    0.0003761119, 0.0004353509, 0.0004897263, 0.0004897583, 0.0004783141, 
    0.0005037931, 0.000555689, 0.0006532025, 0.0008128474, 0.0009215026, 
    0.0009329468, 0.0008809399, 0.0006685725, 0.0005978416, 0.0005748104, 
    0.0005746039, 0.000584522, 0.0005850466, 0.0005674353, 0.0005540045, 
    0.0005499038, 0.0005394607, 0.0005102784, 0.0004931758, 0.0005040795, 
    0.0005317202, 0.0005835523, 0.0006266902, 0.0006712903, 0.0007566127, 
    0.000841283, 0.0008908105, 0.0008882674, 0.0008910964, 0.0008401545, 
    0.0007895622, 0.0007494602, 0.0008927016, 0.0008308083, 0.0007832518, 
    0.000553146, 0.0004915704, 0.0005110095, 0.0003202269, 0.0002706834, 
    0.0002823501, 0.0003293187, 0.0003478832, 0.0004453971, 0.0005296534, 
    0.0005537653, 0.0006597354, 0.000562238, 0.0004317588, 0.0004124474, 
    0.0004378627,
  0.0005383007, 0.0005495218, 0.0005647014, 0.0005684206, 0.0005250447, 
    0.0006682705, 0.0006689064, 0.0006524392, 0.0006432203, 0.0006521686, 
    0.0006323014, 0.0006119879, 0.0005887335, 0.0005949333, 0.0006422191, 
    0.0006615948, 0.0006835291, 0.0006882185, 0.0006606887, 0.0006103665, 
    0.0005945193, 0.0005815654, 0.000582074, 0.0005801987, 0.0005840608, 
    0.000560203, 0.0005635569, 0.000582233, 0.000616152, 0.0006465266, 
    0.0006842921, 0.0006824324, 0.0006396761, 0.0005680071, 0.0004988022, 
    0.0004742927, 0.0004704462, 0.0004779167, 0.0005223738, 0.0005649235, 
    0.0006202048, 0.0006592897, 0.0006795237, 0.0006744056, 0.0005950598, 
    0.0005833457, 0.0006120827, 0.0007231225, 0.0008829265, 0.00137747, 
    0.001192823, 0.001041793, 0.0009564552, 0.0007890213, 0.000730418, 
    0.000683243, 0.0006903954, 0.0007050504, 0.0006780612, 0.0006320941, 
    0.0006091741, 0.000644794, 0.0006888696, 0.0007142372, 0.000742498, 
    0.0007499685, 0.0007756064, 0.0008326201, 0.0008992348, 0.0007453114, 
    0.0008675727, 0.0007985741, 0.0007774659, 0.0006823053, 0.0008550314, 
    0.001002947, 0.0009509552, 0.000916909, 0.0008508512, 0.0006414724, 
    0.000518925, 0.0004622447, 0.0004634369, 0.0003156014, 0.0002314556, 
    0.0001885244, 0.000184058, 0.0002276249, 0.0003047612, 0.0004197266, 
    0.000522994, 0.0005793402, 0.0005441012, 0.0005292092, 0.0005142684, 
    0.0005414477,
  0.0006697811, 0.0006417581, 0.000622144, 0.0006077909, 0.000597714, 
    0.000631188, 0.0007081027, 0.0007804707, 0.0007942193, 0.0007564537, 
    0.0006969757, 0.0006536311, 0.0006452554, 0.0006703048, 0.0006859768, 
    0.0009164482, 0.0009892136, 0.001022576, 0.001019572, 0.0008429677, 
    0.0007506199, 0.0007007429, 0.0006626121, 0.0006351301, 0.0006088562, 
    0.0005899101, 0.0005839334, 0.0005830911, 0.0005936609, 0.0006441262, 
    0.0006853411, 0.0007309744, 0.0007616033, 0.0007820755, 0.0007822184, 
    0.0008835942, 0.0008869637, 0.0008998702, 0.0007990984, 0.0008201112, 
    0.001057767, 0.001059563, 0.001071484, 0.001121218, 0.001159603, 
    0.001177246, 0.001189708, 0.001235055, 0.001317532, 0.001433387, 
    0.001499461, 0.001451634, 0.001352245, 0.001252762, 0.001202773, 
    0.001179535, 0.001176293, 0.001182746, 0.001176293, 0.001161717, 
    0.001151847, 0.00113662, 0.001106595, 0.0009285756, 0.0008864868, 
    0.0008590368, 0.0008526632, 0.0008545546, 0.0008343208, 0.0007402408, 
    0.0007720618, 0.0007573116, 0.0007318647, 0.0008172025, 0.0008974543, 
    0.0009423405, 0.0009916296, 0.001270357, 0.001060532, 0.0007649572, 
    0.0005362502, 0.0004887093, 0.0003070661, 0.0002541689, 0.0002127795, 
    0.0001844077, 0.0001715013, 0.000187078, 0.000238783, 0.0003303993, 
    0.0004841155, 0.0008970089, 0.0008820682, 0.0007395258, 0.0006752473, 
    0.0006892197,
  0.0006155162, 0.0005801977, 0.0005906245, 0.0006284376, 0.0006207451, 
    0.000652153, 0.0007067034, 0.0007645439, 0.0007796595, 0.0008032313, 
    0.0008550477, 0.0009167506, 0.0009910732, 0.001070546, 0.00113139, 
    0.001174385, 0.001197464, 0.00119047, 0.00115946, 0.001102574, 
    0.001023879, 0.0009524334, 0.000886916, 0.0008304267, 0.0008088577, 
    0.0006941785, 0.0006973733, 0.0007169711, 0.0007268892, 0.0007568505, 
    0.0007860647, 0.0009784529, 0.001011577, 0.001022083, 0.001053507, 
    0.001040028, 0.0009906599, 0.0009401469, 0.000894625, 0.0008622953, 
    0.0008502791, 0.0008450657, 0.0008485943, 0.0008563827, 0.0008621365, 
    0.0008623272, 0.0008605312, 0.0008632015, 0.0008737395, 0.0008872023, 
    0.0009051469, 0.0009221385, 0.0009367933, 0.0009434054, 0.0009466956, 
    0.0009482056, 0.0009533394, 0.0009634325, 0.0009826968, 0.001007111, 
    0.001034465, 0.001053332, 0.001056924, 0.001048659, 0.001028521, 
    0.000805059, 0.0007548638, 0.0007153183, 0.0006943057, 0.000694258, 
    0.0007093257, 0.0007747319, 0.0008162009, 0.0008408059, 0.000842745, 
    0.001248263, 0.001256385, 0.001159158, 0.000604358, 0.0004916021, 
    0.0003823587, 0.0002912986, 0.0002193281, 0.0001665899, 0.0001372962, 
    0.0001305568, 0.0001439083, 0.0001795439, 0.0002370664, 0.0003171432, 
    0.000420601, 0.0005652099, 0.0009423243, 0.0009936956, 0.0009722066, 
    0.00079894,
  0.0008837847, 0.000908612, 0.0009118547, 0.0008720706, 0.0007538464, 
    0.0007566758, 0.0007609993, 0.0009392885, 0.0009429124, 0.00093576, 
    0.0009400676, 0.0009477128, 0.000965451, 0.0009819657, 0.0009885936, 
    0.0009849378, 0.0009703942, 0.0009447562, 0.0009290525, 0.0009106308, 
    0.0008919227, 0.0008710851, 0.0008513599, 0.0008248001, 0.0007942189, 
    0.0006690013, 0.0006723868, 0.0007991939, 0.0008115759, 0.0008343051, 
    0.0008519004, 0.0008601338, 0.0008597523, 0.000847291, 0.0008246094, 
    0.000794219, 0.0007624933, 0.0007297187, 0.0006977865, 0.0006712743, 
    0.0006491967, 0.0006298531, 0.0006155161, 0.0006028641, 0.0005939949, 
    0.0005873828, 0.0005824872, 0.0005812157, 0.0005835681, 0.0005874147, 
    0.0005903392, 0.0005913723, 0.0005921035, 0.0005922942, 0.000591865, 
    0.0005909113, 0.0005943445, 0.0006041196, 0.0006228913, 0.0006482113, 
    0.00067795, 0.0007074981, 0.0007327227, 0.0007491576, 0.0007519869, 
    0.0007333267, 0.0007175275, 0.0006927479, 0.0006643126, 0.0006399938, 
    0.0006215084, 0.0004879622, 0.0004722266, 0.0004300106, 0.0003999221, 
    0.0003708828, 0.0003392208, 0.0003070661, 0.0002759922, 0.0002433766, 
    0.0002136219, 0.0001898277, 0.0001727093, 0.0001612334, 0.000159024, 
    0.0001699754, 0.0001928794, 0.0002268779, 0.0002713192, 0.0003282376, 
    0.0003960756, 0.000471559, 0.0006792216, 0.0007493803, 0.0008107808, 
    0.0008580193,
  0.0006212383, 0.0006326347, 0.0006460021, 0.0006546963, 0.0006590038, 
    0.0006676345, 0.0006756614, 0.0006852457, 0.0006919374, 0.0006983428, 
    0.0007045259, 0.0007089127, 0.000711742, 0.0007158109, 0.0007187832, 
    0.0007215966, 0.0007213741, 0.0007204363, 0.0007194985, 0.000719419, 
    0.0007185608, 0.0007175753, 0.0007159061, 0.0007132994, 0.0007087377, 
    0.0007028251, 0.0007030634, 0.0006983428, 0.0006924777, 0.0006846576, 
    0.0006755659, 0.0006646622, 0.000651422, 0.000636497, 0.0006201256, 
    0.0006041992, 0.0005899894, 0.0005773691, 0.0005671647, 0.0005596943, 
    0.000555371, 0.0005544492, 0.0005560544, 0.0005589632, 0.0005623486, 
    0.0005652574, 0.0005675462, 0.0005695806, 0.0005702323, 0.000568325, 
    0.0005652892, 0.0005609023, 0.0005567698, 0.0005524146, 0.0005485523, 
    0.0005460409, 0.0005445786, 0.0005460887, 0.0005517312, 0.0005614746, 
    0.0005734591, 0.0005858408, 0.0005970783, 0.0006073463, 0.0006148327, 
    0.0006184566, 0.0006185044, 0.000614785, 0.0006071555, 0.0005967288, 
    0.0005870649, 0.0005726803, 0.0005616177, 0.000551922, 0.0005414156, 
    0.000539413, 0.0005338022, 0.0005254734, 0.0005188612, 0.0005143313, 
    0.0005028872, 0.0004942088, 0.0004890113, 0.0004880417, 0.0004908073, 
    0.0005019812, 0.0005152532, 0.0005302736, 0.0005424647, 0.0005504756, 
    0.0005604415, 0.0005698987, 0.0005842198, 0.0005953779, 0.0006035157, 
    0.0006102073,
  0.0005550691, 0.0005568652, 0.0005634456, 0.0005716154, 0.0005797058, 
    0.0005866994, 0.0005946308, 0.0006024509, 0.0006084113, 0.0006152619, 
    0.0006212065, 0.0006283112, 0.0006362426, 0.0006418217, 0.0006461926, 
    0.0006490854, 0.000652169, 0.0006537585, 0.0006551413, 0.0006553797, 
    0.0006543784, 0.0006530592, 0.0006514697, 0.0006491014, 0.0006442058, 
    0.0006374984, 0.0006303458, 0.0006223349, 0.0006128936, 0.0006022124, 
    0.0005911975, 0.0005800871, 0.0005679755, 0.0005555776, 0.0005437521, 
    0.0005315769, 0.0005212612, 0.0005118516, 0.0005023944, 0.0004941928, 
    0.0004856893, 0.0004782824, 0.0004714318, 0.0004651534, 0.0004602261, 
    0.0004560618, 0.0004523742, 0.000448782, 0.0004463343, 0.0004430441, 
    0.0004412003, 0.0004394042, 0.000438546, 0.0004381963, 0.0004381963, 
    0.0004387844, 0.0004408348, 0.0004437753, 0.000446827, 0.000449545, 
    0.0004528829, 0.0004576036, 0.0004627217, 0.0004679033, 0.0004722107, 
    0.0004767724, 0.0004830349, 0.0004893292, 0.0004954326, 0.0005007732, 
    0.0005056688, 0.0005102464, 0.0005130756, 0.0005162228, 0.0005193699, 
    0.0005211341, 0.0005233912, 0.000525537, 0.0005273649, 0.0005289225, 
    0.0005293516, 0.0005299557, 0.0005304802, 0.0005323399, 0.0005336591, 
    0.0005360592, 0.0005379824, 0.0005402236, 0.0005433706, 0.0005464224, 
    0.0005484728, 0.0005510319, 0.0005538929, 0.0005554506, 0.0005550374, 
    0.0005553552,
  5.821181e-005, 5.603426e-005, 5.409516e-005, 5.252159e-005, 5.07255e-005, 
    4.943804e-005, 4.818237e-005, 4.711744e-005, 4.622735e-005, 
    4.532134e-005, 4.463788e-005, 4.412925e-005, 4.365241e-005, 
    4.328684e-005, 4.301663e-005, 4.292125e-005, 4.292127e-005, 
    4.296892e-005, 4.293713e-005, 4.296892e-005, 4.30325e-005, 4.315966e-005, 
    4.339807e-005, 4.363649e-005, 4.382725e-005, 4.420872e-005, 4.45584e-005, 
    4.508292e-005, 4.548028e-005, 4.610016e-005, 4.692668e-005, 
    4.764194e-005, 4.859564e-005, 4.953342e-005, 5.066194e-005, 
    5.196528e-005, 5.328453e-005, 5.479452e-005, 5.639985e-005, 
    5.810056e-005, 6.00397e-005, 6.204241e-005, 6.421996e-005, 6.64611e-005, 
    6.873402e-005, 7.099105e-005, 7.318452e-005, 7.518724e-005, 
    7.736476e-005, 7.924033e-005, 8.100463e-005, 8.25146e-005, 8.338879e-005, 
    8.440603e-005, 8.50418e-005, 8.585246e-005, 8.639289e-005, 8.65995e-005, 
    8.640881e-005, 8.615447e-005, 8.604323e-005, 8.566174e-005, 
    8.547102e-005, 8.483525e-005, 8.462858e-005, 8.429482e-005, 
    8.410407e-005, 8.415175e-005, 8.419945e-005, 8.446965e-005, 
    8.488289e-005, 8.540743e-005, 8.613861e-005, 8.597964e-005, 
    8.752142e-005, 8.861814e-005, 8.923802e-005, 9.015991e-005, 
    9.120896e-005, 9.182884e-005, 9.184473e-005, 9.144738e-005, 
    9.087517e-005, 8.996919e-005, 8.868173e-005, 8.707636e-005, 
    8.508953e-005, 8.272124e-005, 8.008274e-005, 7.72535e-005, 7.43448e-005, 
    7.146789e-005, 6.855917e-005, 6.572995e-005, 6.305968e-005, 6.050064e-005,
  7.742835e-005, 7.391567e-005, 7.094338e-005, 6.855918e-005, 6.647699e-005, 
    6.428357e-005, 6.207424e-005, 6.01033e-005, 5.83072e-005, 5.681312e-005, 
    5.557334e-005, 5.447661e-005, 5.36342e-005, 5.303021e-005, 5.258516e-005, 
    5.250567e-005, 5.223547e-005, 5.209243e-005, 5.180632e-005, 
    5.131359e-005, 5.07096e-005, 4.980361e-005, 4.883403e-005, 4.772141e-005, 
    4.665648e-005, 4.575048e-005, 4.497166e-005, 4.452662e-005, 
    4.451071e-005, 4.482859e-005, 4.560743e-005, 4.686312e-005, 
    4.889764e-005, 5.193349e-005, 5.585945e-005, 6.080263e-005, 
    6.687435e-005, 7.413817e-005, 8.18152e-005, 8.984195e-005, 9.753491e-005, 
    0.000104751, 0.0001112838, 0.0001193424, 0.0001249373, 0.0001283865, 
    0.0001374464, 0.0001447262, 0.0001526099, 0.0001582048, 0.0001659137, 
    0.0001746558, 0.0001778982, 0.0001838109, 0.0001795035, 0.0001894535, 
    0.0001867037, 0.0001806002, 0.0001728913, 0.0001637519, 0.000154104, 
    0.0001438679, 0.0001334569, 0.0001240155, 0.0001160046, 0.0001095513, 
    0.0001044014, 9.976016e-005, 9.565937e-005, 9.227381e-005, 9.163804e-005, 
    9.260763e-005, 9.437191e-005, 9.76939e-005, 0.0001032887, 0.000110648, 
    0.0001171331, 0.0001236976, 0.0001275917, 0.000132233, 0.0001354437, 
    0.0001349351, 0.0001362384, 0.0001333932, 0.0001321852, 0.0001296104, 
    0.0001265268, 0.0001228233, 0.0001185635, 0.0001135725, 0.0001081048, 
    0.0001026371, 9.712167e-005, 9.149502e-005, 8.613855e-005, 8.14815e-005,
  6.978307e-005, 6.401334e-005, 5.859332e-005, 5.315738e-005, 4.786449e-005, 
    4.322326e-005, 3.964697e-005, 3.745352e-005, 3.670648e-005, 
    3.716743e-005, 3.799394e-005, 3.974234e-005, 4.226957e-005, 
    4.543259e-005, 4.867509e-005, 5.212419e-005, 5.463556e-005, 
    5.541439e-005, 5.423819e-005, 5.110697e-005, 4.703796e-005, 4.30643e-005, 
    3.95993e-005, 3.743761e-005, 3.681774e-005, 3.781909e-005, 4.007613e-005, 
    4.287357e-005, 4.54167e-005, 4.729225e-005, 4.846846e-005, 4.962877e-005, 
    5.118643e-005, 5.380907e-005, 5.797342e-005, 6.431533e-005, 
    7.275536e-005, 8.380209e-005, 9.675615e-005, 0.000110791, 0.0001247624, 
    0.0001359523, 0.0001459341, 0.0001502257, 0.0001499397, 0.0001510204, 
    0.0001508296, 0.0001533091, 0.0001593809, 0.0001672646, 0.0001773894, 
    0.0001882135, 0.0001992285, 0.0002076845, 0.0002126753, 0.0002116897, 
    0.0002030273, 0.0001904706, 0.0001751641, 0.000160859, 0.0001508931, 
    0.0001431684, 0.0001400214, 0.0001363657, 0.0001348875, 0.0001349828, 
    0.0001336159, 0.0001333616, 0.0001327734, 0.0001321217, 0.0001312475, 
    0.0001315654, 0.0001307389, 0.0001293879, 0.0001304051, 0.0001338384, 
    0.0001343947, 0.0001366676, 0.0001396876, 0.0001400532, 0.0001402279, 
    0.0001401167, 0.0001409591, 0.0001405935, 0.0001400213, 0.0001407365, 
    0.0001420081, 0.0001430095, 0.0001421671, 0.0001389883, 0.0001331072, 
    0.0001229823, 0.0001098692, 9.726471e-005, 8.624981e-005, 7.715815e-005,
  7.062548e-005, 6.290071e-005, 5.70992e-005, 5.174277e-005, 4.705384e-005, 
    4.468556e-005, 4.478091e-005, 4.687901e-005, 5.042351e-005, 5.4572e-005, 
    5.800523e-005, 6.078677e-005, 6.402926e-005, 6.857511e-005, 
    7.528259e-005, 8.439019e-005, 9.384745e-005, 0.0001020967, 0.000104465, 
    9.980792e-005, 8.80936e-005, 7.164272e-005, 5.581175e-005, 4.352526e-005, 
    3.645217e-005, 3.580051e-005, 3.974236e-005, 4.497166e-005, 
    4.899298e-005, 5.107517e-005, 5.212423e-005, 5.22037e-005, 5.325275e-005, 
    5.663828e-005, 6.050068e-005, 6.382262e-005, 6.604788e-005, 6.82095e-005, 
    7.215134e-005, 7.990788e-005, 9.243281e-005, 0.0001072624, 0.0001243651, 
    0.0001409433, 0.0001569332, 0.000171588, 0.0001917738, 0.0001841444, 
    0.0001799166, 0.0001768172, 0.0001729548, 0.000170078, 0.0001683455, 
    0.000164674, 0.0001583319, 0.0001531187, 0.0001438364, 0.0001252712, 
    0.0001202959, 0.000122696, 0.0001275599, 0.0001314222, 0.0001383523, 
    0.0001461248, 0.0001506071, 0.0001551371, 0.0001596828, 0.0001641334, 
    0.0001720648, 0.0001771828, 0.0001795829, 0.0001815856, 0.0001823009, 
    0.0001822214, 0.0001851778, 0.00018877, 0.0001928866, 0.0001963993, 
    0.0001979094, 0.0001989106, 0.0002347687, 0.0002269964, 0.0002297142, 
    0.0002316219, 0.0002445759, 0.0002634746, 0.0002846144, 0.0002995552, 
    0.0003251615, 0.0002652543, 0.0002420803, 0.0002060314, 0.0001652302, 
    0.0001277507, 0.0001008569, 8.259405e-005,
  0.0001287204, 0.0001137794, 0.0001018266, 8.993741e-005, 7.91926e-005, 
    7.364538e-005, 7.617261e-005, 8.202184e-005, 9.182878e-005, 
    9.858399e-005, 9.852037e-005, 8.946049e-005, 7.685611e-005, 
    6.778035e-005, 6.595248e-005, 7.297788e-005, 8.578887e-005, 0.0001002688, 
    0.0001118718, 0.0001143197, 0.0001116017, 9.647006e-005, 7.485336e-005, 
    5.614545e-005, 4.506696e-005, 4.253976e-005, 4.68631e-005, 5.398388e-005, 
    5.794162e-005, 5.790981e-005, 5.512827e-005, 5.465143e-005, 
    6.032581e-005, 7.035525e-005, 8.222851e-005, 8.963537e-005, 
    9.054135e-005, 8.578887e-005, 8.280066e-005, 8.437422e-005, 
    9.197183e-005, 0.0001026372, 0.000112476, 0.0001204552, 0.0001276077, 
    0.0001344424, 0.0001420396, 0.0001367469, 0.0001215995, 0.0001041156, 
    8.671114e-005, 7.464713e-005, 7.026026e-005, 7.469486e-005, 
    8.075067e-005, 8.143391e-005, 8.321414e-005, 9.18447e-005, 0.0001083913, 
    0.0001315179, 0.0001594446, 0.0001814427, 0.000199356, 0.0002085272, 
    0.0002145988, 0.0002248507, 0.0002445284, 0.0002670668, 0.0002889377, 
    0.0002930069, 0.000367457, 0.0003914259, 0.0003804904, 0.000358715, 
    0.0003372891, 0.0003015262, 0.0002952003, 0.0002759201, 0.0002590559, 
    0.0002435427, 0.0002459112, 0.0002225939, 0.0002081774, 0.0002065244, 
    0.0002190175, 0.000240348, 0.0002691331, 0.0002978386, 0.0003238901, 
    0.0003426296, 0.0003603997, 0.000289303, 0.0002577046, 0.0002201458, 
    0.000182587, 0.0001514496,
  0.0003391645, 0.0003187081, 0.0002588648, 0.0002183654, 0.0001836836, 
    0.000166136, 0.0001647373, 0.0001867036, 0.0002080977, 0.0002213378, 
    0.0002237538, 0.0002109111, 0.0001856069, 0.0001559955, 0.0001333774, 
    0.0001259705, 0.0001298806, 0.0001392903, 0.0001478415, 0.0001499713, 
    0.0001543742, 0.0001522283, 0.0001409273, 0.0001216949, 0.0001056255, 
    9.953789e-005, 0.0001073898, 0.0001250328, 0.0001403234, 0.0001421989, 
    0.0001289269, 0.0001118403, 0.0001028599, 0.0001001896, 0.0001020811, 
    0.0001044812, 0.0001003008, 9.494438e-005, 9.885448e-005, 0.0001110455, 
    0.0001253347, 0.0001362861, 0.0001302621, 0.0001129052, 9.200384e-005, 
    6.477651e-005, 4.117307e-005, 1.53603e-005, -4.412839e-006, 
    -1.661992e-005, -1.847977e-005, -1.42674e-005, -3.633788e-006, 
    4.138798e-006, 9.479467e-006, 1.626625e-005, 3.348035e-005, 
    5.223579e-005, 7.577566e-005, 9.494461e-005, 0.0001159729, 0.0001389247, 
    0.0001745762, 0.0002073827, 0.0002361361, 0.0002586904, 0.0002819281, 
    0.0003125572, 0.0003432338, 0.0003668212, 0.0003943983, 0.0004132332, 
    0.0004084331, 0.0003976407, 0.0003760718, 0.0003467305, 0.0003172143, 
    0.0002801323, 0.0003223481, 0.0003274184, 0.0003362877, 0.0003113174, 
    0.0002825165, 0.0002635862, 0.000265239, 0.000284519, 0.0003204409, 
    0.0003448231, 0.0003592236, 0.0003685697, 0.0003754839, 0.0003795048, 
    0.000389089, 0.0003916005, 0.0003809988, 0.0003629907,
  0.0004571658, 0.0004520479, 0.0004477407, 0.000438299, 0.0004272998, 
    0.0004187329, 0.0004155221, 0.0004108651, 0.0004033153, 0.0003903452, 
    0.0003865304, 0.0003939375, 0.0003920459, 0.000377121, 0.0003473505, 
    0.0003270371, 0.0003353023, 0.0003545982, 0.0003746731, 0.0003697774, 
    0.0003533587, 0.0003395145, 0.0003250819, 0.0003119371, 0.0003005246, 
    0.0002817534, 0.0002676073, 0.0002558134, 0.0002482951, 0.0002450051, 
    0.0002488676, 0.000255591, 0.0002494082, 0.0002870464, 0.0002849323, 
    0.0002784792, 0.0002923072, 0.0003008588, 0.0003075502, 0.000303831, 
    0.0002959156, 0.0002829772, 0.0002663357, 0.0002370896, 0.0001878166, 
    0.0001411019, 9.594555e-005, 7.081614e-005, 4.438334e-005, 1.392933e-005, 
    -8.92696e-006, -1.812982e-005, -1.501455e-005, -1.981482e-005, 
    -1.895661e-005, -7.067341e-006, 2.103415e-005, 4.724436e-005, 
    7.032324e-005, 7.924018e-005, 9.567523e-005, 0.0001276233, 0.0001765946, 
    0.000219462, 0.0002570208, 0.0002884921, 0.0003185647, 0.0003584442, 
    0.0003905194, 0.0004347542, 0.0004707235, 0.0005001444, 0.0005171993, 
    0.0005103645, 0.0004928964, 0.0004709777, 0.0004508235, 0.0004390457, 
    0.0004297472, 0.000426457, 0.000396162, 0.000367234, 0.0003418026, 
    0.0003252244, 0.0003327427, 0.0003571732, 0.00039141, 0.0004188281, 
    0.0004280945, 0.0004187645, 0.0004039984, 0.0003963055, 0.0004117868, 
    0.0004411126, 0.000463333, 0.0004639053,
  0.0004144572, 0.0003947001, 0.0003886444, 0.0003898842, 0.000395797, 
    0.0003959236, 0.0003926652, 0.0003855603, 0.0003677902, 0.0003603515, 
    0.0003742434, 0.0004230556, 0.0004799105, 0.0005043729, 0.0004923719, 
    0.0004629828, 0.000457976, 0.0004824696, 0.0004734413, 0.000447724, 
    0.0004152039, 0.0003838597, 0.0003693639, 0.0003575541, 0.0003481444, 
    0.0003303108, 0.0002942937, 0.0002408244, 0.0001950322, 0.0001755932, 
    0.0001744009, 0.0001746709, 0.0001910741, 0.0002215917, 0.0002469276, 
    0.0002969955, 0.0003048473, 0.0003088848, 0.000320758, 0.0003106806, 
    0.0002935147, 0.0002900497, 0.0003052766, 0.0003204083, 0.0003092501, 
    0.0002599135, 0.0002075408, 0.0001555975, 5.883118e-005, -6.147474e-005, 
    -0.0001549984, -0.0001878524, -0.0001755182, -0.0001353528, 
    -7.891119e-005, -2.264418e-005, 4.312955e-006, 1.245085e-005, 
    1.032092e-005, 2.990314e-005, 7.234165e-005, 0.0001188968, 0.0001600955, 
    0.0002058242, 0.0002699271, 0.0003362552, 0.00039942, 0.0004722809, 
    0.000551722, 0.000633579, 0.0007041828, 0.0007536942, 0.000781192, 
    0.0007944002, 0.0008087533, 0.0008163189, 0.0007800316, 0.0006833768, 
    0.0005564268, 0.0004283164, 0.0003486688, 0.0003022407, 0.0002614711, 
    0.0002639031, 0.0002741392, 0.0002832629, 0.000311269, 0.0003489074, 
    0.0003775018, 0.0003930307, 0.0003983874, 0.0004000878, 0.0004067319, 
    0.0004206556, 0.000433197, 0.0004290484,
  0.0003223792, 0.0003051972, 0.0002877924, 0.0002839779, 0.0002994749, 
    0.0003082331, 0.0003098859, 0.0003211552, 0.0003268772, 0.0003226493, 
    0.0003189777, 0.0003520227, 0.0003941432, 0.0004207029, 0.0004436707, 
    0.0004755233, 0.0005099191, 0.0005171353, 0.0004996513, 0.0004869041, 
    0.0004627283, 0.0004237229, 0.0003918861, 0.0003674722, 0.0003334894, 
    0.000295104, 0.000239314, 0.000183715, 0.0001612082, 0.0001725887, 
    0.0001904382, 0.0001983061, 0.0002096391, 0.0002125476, 0.0002168396, 
    0.0002416824, 0.0003147973, 0.0003842884, 0.0004254079, 0.0004316864, 
    0.0004355328, 0.0004979346, 0.0006129004, 0.0006773369, 0.0006507612, 
    0.0006075278, 0.0005101576, 0.0003366689, 0.0001561698, -6.342959e-005, 
    -0.0001882501, -0.000188075, -0.0001735948, -0.0001841486, -0.000211122, 
    -0.0002000113, -0.0001912541, -0.0001947191, -0.0001134179, 
    4.125154e-005, 0.0001782314, 0.0002693231, 0.000353565, 0.0004546861, 
    0.0005537886, 0.0006172559, 0.0006827409, 0.0007459535, 0.0007817643, 
    0.0008131401, 0.0008497611, 0.0008914527, 0.000924068, 0.0009322856, 
    0.0009108912, 0.0008645901, 0.0007704627, 0.0007118913, 0.0006711222, 
    0.0006401436, 0.000583082, 0.0004872533, 0.0003692205, 0.0002935305, 
    0.0002682898, 0.0002538734, 0.0002515528, 0.0002835963, 0.0002848201, 
    0.0002975517, 0.000320917, 0.0003476199, 0.0003549312, 0.0003390207, 
    0.0003174995, 0.0003219023,
  0.000336573, 0.0003585711, 0.0004175401, 0.0004896536, 0.0005127962, 
    0.0005165313, 0.000529072, 0.0005545989, 0.0005730689, 0.000569683, 
    0.0005486228, 0.0005402304, 0.0005384504, 0.0005530573, 0.0005914746, 
    0.0006435451, 0.0006948214, 0.0007504681, 0.0007417419, 0.0006023622, 
    0.0004845196, 0.0004385686, 0.000415124, 0.0004221334, 0.0004328466, 
    0.0004294452, 0.000429827, 0.0004402532, 0.0004642699, 0.0004880168, 
    0.0004786863, 0.0004461664, 0.0004281262, 0.0004009781, 0.0003744815, 
    0.0003926968, 0.0004632049, 0.0005534389, 0.00061282, 0.000617207, 
    0.0006254409, 0.000686158, 0.0007760259, 0.0007861028, 0.0007530111, 
    0.0007406455, 0.0007124157, 0.0006115008, 0.0004944853, 0.000334077, 
    0.000221909, 0.0001767208, 0.0001290371, 7.216632e-005, 2.834573e-005, 
    1.947582e-005, 2.637412e-005, 4.166458e-005, 0.0001089303, 0.0002023592, 
    0.0002928465, 0.0003560116, 0.0004288885, 0.0005142423, 0.0005705245, 
    0.0005943668, 0.0006432896, 0.000706932, 0.0007504513, 0.000787613, 
    0.0008270792, 0.0008474085, 0.0008517792, 0.0008368068, 0.0007792525, 
    0.0006770189, 0.0006763195, 0.0008165091, 0.0008813115, 0.00073737, 
    0.0007226197, 0.0006519365, 0.0005355575, 0.000415442, 0.0003446797, 
    0.0003477631, 0.0003855922, 0.0004037751, 0.0004030124, 0.0004013912, 
    0.000397624, 0.000410324, 0.0004064932, 0.0003803466, 0.0003592863, 
    0.0003451877,
  0.0006036176, 0.0006496962, 0.0007055178, 0.0007462557, 0.0007658377, 
    0.0007729265, 0.0007927474, 0.0008113594, 0.0008241073, 0.0008408441, 
    0.0008409875, 0.0008286531, 0.0008276836, 0.0008215802, 0.0008291141, 
    0.000854434, 0.0008982234, 0.0009701466, 0.001009041, 0.0009374353, 
    0.0008495864, 0.0008402723, 0.0008415589, 0.0008033807, 0.0007643439, 
    0.0007550297, 0.0007618004, 0.0007475107, 0.0007430604, 0.0007505468, 
    0.000748687, 0.0007204269, 0.0006734589, 0.0006164452, 0.0005921423, 
    0.0006198464, 0.0006583747, 0.0006791493, 0.0007038177, 0.0007600207, 
    0.0008362038, 0.0009028492, 0.0009140549, 0.0009028655, 0.0009320001, 
    0.000950072, 0.0009052497, 0.0008247914, 0.0007656477, 0.0007101116, 
    0.0006344379, 0.0005225241, 0.00042002, 0.0003737193, 0.0003704447, 
    0.0003700475, 0.0003819684, 0.0004082583, 0.0004513958, 0.000501893, 
    0.0005302648, 0.0005610203, 0.0006084819, 0.0006308611, 0.0006352803, 
    0.000660012, 0.0006839493, 0.0006817877, 0.0006881137, 0.0007161996, 
    0.0007401528, 0.0007353048, 0.0007139901, 0.0006851573, 0.0006505069, 
    0.0006550848, 0.0007365448, 0.0007802704, 0.0007651863, 0.0007347167, 
    0.000674508, 0.0006146175, 0.0005511651, 0.000466702, 0.0004384415, 
    0.0005065026, 0.0005827006, 0.0006253454, 0.0006344211, 0.0006640493, 
    0.0006564828, 0.0006117877, 0.000594208, 0.0005802691, 0.0005626576, 
    0.0005689999,
  0.0007683807, 0.0008197832, 0.0008523199, 0.0008903076, 0.0009292495, 
    0.0009755827, 0.001056867, 0.001125357, 0.001154396, 0.001186233, 
    0.001223569, 0.001243231, 0.00122891, 0.001177094, 0.001129219, 
    0.00111501, 0.001138057, 0.001163568, 0.001187536, 0.001261685, 
    0.001428307, 0.001567862, 0.001553287, 0.001415243, 0.001308066, 
    0.00123964, 0.001153348, 0.001037556, 0.0009417115, 0.0008900226, 
    0.00086537, 0.0008024913, 0.0007462879, 0.0007305681, 0.0007471945, 
    0.0007737698, 0.0007735309, 0.0007466055, 0.0007434911, 0.0007968172, 
    0.0009279316, 0.001045457, 0.001087466, 0.00107332, 0.001147564, 
    0.00121324, 0.00110406, 0.001075624, 0.001041656, 0.001021502, 
    0.001000665, 0.0009358628, 0.0008384129, 0.0007715919, 0.0007386748, 
    0.0007245285, 0.0007229871, 0.0007316815, 0.0007308703, 0.0007379758, 
    0.0007286612, 0.0007220171, 0.000736529, 0.0007012426, 0.000686985, 
    0.000690069, 0.000656595, 0.0006288271, 0.0006314656, 0.0006304323, 
    0.0006421786, 0.000658677, 0.0006521125, 0.0006276192, 0.0006159046, 
    0.0006375373, 0.0007248144, 0.0007925094, 0.0006710114, 0.0007383088, 
    0.0006633978, 0.0006380775, 0.0006669583, 0.0006782273, 0.0006569922, 
    0.0006653843, 0.0006925166, 0.0006950917, 0.0007099686, 0.0007360829, 
    0.0007154993, 0.0006782585, 0.0006717574, 0.0006828359, 0.000685649, 
    0.0007183282,
  0.0009347182, 0.001009979, 0.001075464, 0.0011286, 0.00119148, 0.001309958, 
    0.001533197, 0.001747662, 0.0018735, 0.001945947, 0.002002929, 
    0.001996142, 0.001869845, 0.001732834, 0.001642075, 0.001598699, 
    0.001576239, 0.001552239, 0.001575095, 0.001647335, 0.001669015, 
    0.001625798, 0.001479647, 0.001325532, 0.00122883, 0.001127392, 
    0.001010932, 0.0009350036, 0.0008796589, 0.0008164463, 0.0007914766, 
    0.0007887743, 0.0008071014, 0.0008196733, 0.0007994715, 0.000788887, 
    0.0007944326, 0.0008054785, 0.0008683577, 0.0009321431, 0.001127677, 
    0.001266611, 0.001328854, 0.001313405, 0.001383548, 0.001469474, 
    0.001420233, 0.001401238, 0.001455391, 0.00151703, 0.001585312, 
    0.001523658, 0.001365285, 0.001243962, 0.001161247, 0.001069646, 
    0.001019308, 0.0009504049, 0.0008703452, 0.0008494765, 0.0008384446, 
    0.0008380637, 0.0008218032, 0.0007857229, 0.0007640268, 0.0007511522, 
    0.0007209829, 0.0007251804, 0.0007270416, 0.0007073795, 0.0007079039, 
    0.0007379283, 0.0007546176, 0.0007212395, 0.0006619045, 0.0006489656, 
    0.0007076645, 0.0007744213, 0.0005645812, 0.0008126795, 0.0006952505, 
    0.0006796098, 0.0007661404, 0.0008585192, 0.0008563418, 0.0007853252, 
    0.0007721009, 0.000798041, 0.000810375, 0.0008364101, 0.0008370937, 
    0.0008187196, 0.0007977863, 0.0007794914, 0.0008118851, 0.0008740807,
  0.001098703, 0.001116551, 0.001108842, 0.00114052, 0.001281854, 0.00152396, 
    0.001689296, 0.001912504, 0.002100742, 0.002155023, 0.0019788, 
    0.001797633, 0.00163554, 0.001514615, 0.001425017, 0.00135942, 
    0.001356368, 0.001354349, 0.001301786, 0.001267455, 0.00123104, 
    0.001193512, 0.001144731, 0.001054276, 0.0009695739, 0.0009093331, 
    0.0008762097, 0.0008575171, 0.000835917, 0.0008716797, 0.0009476719, 
    0.0009436188, 0.000925133, 0.0008698674, 0.0008376334, 0.0008969363, 
    0.0009575412, 0.001001824, 0.001022472, 0.001537391, 0.001386775, 
    0.001743354, 0.001846175, 0.001786364, 0.001756911, 0.001746723, 
    0.00172978, 0.001711453, 0.001706145, 0.001638274, 0.001494476, 
    0.001386235, 0.001301612, 0.00120777, 0.001120477, 0.001054896, 
    0.001010773, 0.000940185, 0.0009075059, 0.0009236699, 0.0009475918, 
    0.0009410903, 0.0009004008, 0.00085124, 0.0008722674, 0.0008881781, 
    0.0008727293, 0.000885237, 0.0008792607, 0.0008431971, 0.0008561509, 
    0.0008593937, 0.0007886468, 0.0007283902, 0.0006523663, 0.0006585969, 
    0.0007365765, 0.0007827817, 0.000954729, 0.00118237, 0.0008558007, 
    0.0008490141, 0.001029355, 0.001139995, 0.001149135, 0.001046409, 
    0.001009041, 0.0009878371, 0.0009696539, 0.001006831, 0.001025984, 
    0.001050303, 0.001030132, 0.0009866925, 0.001015732, 0.00107014,
  0.001151661, 0.001157734, 0.001129172, 0.001236348, 0.001487593, 
    0.00170136, 0.001946691, 0.002089361, 0.002216946, 0.002058334, 
    0.001656153, 0.001480677, 0.001449954, 0.001416098, 0.001394115, 
    0.00131868, 0.001294537, 0.001285351, 0.001181798, 0.001109128, 
    0.001043945, 0.0009973738, 0.001006354, 0.0009871852, 0.000972514, 
    0.0009875344, 0.001020183, 0.001054863, 0.001092932, 0.001218149, 
    0.001173533, 0.001180225, 0.001182624, 0.00112639, 0.001112101, 
    0.001129649, 0.001061094, 0.001703315, 0.001856968, 0.001881192, 
    0.002131323, 0.002421828, 0.002541467, 0.002249277, 0.002055665, 
    0.001941193, 0.001805788, 0.001679043, 0.001568513, 0.001420153, 
    0.001254802, 0.001195675, 0.001155429, 0.001067644, 0.001038207, 
    0.001044421, 0.001033041, 0.001006115, 0.001017417, 0.001083602, 
    0.001105504, 0.001088115, 0.001042927, 0.001003763, 0.0009725466, 
    0.0009455094, 0.0009161048, 0.0009041512, 0.0008525737, 0.0008149827, 
    0.000789552, 0.0007151496, 0.0006553698, 0.0006845044, 0.0006172387, 
    0.000704214, 0.0008035069, 0.001625749, 0.001335643, 0.001345576, 
    0.001184626, 0.001234664, 0.001468218, 0.001744082, 0.001698767, 
    0.001472779, 0.001424665, 0.001402304, 0.001329141, 0.001284763, 
    0.001205401, 0.0011622, 0.001133923, 0.001084253, 0.001090086, 0.001110718,
  0.001267533, 0.001251051, 0.001226987, 0.001374504, 0.00155238, 0.00166935, 
    0.002191311, 0.002891958, 0.002926782, 0.002392406, 0.002109864, 
    0.0020889, 0.002077407, 0.0019616, 0.001860781, 0.001793086, 0.001739171, 
    0.001670188, 0.001543286, 0.00147974, 0.001446981, 0.001384913, 
    0.001369242, 0.001372547, 0.001422157, 0.001415942, 0.001427162, 
    0.001504267, 0.001479663, 0.001427432, 0.001392462, 0.001859445, 
    0.00158722, 0.001367988, 0.001163808, 0.001238337, 0.001607233, 
    0.001767004, 0.001950299, 0.002124617, 0.002432111, 0.002183774, 
    0.001876707, 0.001726456, 0.00179822, 0.001797044, 0.001679312, 
    0.001484763, 0.001375853, 0.001357176, 0.00131709, 0.001263765, 
    0.001207403, 0.001131553, 0.001119205, 0.00109541, 0.001098542, 
    0.001146924, 0.001209326, 0.001261524, 0.001216701, 0.001168191, 
    0.001109475, 0.001031831, 0.0009853235, 0.0009525809, 0.00091046, 
    0.0008104825, 0.0007936824, 0.0007355101, 0.0006459914, 0.0007133214, 
    0.0006874604, 0.0006824229, 0.0006065266, 0.0006963303, 0.0008323397, 
    0.0008943602, 0.00142551, 0.001891949, 0.001736787, 0.00207097, 
    0.002104429, 0.002046334, 0.002025114, 0.001752475, 0.001675561, 
    0.001599267, 0.001480026, 0.001449063, 0.001372483, 0.001343158, 
    0.00134025, 0.001318919, 0.001310114, 0.001255786,
  0.001297207, 0.001280962, 0.001337547, 0.00147993, 0.001821314, 
    0.002306355, 0.002800945, 0.003089018, 0.002903878, 0.002505816, 
    0.002507039, 0.002537811, 0.002584811, 0.002463043, 0.002329784, 
    0.002249784, 0.002172775, 0.002032346, 0.00194197, 0.001854836, 
    0.001740935, 0.001743781, 0.00172075, 0.001692028, 0.001712849, 
    0.001658125, 0.001591876, 0.001563092, 0.001558243, 0.001662781, 
    0.00175772, 0.002404454, 0.002208937, 0.001140108, 0.0009582727, 
    0.001418422, 0.00164023, 0.001656314, 0.002190769, 0.002239327, 
    0.002488934, 0.001784169, 0.0016017, 0.001629991, 0.001758404, 
    0.001811952, 0.001807201, 0.001788221, 0.001727489, 0.001710053, 
    0.001675544, 0.001536452, 0.001402635, 0.001305329, 0.001259663, 
    0.001231546, 0.001280231, 0.001337198, 0.001331174, 0.001284825, 
    0.001211932, 0.00117048, 0.00108263, 0.001017049, 0.0009937789, 
    0.000977519, 0.001014872, 0.000936877, 0.0009306148, 0.0008624103, 
    0.0008019153, 0.0008624736, 0.0007004933, 0.000720012, 0.0007049926, 
    0.000774961, 0.001165617, 0.0007714164, 0.002013164, 0.002555946, 
    0.002477237, 0.002716832, 0.002948813, 0.002734761, 0.002396253, 
    0.002128733, 0.002058065, 0.001974809, 0.001839085, 0.001752888, 
    0.001689977, 0.001691837, 0.001664562, 0.001547704, 0.001440497, 
    0.001303867,
  0.001435903, 0.001431548, 0.001616258, 0.001945593, 0.002117019, 
    0.003146556, 0.003090082, 0.003089034, 0.003093867, 0.00275892, 
    0.002916532, 0.002875891, 0.003104455, 0.002597416, 0.00238392, 
    0.002330451, 0.002233779, 0.002141321, 0.002034349, 0.001965622, 
    0.001856489, 0.001883351, 0.001902567, 0.001877057, 0.00182427, 
    0.001780481, 0.001765191, 0.001797647, 0.001857602, 0.002007154, 
    0.002130321, 0.00249259, 0.001988924, 0.001054324, 0.001087051, 
    0.001727365, 0.001673594, 0.002011828, 0.002458972, 0.002482068, 
    0.002378913, 0.001901598, 0.00200771, 0.002156578, 0.002173379, 
    0.002170295, 0.002112917, 0.002093493, 0.002041645, 0.001908323, 
    0.001791815, 0.001568083, 0.001429356, 0.001333924, 0.001342968, 
    0.001424237, 0.001475339, 0.001528474, 0.001483398, 0.001436174, 
    0.001396358, 0.001379669, 0.001354349, 0.001272762, 0.001240098, 
    0.001238684, 0.001251526, 0.00119208, 0.001115579, 0.001049935, 
    0.001013441, 0.0009764861, 0.0008802125, 0.000882946, 0.0008329591, 
    0.001147003, 0.00191603, 0.001093091, 0.001833619, 0.003085076, 
    0.003042561, 0.003067611, 0.003275194, 0.003036044, 0.002928199, 
    0.002482038, 0.002526716, 0.002359633, 0.002163573, 0.0020601, 
    0.001961377, 0.001800301, 0.001661177, 0.001512705, 0.001428242, 
    0.001348339,
  0.001747691, 0.00175532, 0.001956783, 0.002263152, 0.002609526, 
    0.003458821, 0.003400763, 0.003318458, 0.003312879, 0.002726051, 
    0.003105598, 0.003227685, 0.002927134, 0.002649487, 0.002464918, 
    0.002410481, 0.002270164, 0.002286057, 0.002185667, 0.002130927, 
    0.002153686, 0.002177688, 0.002165561, 0.002165512, 0.002111693, 
    0.002100105, 0.002091237, 0.002154037, 0.002271656, 0.002444494, 
    0.002595684, 0.00274147, 0.002430649, 0.0007538055, 0.001320748, 
    0.001600637, 0.001885595, 0.002635339, 0.002967458, 0.002275773, 
    0.002124362, 0.002314794, 0.002410845, 0.002471816, 0.002540276, 
    0.002592633, 0.002587721, 0.002463281, 0.0023953, 0.002230171, 
    0.002099263, 0.00194631, 0.001876501, 0.001880554, 0.001899628, 
    0.001999192, 0.002045127, 0.002073053, 0.002103904, 0.00215197, 
    0.002157183, 0.002090793, 0.002039978, 0.001928619, 0.001793626, 
    0.001716029, 0.00157274, 0.00147564, 0.001404051, 0.001356224, 
    0.001274748, 0.001252861, 0.001275845, 0.001207847, 0.001286017, 
    0.001587013, 0.002282177, 0.001661911, 0.002308962, 0.003272236, 
    0.003306219, 0.003258059, 0.003391191, 0.003336278, 0.003398933, 
    0.00293079, 0.002502479, 0.002367883, 0.002174572, 0.002051738, 
    0.001950602, 0.001755066, 0.001674067, 0.001592925, 0.001581338, 
    0.001613811,
  0.002150125, 0.002168277, 0.002214165, 0.002371871, 0.002805143, 
    0.003198151, 0.003306968, 0.003077482, 0.003306983, 0.002677381, 
    0.002547491, 0.003089862, 0.003052367, 0.002691098, 0.002540229, 
    0.002622673, 0.0024962, 0.002569031, 0.002574768, 0.002573702, 
    0.00258556, 0.00259826, 0.002577976, 0.00260646, 0.002574067, 
    0.002588324, 0.002627362, 0.00271127, 0.002808116, 0.002886271, 
    0.003032165, 0.003449382, 0.003624031, 0.003628625, 0.003666281, 
    0.002883246, 0.002535379, 0.002588263, 0.002849998, 0.002366357, 
    0.002536494, 0.002656434, 0.002715338, 0.002759112, 0.002896966, 
    0.00298316, 0.003045198, 0.002945619, 0.002829717, 0.002660105, 
    0.00262199, 0.002634516, 0.002703609, 0.002751261, 0.002793333, 
    0.002902402, 0.00297555, 0.002986517, 0.003004158, 0.002974721, 
    0.002882821, 0.002779951, 0.002633115, 0.002500365, 0.002320278, 
    0.002219298, 0.002070542, 0.001993787, 0.001928413, 0.001854375, 
    0.001823635, 0.00184673, 0.001801017, 0.001730413, 0.00176384, 
    0.001953382, 0.002258449, 0.002402565, 0.002565372, 0.003652087, 
    0.003473446, 0.003241941, 0.0034013, 0.002969764, 0.003122257, 
    0.002665397, 0.002530772, 0.002361063, 0.002240789, 0.0021582, 
    0.00208906, 0.002013464, 0.002038372, 0.00200523, 0.002099501, 0.002126014,
  0.002434766, 0.002501364, 0.002624356, 0.002876954, 0.003296953, 
    0.003166793, 0.00320103, 0.003017542, 0.002904166, 0.002328415, 
    0.002320706, 0.002867799, 0.002839936, 0.0026547, 0.002877846, 
    0.002931982, 0.002988297, 0.002981208, 0.002978999, 0.002973624, 
    0.002987532, 0.002990203, 0.002988122, 0.002986787, 0.002983337, 
    0.002958097, 0.003043482, 0.003180938, 0.003273541, 0.003315471, 
    0.003283283, 0.003513565, 0.003805708, 0.003625907, 0.003540093, 
    0.00361618, 0.003160482, 0.00281382, 0.00271046, 0.002636706, 
    0.002839539, 0.002905374, 0.002942266, 0.002978157, 0.003126627, 
    0.003206242, 0.003255961, 0.003201062, 0.003139867, 0.003150851, 
    0.003167206, 0.003287226, 0.003329329, 0.003350344, 0.003500579, 
    0.003556481, 0.003628133, 0.003566382, 0.00346658, 0.003312785, 
    0.003150182, 0.003052112, 0.002904929, 0.00282819, 0.00269668, 
    0.002568727, 0.002482419, 0.002416264, 0.002403088, 0.002376655, 
    0.002354785, 0.002310996, 0.002260084, 0.002251375, 0.00225743, 
    0.002782857, 0.003226076, 0.002642286, 0.002800452, 0.003766257, 
    0.003415924, 0.002994051, 0.003233805, 0.003077308, 0.002929993, 
    0.002354626, 0.002684487, 0.002579123, 0.002557427, 0.002493832, 
    0.002464713, 0.002424325, 0.002436038, 0.002441888, 0.002484803, 
    0.002486137,
  0.002804999, 0.002830654, 0.002963819, 0.002883632, 0.002879704, 
    0.00322589, 0.003238399, 0.00320413, 0.002816047, 0.002534823, 
    0.002356232, 0.002896395, 0.002940534, 0.003158018, 0.003248347, 
    0.003281964, 0.003402047, 0.003370911, 0.003316265, 0.003188394, 
    0.003196498, 0.00320467, 0.003223123, 0.003200727, 0.003207339, 
    0.00319572, 0.003249127, 0.003318347, 0.003262844, 0.003306538, 
    0.003445202, 0.003355842, 0.003355304, 0.003340553, 0.003346767, 
    0.003166094, 0.003089037, 0.002927404, 0.002544012, 0.0026832, 
    0.002935225, 0.003055738, 0.003128838, 0.003148593, 0.003156191, 
    0.003132906, 0.003062032, 0.003071267, 0.003129344, 0.003320573, 
    0.003347147, 0.003426621, 0.003553746, 0.003675435, 0.003783185, 
    0.003761061, 0.003769657, 0.003675928, 0.003570547, 0.003420867, 
    0.003314866, 0.003225109, 0.003168762, 0.00307419, 0.003002046, 
    0.002878895, 0.002834264, 0.002821578, 0.002823675, 0.002816412, 
    0.002794797, 0.002805952, 0.002835182, 0.002881788, 0.002938132, 
    0.003247711, 0.002616789, 0.002418823, 0.002974564, 0.003361406, 
    0.002991108, 0.002817415, 0.002790599, 0.003524326, 0.002851589, 
    0.002742995, 0.002560508, 0.002882835, 0.002958924, 0.00280791, 
    0.00280834, 0.002783876, 0.00275708, 0.0027868, 0.002768665, 0.002774926,
  0.003197836, 0.003137086, 0.003263829, 0.003141709, 0.003137676, 
    0.00318566, 0.003152933, 0.00297164, 0.002841908, 0.002700841, 
    0.003005318, 0.002995307, 0.003166905, 0.003378015, 0.003483666, 
    0.003544003, 0.003522117, 0.00350506, 0.003513502, 0.003408533, 
    0.00336986, 0.003372803, 0.003444821, 0.003438719, 0.003414938, 
    0.003398949, 0.003452146, 0.003468998, 0.003443945, 0.003319651, 
    0.003320843, 0.003338391, 0.003357369, 0.003205338, 0.003141187, 
    0.003169511, 0.00304763, 0.002812617, 0.002579486, 0.002689416, 
    0.003031245, 0.003091771, 0.003155667, 0.003173739, 0.003197184, 
    0.003340075, 0.003417816, 0.00366752, 0.003915697, 0.004127858, 
    0.004228789, 0.004248131, 0.004292464, 0.004344167, 0.004335998, 
    0.004258161, 0.004192088, 0.004068237, 0.003982455, 0.003806723, 
    0.003739968, 0.003626939, 0.003561391, 0.003443899, 0.00340626, 
    0.003306713, 0.003260015, 0.003257917, 0.003240148, 0.003263846, 
    0.003283825, 0.003280138, 0.003239336, 0.003211569, 0.003352694, 
    0.003418945, 0.002396318, 0.003209898, 0.003689375, 0.003123719, 
    0.002415916, 0.00180221, 0.001997394, 0.002707596, 0.003103534, 
    0.002951184, 0.003189759, 0.003250096, 0.003243644, 0.003204953, 
    0.003198897, 0.003179874, 0.003098002, 0.003084188, 0.003088146, 
    0.003115771,
  0.003438238, 0.003405338, 0.003362359, 0.003101721, 0.003157875, 
    0.002890211, 0.003032451, 0.002755092, 0.002690366, 0.002733886, 
    0.002845451, 0.00335988, 0.003148403, 0.003303375, 0.003416225, 
    0.003416482, 0.00329894, 0.003251621, 0.003252847, 0.003298828, 
    0.003384104, 0.003401667, 0.003399808, 0.003447397, 0.003473798, 
    0.003458712, 0.00355063, 0.003144443, 0.003260316, 0.003482936, 
    0.003085872, 0.002858517, 0.00281789, 0.003119094, 0.003223171, 
    0.003219912, 0.002875715, 0.00301268, 0.003107838, 0.003160339, 
    0.003166554, 0.003163328, 0.003186248, 0.003285239, 0.003431089, 
    0.003772678, 0.004192915, 0.004607175, 0.004787944, 0.004720423, 
    0.004657354, 0.004533043, 0.004391404, 0.004308483, 0.004186809, 
    0.004073957, 0.003964938, 0.003877884, 0.003834493, 0.003768481, 
    0.00381119, 0.003796043, 0.003787477, 0.003758978, 0.003727823, 
    0.003661146, 0.003616609, 0.00358358, 0.003554875, 0.003501248, 
    0.003515011, 0.003409917, 0.003400076, 0.003321512, 0.003170302, 
    0.003420994, 0.002894233, 0.003497733, 0.003514852, 0.002443431, 
    0.001663737, 0.001450653, 0.00187828, 0.002419109, 0.002690354, 
    0.003293505, 0.0032802, 0.003356177, 0.003372468, 0.003426015, 
    0.00333265, 0.003362151, 0.003360085, 0.003402047, 0.003351804, 
    0.003343984,
  0.003171671, 0.003401777, 0.003366111, 0.003036585, 0.00319054, 
    0.003290581, 0.003108429, 0.002813439, 0.002855242, 0.003036934, 
    0.002928168, 0.003211122, 0.003410265, 0.003277848, 0.003385598, 
    0.00349538, 0.00345787, 0.003348324, 0.003339695, 0.003257392, 
    0.00324377, 0.003220532, 0.003121635, 0.00320629, 0.003305648, 0.0033643, 
    0.00347076, 0.00286041, 0.003180303, 0.003265705, 0.003180429, 
    0.002847121, 0.00267333, 0.00296169, 0.002973834, 0.003001092, 
    0.002955221, 0.003034057, 0.003203971, 0.003248585, 0.003232628, 
    0.003269853, 0.003208168, 0.003303835, 0.003429897, 0.003719226, 
    0.00416211, 0.004538748, 0.004764689, 0.004747493, 0.004727624, 
    0.004694181, 0.004592583, 0.004483005, 0.004337078, 0.004206792, 
    0.004113283, 0.004036702, 0.003969086, 0.003952747, 0.003898244, 
    0.003891204, 0.003852502, 0.003806151, 0.003780244, 0.003739027, 
    0.003697256, 0.003609629, 0.003594544, 0.003511019, 0.003505282, 
    0.003304901, 0.003156079, 0.003041655, 0.002803586, 0.003132856, 
    0.003050175, 0.002735447, 0.002840254, 0.001774728, 0.002020014, 
    0.001937217, 0.002308533, 0.00311698, 0.003033563, 0.003084714, 
    0.003034376, 0.003129536, 0.003153395, 0.003135623, 0.003217608, 
    0.003305601, 0.0032205, 0.003251368, 0.003230514, 0.003217211,
  0.00323269, 0.003487688, 0.002567137, 0.002493514, 0.002664633, 
    0.003159544, 0.003381035, 0.002877639, 0.002949166, 0.003175043, 
    0.002809068, 0.003148783, 0.003295492, 0.003339376, 0.003313515, 
    0.003532654, 0.003648637, 0.003635539, 0.003649527, 0.003517918, 
    0.003422918, 0.003432916, 0.003257662, 0.003149658, 0.003076496, 
    0.003099939, 0.002901861, 0.00255703, 0.003073586, 0.003055213, 
    0.003096538, 0.003143346, 0.003104661, 0.003123004, 0.003112799, 
    0.0030853, 0.003069581, 0.003075749, 0.003173469, 0.003267707, 
    0.003268978, 0.003243104, 0.00311075, 0.003043927, 0.00305224, 
    0.003088098, 0.003192637, 0.003295492, 0.003524214, 0.003720036, 
    0.003916413, 0.004079124, 0.004172696, 0.00423076, 0.004259782, 
    0.004236879, 0.004146231, 0.004033938, 0.003914697, 0.003843967, 
    0.003707495, 0.003687404, 0.00362106, 0.003568862, 0.00355381, 
    0.00350271, 0.003480075, 0.003466677, 0.0034998, 0.003468441, 
    0.003375124, 0.003295111, 0.003260603, 0.003182704, 0.003057629, 
    0.003192621, 0.003129791, 0.002764946, 0.002888544, 0.001275385, 
    0.002194807, 0.002791619, 0.002957445, 0.00307769, 0.003010184, 
    0.002951961, 0.002884442, 0.002971655, 0.002918312, 0.002919473, 
    0.003008436, 0.003049618, 0.003121255, 0.003266102, 0.003007386, 
    0.003182195,
  0.002709519, 0.002530927, 0.001970898, 0.001605561, 0.001704744, 
    0.002119576, 0.002333246, 0.002142337, 0.002559475, 0.003067055, 
    0.00297952, 0.003296824, 0.003573009, 0.003283155, 0.003303723, 
    0.003412412, 0.003548581, 0.003561057, 0.003595183, 0.003614988, 
    0.003342874, 0.003192047, 0.003274892, 0.003080977, 0.002947431, 
    0.002905359, 0.002703132, 0.002737209, 0.002856309, 0.002938515, 
    0.00297752, 0.003043689, 0.003096443, 0.00297752, 0.003015969, 
    0.003077006, 0.003154473, 0.003192192, 0.003219228, 0.003243197, 
    0.003239684, 0.003195593, 0.00314907, 0.003098384, 0.003072793, 
    0.003012234, 0.002907839, 0.002887318, 0.002899129, 0.002900623, 
    0.002878465, 0.002904484, 0.002950039, 0.002995068, 0.00299111, 
    0.002993511, 0.002947129, 0.002911575, 0.00293443, 0.003048124, 
    0.003140122, 0.003208341, 0.003331557, 0.003385756, 0.003425922, 
    0.003458299, 0.003464673, 0.003521465, 0.003533797, 0.003571484, 
    0.003572041, 0.003586473, 0.003435507, 0.003346194, 0.003217099, 
    0.003307745, 0.003165888, 0.002840145, 0.002787359, 0.002727563, 
    0.002863685, 0.002756156, 0.002843259, 0.002764454, 0.002697125, 
    0.002694009, 0.002768045, 0.002923321, 0.0030383, 0.003130505, 
    0.003157988, 0.00326696, 0.003255088, 0.003199297, 0.002763132, 
    0.002638057,
  0.001945564, 0.001889664, 0.001759931, 0.001812033, 0.002050596, 
    0.002163956, 0.001995616, 0.002368423, 0.002476504, 0.003592542, 
    0.003591669, 0.003422058, 0.003623506, 0.00327802, 0.003266465, 
    0.003333321, 0.003421504, 0.00352137, 0.003599841, 0.003703838, 
    0.003120189, 0.00299761, 0.00316274, 0.002979841, 0.002709839, 
    0.002526114, 0.002155595, 0.001927618, 0.002038896, 0.002427122, 
    0.002906868, 0.002900479, 0.002885904, 0.002939435, 0.003026333, 
    0.003040589, 0.003088718, 0.003145002, 0.003134511, 0.00316228, 
    0.003184577, 0.003181271, 0.003183801, 0.003174072, 0.003127106, 
    0.003123958, 0.003102658, 0.003120603, 0.003125865, 0.00316851, 
    0.003119618, 0.003102928, 0.003079865, 0.003068961, 0.003027795, 
    0.003013441, 0.002991602, 0.002926085, 0.002896935, 0.002922986, 
    0.00299092, 0.00301748, 0.00314961, 0.003226509, 0.003402272, 
    0.003628116, 0.0036439, 0.003784709, 0.003828706, 0.00378808, 
    0.003904331, 0.003762871, 0.003202382, 0.002901243, 0.003028462, 
    0.00306928, 0.002917534, 0.002820021, 0.002806703, 0.002760988, 
    0.002715658, 0.002651569, 0.002706645, 0.002590088, 0.002726067, 
    0.002718693, 0.002785258, 0.002867578, 0.002981097, 0.00300017, 
    0.003161483, 0.003110606, 0.00245945, 0.002215294, 0.002034461, 
    0.001515855,
  0.001254389, 0.001282125, 0.001351712, 0.001288817, 0.001035315, 
    0.001182291, 0.001254803, 0.001137325, 0.001242771, 0.002275105, 
    0.003766396, 0.003457566, 0.002954424, 0.003036647, 0.003202697, 
    0.003190825, 0.003308795, 0.003433201, 0.003550978, 0.003701165, 
    0.003281151, 0.002988867, 0.003293948, 0.003152598, 0.002777616, 
    0.002427105, 0.001732877, 0.001183671, 0.001142187, 0.002000146, 
    0.002763085, 0.002877669, 0.002825711, 0.002764661, 0.003004652, 
    0.002983941, 0.003021453, 0.003133764, 0.003151231, 0.003119508, 
    0.003095459, 0.003142267, 0.003116138, 0.003122671, 0.003081724, 
    0.003046406, 0.002950436, 0.00291248, 0.002913067, 0.002899589, 
    0.002906233, 0.002924051, 0.002933696, 0.002923794, 0.002939865, 
    0.002918584, 0.002876891, 0.00280109, 0.002707662, 0.002594447, 
    0.002527671, 0.002506245, 0.002497822, 0.002622766, 0.002882754, 
    0.003188618, 0.003526138, 0.003695002, 0.003574265, 0.002986338, 
    0.00294735, 0.002821211, 0.002480463, 0.003055977, 0.003214698, 
    0.002975501, 0.002876796, 0.002821069, 0.002786579, 0.002663204, 
    0.002671834, 0.002584619, 0.002493769, 0.00245985, 0.002484327, 
    0.00238481, 0.002505688, 0.002512173, 0.002686268, 0.002669483, 
    0.002872568, 0.002785036, 0.001698609, 0.00127181, 0.001069536, 
    0.0009766794,
  0.0009068227, 0.0009178058, 0.0008619684, 0.0009839106, 0.0006495698, 
    0.0009761231, 0.0009673811, 0.001071156, 0.0008348203, 0.001734977, 
    0.00361483, 0.002759349, 0.002227583, 0.001867475, 0.00195569, 0.0026482, 
    0.00319742, 0.003197644, 0.003147259, 0.003191302, 0.002997703, 
    0.002723729, 0.002835086, 0.002770633, 0.002723126, 0.002342467, 
    0.001847143, 0.001379813, 0.0008090064, 0.001136067, 0.002069301, 
    0.00250542, 0.002647515, 0.002556138, 0.002746716, 0.002897285, 
    0.002972163, 0.003023695, 0.003043959, 0.003078021, 0.003091278, 
    0.003101291, 0.003091151, 0.003110779, 0.003019258, 0.002964884, 
    0.00288263, 0.002875699, 0.00285014, 0.002772352, 0.002771989, 
    0.002776215, 0.002805144, 0.002753073, 0.002761466, 0.002695645, 
    0.00261474, 0.002548445, 0.002461933, 0.002373604, 0.002251757, 
    0.002169152, 0.002048432, 0.002082095, 0.002188927, 0.00248215, 
    0.003087111, 0.003144156, 0.002594935, 0.00214415, 0.002199844, 
    0.002436863, 0.002159282, 0.003058406, 0.003217768, 0.003145875, 
    0.003027063, 0.002867082, 0.002798053, 0.002746506, 0.002660884, 
    0.002470039, 0.002423737, 0.002332723, 0.00225578, 0.002251423, 
    0.002310358, 0.00224357, 0.002337125, 0.002308914, 0.002461899, 
    0.002420158, 0.001080439, 0.0007171051, 0.000346873, 0.0003820322,
  0.001027208, 0.0008759077, 0.000740136, 0.0007444913, 0.0008700746, 
    0.001000267, 0.0008136167, 0.00110285, 0.0008351698, 0.001446714, 
    0.003023962, 0.002029838, 0.001982822, 0.001920722, 0.00155254, 
    0.002103589, 0.002946063, 0.002906596, 0.002289808, 0.002029394, 
    0.002172635, 0.002475474, 0.002078745, 0.001673321, 0.001885846, 
    0.002018279, 0.001817215, 0.001641072, 0.0009350991, 0.0007367195, 
    0.001201809, 0.001571134, 0.002279048, 0.002326842, 0.002400467, 
    0.002553008, 0.002666827, 0.00274967, 0.002793541, 0.002840986, 
    0.002832435, 0.002863493, 0.002908746, 0.00291766, 0.002876144, 
    0.002858007, 0.002789151, 0.002706597, 0.002631782, 0.002585972, 
    0.002547493, 0.00248679, 0.002520423, 0.002485296, 0.002500951, 
    0.002439343, 0.002345471, 0.002256476, 0.002151255, 0.002133135, 
    0.002056077, 0.001996504, 0.001910388, 0.001811285, 0.001789176, 
    0.001927285, 0.00224303, 0.001830932, 0.001811047, 0.001888884, 
    0.00222405, 0.003054546, 0.003003014, 0.003028668, 0.003090579, 
    0.003114993, 0.003014587, 0.003006766, 0.002950929, 0.00282657, 
    0.002758587, 0.002697887, 0.002572145, 0.002359077, 0.002330515, 
    0.002242887, 0.002192836, 0.002249165, 0.002259943, 0.002195997, 
    0.00218166, 0.002276932, 0.001132733, 0.0007072347, 0.0007634377, 
    0.0007489258,
  0.0005095534, 0.0009580352, 0.0008826945, 0.0008701854, 0.001332765, 
    0.001534404, 0.001190525, 0.001330953, 0.001148293, 0.000781239, 
    0.001235235, 0.001399491, 0.002153768, 0.002290001, 0.002122535, 
    0.001823877, 0.001740811, 0.001625051, 0.001448922, 0.001327998, 
    0.001528747, 0.001604436, 0.001433569, 0.0009921289, 0.00133472, 
    0.001432728, 0.001313438, 0.001454567, 0.0009636618, 0.0005818428, 
    0.000548623, 0.0007340973, 0.001231962, 0.001945929, 0.002066774, 
    0.002139778, 0.002258463, 0.002389071, 0.002410051, 0.002403487, 
    0.002399735, 0.002448276, 0.002475251, 0.002497282, 0.002523713, 
    0.002554009, 0.002501668, 0.002416283, 0.002380884, 0.002373224, 
    0.002366357, 0.002333835, 0.00233603, 0.002286232, 0.002262343, 
    0.002213434, 0.002150268, 0.00207612, 0.001938457, 0.001920226, 
    0.001851959, 0.001811269, 0.00173701, 0.001651831, 0.001656742, 
    0.001555827, 0.001043198, 0.001058425, 0.001250861, 0.001532655, 
    0.002007378, 0.002828728, 0.003058281, 0.003019559, 0.002854048, 
    0.002833118, 0.002831209, 0.002857515, 0.002822421, 0.002714624, 
    0.002633052, 0.002545965, 0.002444129, 0.002377657, 0.002353163, 
    0.002219141, 0.002237117, 0.002217582, 0.002123772, 0.002097816, 
    0.001979657, 0.00211592, 0.002120053, 0.0008266354, 0.0003491142, 
    5.781441e-005,
  0.0003467933, 0.0004296037, 0.0004519997, 0.001258125, 0.001583073, 
    0.00189354, 0.001256202, 0.001464183, 0.001972567, 0.0008035405, 
    0.0006962032, 0.0009742947, 0.001468107, 0.001661751, 0.001657586, 
    0.001555956, 0.001302645, 0.001187107, 0.00124277, 0.001078198, 
    0.0007050895, 0.0009045028, 0.0009468456, 0.0007665695, 0.0008585041, 
    0.0008975561, 0.0009855961, 0.001324119, 0.001080662, 0.0008499511, 
    0.0006438466, 0.0005016215, 0.00073459, 0.001286527, 0.001491169, 
    0.001772502, 0.00192555, 0.001952428, 0.001984965, 0.001952079, 
    0.001898769, 0.001904427, 0.001926568, 0.001940222, 0.001984456, 
    0.002041216, 0.002060132, 0.002049847, 0.002066552, 0.002092619, 
    0.00212746, 0.002171249, 0.002209777, 0.002269127, 0.002301124, 
    0.002260814, 0.002156118, 0.002034031, 0.001893158, 0.001832521, 
    0.001694412, 0.001603972, 0.001528583, 0.001433439, 0.001391032, 
    0.00111865, 0.0008847774, 0.000771306, 0.0008826316, 0.001119651, 
    0.001349202, 0.00196362, 0.002198572, 0.002119449, 0.00231675, 
    0.002498932, 0.002507214, 0.002412022, 0.002349445, 0.002263741, 
    0.002232143, 0.002238517, 0.002220666, 0.002171664, 0.002104684, 
    0.002099867, 0.002192995, 0.002142782, 0.002114346, 0.002046286, 
    0.001823873, 0.001855837, 0.001913121, 0.001741396, 0.0004890184, 
    0.0001234105,
  0.0002850271, 0.0006388091, 0.0009539509, 0.001931241, 0.001948852, 
    0.00185536, 0.001616274, 0.001487353, 0.001708018, 0.001652721, 
    0.0007393416, 0.0008301949, 0.0009873919, 0.001047616, 0.001308685, 
    0.001310624, 0.001277245, 0.001273844, 0.001102597, 0.001044772, 
    0.0008251413, 0.0008304501, 0.0007334771, 0.0006299879, 0.0007239722, 
    0.0008190854, 0.0008077836, 0.0009459234, 0.0009862799, 0.0009297584, 
    0.0007262921, 0.0006102298, 0.0007729898, 0.001059189, 0.0007068999, 
    0.001366843, 0.001230771, 0.001219469, 0.001648209, 0.001691297, 
    0.001612095, 0.001588873, 0.001576476, 0.001554763, 0.001532462, 
    0.001516473, 0.001533669, 0.001586075, 0.001680695, 0.001738726, 
    0.001771739, 0.001869299, 0.001957531, 0.002032219, 0.002078123, 
    0.002097466, 0.002028326, 0.001887626, 0.001795391, 0.001745593, 
    0.001590716, 0.001472302, 0.001412841, 0.001218865, 0.0007846416, 
    0.0006741579, 0.0007548067, 0.0008017435, 0.0008019181, 0.0006340719, 
    0.0009209216, 0.00135095, 0.001627754, 0.001763415, 0.001804486, 
    0.001912106, 0.002189306, 0.002157246, 0.002094256, 0.001986617, 
    0.001897099, 0.001849861, 0.001833204, 0.001823238, 0.001795375, 
    0.001775745, 0.001804021, 0.001966416, 0.002114029, 0.002005898, 
    0.001823906, 0.001689008, 0.001584946, 0.001735308, 0.001624429, 
    0.0004281742,
  0.0008735717, 0.001727902, 0.001879219, 0.001885354, 0.001855821, 
    0.001830455, 0.001395295, 0.00087106, 0.0007139095, 0.0006598532, 
    0.0006501093, 0.000683615, 0.0008841888, 0.001232265, 0.00146434, 
    0.001157177, 0.0009370542, 0.000914786, 0.001003319, 0.0009769818, 
    0.0009402973, 0.0008853181, 0.0007168194, 0.0006880661, 0.0008024916, 
    0.0008180204, 0.0006935024, 0.0006616015, 0.0006344533, 0.0006474708, 
    0.0005713676, 0.000613075, 0.0006755725, 0.0007046596, 0.000694185, 
    0.001258062, 0.00129322, 0.000962819, 0.001272812, 0.001358593, 
    0.001385948, 0.001384215, 0.001375695, 0.001425304, 0.001435492, 
    0.001373217, 0.001335498, 0.001349995, 0.001387919, 0.001399205, 
    0.001397408, 0.001451799, 0.001528173, 0.001596916, 0.001638783, 
    0.001664866, 0.001682684, 0.001666885, 0.001644108, 0.001585742, 
    0.001448653, 0.001305046, 0.001229275, 0.000975138, 0.0006618709, 
    0.0005490833, 0.0006469782, 0.0006129637, 0.0007218099, 0.000792319, 
    0.0009306646, 0.001058536, 0.001199776, 0.001354812, 0.001444632, 
    0.001501789, 0.001614387, 0.002077077, 0.0020652, 0.001943957, 
    0.001769847, 0.00161672, 0.001637033, 0.001696637, 0.001657155, 
    0.001545448, 0.001471109, 0.001509972, 0.001653897, 0.001733258, 
    0.0017595, 0.001655772, 0.001460986, 0.001438177, 0.0009327624, 
    0.0004275539,
  0.001134258, 0.001586315, 0.001671319, 0.001308845, 0.001685131, 
    0.001404752, 0.001348024, 0.00118973, 0.001019833, 0.0008564363, 
    0.0008236617, 0.0008420998, 0.0009259912, 0.001198902, 0.001138995, 
    0.0009374672, 0.000910606, 0.0008901651, 0.0008650515, 0.0009964367, 
    0.0009446207, 0.0007890924, 0.0006969356, 0.000706234, 0.0006190361, 
    0.0005127012, 0.0004921813, 0.0005348581, 0.0006875099, 0.0007485931, 
    0.0007298215, 0.0006863656, 0.0007635815, 0.0007587021, 0.0006776714, 
    0.0007427598, 0.001014524, 0.001088593, 0.0008466137, 0.00105682, 
    0.0009923992, 0.0009720381, 0.0009567947, 0.0009809393, 0.001008675, 
    0.001034504, 0.001083555, 0.001098845, 0.001110115, 0.001165921, 
    0.001219899, 0.001241579, 0.001263323, 0.001284718, 0.001304014, 
    0.001281571, 0.001268283, 0.001305872, 0.001324436, 0.001326899, 
    0.001277038, 0.001162534, 0.001080471, 0.0008650203, 0.0006952817, 
    0.0006034905, 0.0005606704, 0.000480101, 0.0005889947, 0.0007749456, 
    0.0009280262, 0.0008858258, 0.0009034048, 0.001094712, 0.001343876, 
    0.001132001, 0.001116344, 0.00130708, 0.00168178, 0.001730956, 
    0.001648082, 0.001513471, 0.001472844, 0.00133952, 0.001253864, 
    0.001252387, 0.001162645, 0.001077116, 0.001179923, 0.00135791, 
    0.001495413, 0.001497719, 0.001396836, 0.001359849, 0.001134735, 
    0.0009713541,
  0.001076196, 0.0009288685, 0.0008343426, 0.0008798488, 0.0009771721, 
    0.001038874, 0.001042769, 0.001050557, 0.001019118, 0.0009308236, 
    0.0009018164, 0.0008064169, 0.0007885511, 0.0008931055, 0.0009113047, 
    0.00079022, 0.0007933518, 0.0008656397, 0.000809548, 0.0009038509, 
    0.0009878059, 0.0008613332, 0.0007286771, 0.0006170335, 0.0005077104, 
    0.0004657966, 0.0004515388, 0.0004498861, 0.0004690232, 0.0005139095, 
    0.0005317591, 0.0005404375, 0.0006002967, 0.000682503, 0.0006729664, 
    0.0006150942, 0.0006272695, 0.000861682, 0.0008610939, 0.0008041915, 
    0.0007775521, 0.0007693027, 0.0007577157, 0.000757413, 0.0007663937, 
    0.0008165101, 0.0008685323, 0.0008791503, 0.0009174715, 0.0009853737, 
    0.001021311, 0.001044009, 0.001076847, 0.001114581, 0.00115036, 
    0.001169863, 0.001164252, 0.001181784, 0.001189508, 0.001167623, 
    0.001116091, 0.001044518, 0.001014032, 0.0007997416, 0.0007021483, 
    0.0005875484, 0.0005118425, 0.0005248284, 0.000642766, 0.0007760897, 
    0.0008909439, 0.000630066, 0.0006747299, 0.001081694, 0.001016162, 
    0.0009728326, 0.0009169632, 0.0009873922, 0.001082664, 0.001171339, 
    0.001300659, 0.001181672, 0.0009181397, 0.0008216123, 0.0008607609, 
    0.0009543477, 0.0008489517, 0.0007120683, 0.0007332386, 0.0008784188, 
    0.0010346, 0.001177062, 0.001168096, 0.001123291, 0.001199394, 0.001129474,
  0.0008885763, 0.0009153578, 0.0008681985, 0.0007755333, 0.0007302179, 
    0.0007541552, 0.000774119, 0.0007862307, 0.0008219297, 0.0008305924, 
    0.0008536715, 0.0007937804, 0.0007105565, 0.0007396278, 0.0007356699, 
    0.0006018535, 0.0005757553, 0.0005936367, 0.0005423289, 0.0005511189, 
    0.0006676896, 0.0007341765, 0.0006629211, 0.0005564117, 0.0004967116, 
    0.0004132965, 0.0003926494, 0.0003900587, 0.000498301, 0.0005480828, 
    0.0005311868, 0.0005562684, 0.0006132979, 0.0006047945, 0.0005726396, 
    0.0005264499, 0.000507901, 0.0005074719, 0.0005734817, 0.0006008202, 
    0.0006666239, 0.0006798797, 0.0006840124, 0.0006704386, 0.0006794031, 
    0.000756253, 0.0008132346, 0.0008370928, 0.0008660848, 0.0009089364, 
    0.0009343997, 0.0009844834, 0.001049238, 0.00108775, 0.001094569, 
    0.001092519, 0.001077848, 0.001082569, 0.001077642, 0.001035633, 
    0.0009958488, 0.000988394, 0.0008468358, 0.0007651227, 0.0006845051, 
    0.0006143146, 0.000619258, 0.000677448, 0.0007338577, 0.0006966325, 
    0.0006305589, 0.0006036812, 0.0006103572, 0.000655879, 0.0007398501, 
    0.0008233124, 0.0008533054, 0.000830322, 0.0008307192, 0.0009089208, 
    0.00111733, 0.0009888385, 0.0008044136, 0.0007850225, 0.0007872474, 
    0.0007014014, 0.0005182163, 0.0002931021, 0.0002087969, 0.0003068349, 
    0.0005149744, 0.0007186644, 0.0007746448, 0.000748069, 0.0007916996, 
    0.0009410609,
  0.0006030132, 0.0008499208, 0.0008842833, 0.000855817, 0.000763851, 
    0.0007535513, 0.0007883923, 0.0007304407, 0.0006579452, 0.0006298916, 
    0.0006449595, 0.0006148871, 0.0005549327, 0.0005565542, 0.0005460642, 
    0.0005308215, 0.0005190913, 0.000542806, 0.0004928494, 0.0004540667, 
    0.0005326176, 0.0005736733, 0.0005433464, 0.0005014164, 0.0004787666, 
    0.0004591845, 0.0004700405, 0.0004790208, 0.0004862049, 0.0004681009, 
    0.0004162051, 0.000428142, 0.000471407, 0.0004468341, 0.0003810784, 
    0.0003396253, 0.0003521343, 0.0004141228, 0.0005188042, 0.0005509588, 
    0.0006166832, 0.0006583428, 0.0005179946, 0.0006146329, 0.0006058111, 
    0.0006709313, 0.0007271185, 0.0007834169, 0.0008365689, 0.000882742, 
    0.0009102393, 0.0009609121, 0.001028082, 0.001074701, 0.001081837, 
    0.00107405, 0.001061254, 0.001059077, 0.001075226, 0.001065785, 
    0.001018752, 0.0009499127, 0.000872649, 0.000737895, 0.0006446897, 
    0.0006148552, 0.0006157295, 0.0006593917, 0.0006639375, 0.0006547188, 
    0.0006326579, 0.0006396673, 0.0006684682, 0.0007137673, 0.0007699544, 
    0.0008929945, 0.0009226699, 0.0009137217, 0.0009047093, 0.0009292667, 
    0.000945224, 0.0007440303, 0.0006714237, 0.0006160312, 0.0006121048, 
    0.0006044442, 0.0004924187, 0.0002905419, 0.0001056087, 6.202655e-005, 
    0.000202137, 0.0003772955, 0.0004715342, 0.0005350974, 0.0005321875, 
    0.0005467143,
  0.000572592, 0.0006939792, 0.0006883838, 0.0006172713, 0.0006032996, 
    0.0007515643, 0.0007584151, 0.0006756522, 0.0006291762, 0.0006018851, 
    0.000633277, 0.0006098642, 0.0005599237, 0.0005363366, 0.0005608462, 
    0.0005872946, 0.0005654874, 0.0005562687, 0.0005322044, 0.0005149269, 
    0.0005008917, 0.0005053106, 0.0005371473, 0.000551071, 0.0005373699, 
    0.0004974585, 0.0004858077, 0.000486952, 0.0004723447, 0.0004201949, 
    0.0003664395, 0.0003620368, 0.0003825088, 0.0003638805, 0.0003173571, 
    0.0002969007, 0.000311937, 0.0003692688, 0.0004668294, 0.0004787976, 
    0.0005072171, 0.0005137818, 0.0004164599, 0.0004356607, 0.0005795057, 
    0.0006873028, 0.0007673476, 0.00079022, 0.0008474723, 0.0009128468, 
    0.0009594494, 0.0009816387, 0.0009947829, 0.001041433, 0.0009308234, 
    0.001024124, 0.001002508, 0.001003827, 0.001027844, 0.001023091, 
    0.0009450337, 0.0008998925, 0.0007481477, 0.0006831549, 0.0006566904, 
    0.0006667352, 0.00062951, 0.0005839569, 0.000593001, 0.0006258711, 
    0.0006515725, 0.0006952826, 0.0007707332, 0.0008226288, 0.0008877013, 
    0.0009789679, 0.001037811, 0.00100591, 0.0009946885, 0.0009385491, 
    0.0006866509, 0.0006387134, 0.0005826526, 0.0005552028, 0.0005867851, 
    0.0005603367, 0.0005327282, 0.0004324331, 0.0003002058, 0.0002606446, 
    0.0003130813, 0.0003882153, 0.0004332447, 0.0004835981, 0.0005432349, 
    0.0005346029,
  0.0005277218, 0.0006349306, 0.0004825012, 0.0005504664, 0.0005806182, 
    0.0006454047, 0.0005485276, 0.0004808959, 0.0004394108, 0.000440476, 
    0.000497649, 0.0005529942, 0.0005778533, 0.0005854828, 0.0006053988, 
    0.0006114386, 0.0006032848, 0.000580349, 0.0005714954, 0.0005671403, 
    0.0005740387, 0.0005538366, 0.0005260051, 0.0005036254, 0.0004675448, 
    0.0004428445, 0.0004436233, 0.0004519363, 0.0004520317, 0.0004255992, 
    0.0004120569, 0.0003826997, 0.0003627838, 0.0003260832, 0.0002901137, 
    0.0002446233, 0.0002120236, 0.0002005, 0.0001963197, 0.0002046803, 
    0.0002344986, 0.0002487244, 0.0002543351, 0.0002790829, 0.000329898, 
    0.0004214663, 0.0005571109, 0.0007078224, 0.000850826, 0.0009709259, 
    0.001028639, 0.00101578, 0.0009399001, 0.0009193802, 0.0009184424, 
    0.0009030246, 0.0008478547, 0.0007743263, 0.0006772422, 0.0006477896, 
    0.0006780687, 0.0006753666, 0.0006290021, 0.0005516752, 0.00055096, 
    0.0005961959, 0.0006329124, 0.000637013, 0.0006388249, 0.0006596785, 
    0.0007295195, 0.000779476, 0.0008421005, 0.0009274383, 0.001067422, 
    0.00114939, 0.001073097, 0.001018022, 0.001064482, 0.0008282722, 
    0.0006337697, 0.0005510862, 0.0004693882, 0.0003988796, 0.0004329425, 
    0.0003879128, 0.0004978874, 0.0004868563, 0.0004473901, 0.0004075421, 
    0.0003984659, 0.0003950968, 0.0003537708, 0.0003379402, 0.0004085433, 
    0.000468005,
  0.0003443928, 0.0003822851, 0.0003537862, 0.0003537869, 0.0003673451, 
    0.0003826991, 0.0004496155, 0.0004343407, 0.0004745864, 0.0005340956, 
    0.0005963545, 0.0006360118, 0.0006501897, 0.0006556893, 0.0006482187, 
    0.0006333092, 0.0005958779, 0.0005576195, 0.0005398492, 0.0005466997, 
    0.0005720198, 0.0005774557, 0.0005571424, 0.0005090771, 0.000446723, 
    0.000393826, 0.0003723683, 0.00037089, 0.0003719708, 0.0003711125, 
    0.0003435513, 0.0003280223, 0.0003120959, 0.0002845507, 0.0002438127, 
    0.0002158224, 0.0002051094, 0.0001848598, 0.0001692672, 0.0001577595, 
    0.0001695851, 0.0002118011, 0.0002416988, 0.0002598028, 0.0002718668, 
    0.0002997458, 0.0003738623, 0.0004789572, 0.0006735066, 0.0009217162, 
    0.001146068, 0.001169211, 0.0009602293, 0.0007713694, 0.0006578983, 
    0.0005960364, 0.0005488455, 0.0004788141, 0.0004129627, 0.0004032035, 
    0.000430272, 0.0004793545, 0.0004942956, 0.0004579766, 0.0004265369, 
    0.0004415414, 0.0004886845, 0.0005459208, 0.0005929688, 0.000634247, 
    0.0006697237, 0.0007241784, 0.0008365849, 0.00100041, 0.001450354, 
    0.001450767, 0.001379576, 0.0009144365, 0.0008210557, 0.0008185131, 
    0.0007031662, 0.0005551078, 0.0004531287, 0.0002745687, 0.0002007859, 
    0.0001821736, 0.00020298, 0.0002200976, 0.0002587694, 0.000256401, 
    0.0002929741, 0.0003555038, 0.0003456655, 0.0002843123, 0.0002797665, 
    0.0002901605,
  0.0003289282, 0.0003041807, 0.0003027502, 0.0003307397, 0.00035509, 
    0.0003605101, 0.0004088776, 0.0004567208, 0.0005035463, 0.0005572382, 
    0.0006118361, 0.0005619263, 0.0005525802, 0.0005707478, 0.0006502373, 
    0.0006804526, 0.0006838861, 0.0006692628, 0.0006439904, 0.0006111045, 
    0.0005658845, 0.0005186457, 0.0004758578, 0.0004381877, 0.000404046, 
    0.0003645957, 0.000342693, 0.0003289601, 0.0003079157, 0.0002771913, 
    0.000255225, 0.0002366761, 0.0002239763, 0.0002065082, 0.0002079069, 
    0.0002271553, 0.0002408564, 0.0002694507, 0.0002605974, 0.0002700547, 
    0.0002831041, 0.0002969324, 0.0003271799, 0.0003258607, 0.0003101409, 
    0.0003127794, 0.0003443937, 0.0004381398, 0.0006156504, 0.001328554, 
    0.001662976, 0.001610603, 0.001497704, 0.0008305926, 0.0006790538, 
    0.0006085295, 0.0005886295, 0.0005927621, 0.0005568085, 0.0005473195, 
    0.0005263863, 0.0005067724, 0.0004768111, 0.0004377265, 0.0004332761, 
    0.0004573563, 0.0005244472, 0.0006465493, 0.0007603546, 0.001122131, 
    0.0008502862, 0.0008367121, 0.0008466939, 0.001370325, 0.0009043275, 
    0.001140966, 0.0009143887, 0.0009158354, 0.0009239413, 0.001194865, 
    0.0009022775, 0.0006299082, 0.0003183741, 0.0001604776, 8.893598e-005, 
    7.37567e-005, 8.686967e-005, 0.0001283707, 0.0001940787, 0.0002773025, 
    0.0005318702, 0.0005794421, 0.0005564585, 0.0005711454, 0.0004602331, 
    0.0003812844,
  0.0005815562, 0.0005018925, 0.000440333, 0.0004097517, 0.0003786618, 
    0.0003851943, 0.000467926, 0.0005743401, 0.0006391103, 0.000655116, 
    0.000637616, 0.0006186857, 0.000644753, 0.0007733239, 0.0009440961, 
    0.000865497, 0.001198266, 0.00124932, 0.001211475, 0.0007690489, 
    0.0006597102, 0.0005600034, 0.0004833282, 0.0004200359, 0.0003746888, 
    0.0003421526, 0.0003139238, 0.0002835651, 0.0002598504, 0.0002471188, 
    0.0002350708, 0.0002500434, 0.0002812445, 0.0003310899, 0.0003857514, 
    0.0006411771, 0.0007121782, 0.0007489105, 0.0004069548, 0.0003759126, 
    0.0005043091, 0.0004839004, 0.0004725993, 0.0004760961, 0.0004741253, 
    0.0004630308, 0.0004566094, 0.0004751742, 0.0005265613, 0.0006123761, 
    0.0006890038, 0.0007109541, 0.0007017194, 0.0006813585, 0.000669978, 
    0.0006761292, 0.0006986675, 0.0007257361, 0.0007466691, 0.0007485609, 
    0.0007251003, 0.0006693264, 0.0005961796, 0.000420942, 0.0003998022, 
    0.0004157922, 0.0004659236, 0.0005480031, 0.0006382207, 0.001222569, 
    0.0007395644, 0.0007209043, 0.001210521, 0.0006667353, 0.000679626, 
    0.0007186789, 0.0007947821, 0.001234522, 0.001302217, 0.001204195, 
    0.0009786986, 0.0004529377, 0.0002544146, 0.0001394809, 8.475568e-005, 
    6.563458e-005, 6.776447e-005, 8.691743e-005, 0.0001342197, 0.0002170781, 
    0.0003539941, 0.0007840217, 0.0009666188, 0.000957543, 0.0007457789, 
    0.0006558155,
  0.0006505393, 0.0005031801, 0.000507996, 0.0005270536, 0.0004888272, 
    0.0005472079, 0.0007149596, 0.0008999093, 0.001017497, 0.001055612, 
    0.001081537, 0.001103551, 0.001136325, 0.001147149, 0.001111593, 
    0.001091279, 0.001089467, 0.001070029, 0.001023823, 0.0009510578, 
    0.0008726973, 0.0007845302, 0.0007126548, 0.0006334521, 0.0005649944, 
    0.0004306377, 0.0003910919, 0.0003351272, 0.0003017962, 0.0002917032, 
    0.0002836128, 0.0003548206, 0.0003867369, 0.0004299701, 0.0004648905, 
    0.0004760962, 0.0004658283, 0.0004334829, 0.0003881038, 0.0003567756, 
    0.0003381949, 0.0003344279, 0.0003425023, 0.0003549954, 0.0003643732, 
    0.0003671389, 0.0003621321, 0.0003550113, 0.000352039, 0.0003574114, 
    0.0003725271, 0.0003952405, 0.000418526, 0.000438124, 0.0004524768, 
    0.0004620294, 0.0004681329, 0.000474157, 0.0004799743, 0.0004882396, 
    0.0004953285, 0.0004974107, 0.0004923881, 0.0004845521, 0.0004771451, 
    0.0004086714, 0.0004131695, 0.0004211963, 0.0004328152, 0.0004454355, 
    0.0004573405, 0.0004687051, 0.0004710575, 0.0004781306, 0.0004814844, 
    0.0005891384, 0.0006179869, 0.0006579299, 0.0004169206, 0.0003532788, 
    0.0002820393, 0.0002118488, 0.0001547077, 0.0001126507, 8.281664e-005, 
    6.887707e-005, 6.995793e-005, 8.483522e-005, 0.000115623, 0.0001664379, 
    0.0002327183, 0.0003250819, 0.0004722815, 0.000596068, 0.0007175506, 
    0.0007946555,
  0.0004985072, 0.0005207438, 0.0005318698, 0.0005316791, 0.0004575787, 
    0.0004654147, 0.0004743474, 0.0005491792, 0.0005707481, 0.0005883433, 
    0.000605589, 0.0006251551, 0.0006460724, 0.0006581523, 0.0006602186, 
    0.0006525256, 0.000637235, 0.0006139018, 0.0005879779, 0.0005596221, 
    0.0005302649, 0.0005031963, 0.0004812141, 0.0004657169, 0.0004599472, 
    0.0003627519, 0.0003521185, 0.0003988803, 0.0003874521, 0.0003810148, 
    0.0003744822, 0.0003641824, 0.0003583014, 0.0003517688, 0.000341326, 
    0.000328356, 0.0003141304, 0.0002993166, 0.0002850592, 0.0002749502, 
    0.0002680997, 0.0002653817, 0.0002655406, 0.0002689421, 0.000274823, 
    0.0002823412, 0.0002890487, 0.0002943735, 0.0002995869, 0.000303799, 
    0.0003071527, 0.0003085196, 0.0003063262, 0.0003014307, 0.0002950887, 
    0.0002889692, 0.0002851228, 0.0002852658, 0.0002907176, 0.0003023685, 
    0.0003201862, 0.0003412466, 0.0003612419, 0.0003780107, 0.0003884057, 
    0.000388962, 0.0003922363, 0.0003903131, 0.0003798386, 0.000373592, 
    0.000372845, 0.0002821664, 0.0002805293, 0.0002618213, 0.0002501547, 
    0.0002374073, 0.0002222915, 0.0002043466, 0.0001864333, 0.000168838, 
    0.0001525461, 0.0001397828, 0.0001317719, 0.0001263836, 0.0001233637, 
    0.0001231729, 0.0001283705, 0.0001372555, 0.0001512428, 0.0001730342, 
    0.0002043306, 0.0002427479, 0.0003282289, 0.0003756425, 0.0004253766, 
    0.0004698018,
  0.0003271163, 0.0003363194, 0.0003474773, 0.0003562829, 0.0003617029, 
    0.0003719073, 0.0003827951, 0.0003935238, 0.0004026315, 0.000410849, 
    0.000418669, 0.0004259805, 0.0004306535, 0.0004317503, 0.0004304945, 
    0.0004260918, 0.0004189552, 0.0004101655, 0.0004002631, 0.0003889939, 
    0.0003781061, 0.0003678382, 0.0003586512, 0.0003507833, 0.000345252, 
    0.0003400386, 0.0003411989, 0.000337114, 0.0003341417, 0.0003345391, 
    0.0003354769, 0.0003349523, 0.0003342212, 0.0003329815, 0.0003308038, 
    0.0003269256, 0.0003219187, 0.0003170391, 0.0003131608, 0.0003093462, 
    0.0003054201, 0.000302416, 0.0003003339, 0.0002976159, 0.0002950251, 
    0.0002922594, 0.0002881745, 0.0002837082, 0.0002784153, 0.0002730906, 
    0.0002669393, 0.0002606927, 0.0002554317, 0.0002511084, 0.0002486129, 
    0.0002475797, 0.0002478182, 0.0002509335, 0.0002563218, 0.0002637287, 
    0.0002732495, 0.0002831519, 0.0002920846, 0.0003007631, 0.0003077567, 
    0.000312684, 0.0003166576, 0.0003185491, 0.000319312, 0.0003193756, 
    0.0003181676, 0.0003115714, 0.0003123025, 0.0003138761, 0.0003124615, 
    0.0003146867, 0.0003137013, 0.0003108879, 0.000307566, 0.0003035128, 
    0.0002934039, 0.0002857904, 0.0002771755, 0.0002693553, 0.0002638717, 
    0.0002608517, 0.0002602636, 0.000262012, 0.0002654771, 0.0002703727, 
    0.0002775093, 0.0002882541, 0.0002940079, 0.0003017803, 0.0003099184, 
    0.0003189624,
  0.000299428, 0.0003006995, 0.0003036241, 0.0003067713, 0.0003104428, 
    0.0003151477, 0.0003190578, 0.0003224751, 0.0003257812, 0.0003291667, 
    0.0003320278, 0.0003345073, 0.0003373206, 0.0003395618, 0.0003404995, 
    0.0003406426, 0.0003399432, 0.0003385127, 0.0003371299, 0.000335906, 
    0.0003344596, 0.0003327112, 0.0003306926, 0.0003283879, 0.0003257812, 
    0.0003231109, 0.0003204247, 0.000317818, 0.0003155769, 0.000312843, 
    0.0003108879, 0.0003089011, 0.0003066918, 0.0003045778, 0.0003027817, 
    0.0003009538, 0.0002986491, 0.0002961855, 0.0002937854, 0.0002913535, 
    0.0002886991, 0.0002862354, 0.0002842168, 0.0002816895, 0.0002791941, 
    0.0002763965, 0.0002732812, 0.0002711673, 0.0002691963, 0.0002673526, 
    0.0002658108, 0.0002636333, 0.0002616306, 0.0002602001, 0.0002588967, 
    0.0002580066, 0.0002580861, 0.0002577523, 0.0002577205, 0.0002579748, 
    0.0002585471, 0.0002605657, 0.0002616941, 0.0002633313, 0.0002641896, 
    0.0002652864, 0.0002670824, 0.0002681951, 0.0002689421, 0.0002700865, 
    0.0002710561, 0.0002718031, 0.0002724866, 0.0002737264, 0.000275284, 
    0.0002758721, 0.0002766192, 0.0002765238, 0.0002765397, 0.0002769211, 
    0.0002770483, 0.000277096, 0.0002768258, 0.0002768735, 0.0002772867, 
    0.0002779066, 0.0002788763, 0.0002808154, 0.0002834062, 0.0002854566, 
    0.0002869348, 0.000288413, 0.0002903203, 0.0002916555, 0.000293086, 
    0.0002952318,
  9.013433e-005, 8.579512e-005, 8.198043e-005, 7.846771e-005, 7.557485e-005, 
    7.279334e-005, 7.055223e-005, 6.880378e-005, 6.759577e-005, 
    6.653086e-005, 6.560891e-005, 6.498912e-005, 6.497322e-005, 
    6.537055e-005, 6.605397e-005, 6.67533e-005, 6.778646e-005, 6.88514e-005, 
    7.002763e-005, 7.134685e-005, 7.280914e-005, 7.436681e-005, 
    7.590858e-005, 7.751398e-005, 7.907161e-005, 8.042267e-005, 
    8.161477e-005, 8.239356e-005, 8.306114e-005, 8.358565e-005, 
    8.412611e-005, 8.458708e-005, 8.501625e-005, 8.56361e-005, 8.614472e-005, 
    8.682825e-005, 8.797261e-005, 8.914887e-005, 9.034091e-005, 
    9.183504e-005, 9.390141e-005, 9.620615e-005, 9.886042e-005, 0.0001018805, 
    0.0001049321, 0.0001080792, 0.0001109563, 0.0001141511, 0.0001170756, 
    0.0001199843, 0.0001232903, 0.0001259447, 0.00012817, 0.0001302998, 
    0.0001318416, 0.0001328111, 0.0001333674, 0.0001333834, 0.0001327317, 
    0.000131778, 0.0001303316, 0.0001283765, 0.0001269937, 0.0001248003, 
    0.0001225751, 0.0001204293, 0.0001184902, 0.0001171232, 0.0001168372, 
    0.000116853, 0.0001173776, 0.0001182358, 0.0001195074, 0.0001206201, 
    0.0001249911, 0.0001285992, 0.0001312377, 0.0001338444, 0.0001376272, 
    0.0001406154, 0.0001428407, 0.0001443825, 0.0001449388, 0.0001449705, 
    0.0001439215, 0.0001420141, 0.0001391372, 0.0001354974, 0.000131031, 
    0.0001261355, 0.0001208744, 0.0001154226, 0.0001098595, 0.0001045348, 
    9.946455e-005, 9.469606e-005,
  0.0001089852, 0.0001063945, 0.0001031997, 9.97188e-005, 9.612663e-005, 
    9.294768e-005, 8.959387e-005, 8.596992e-005, 8.209166e-005, 
    7.851535e-005, 7.493899e-005, 7.155348e-005, 6.905803e-005, 
    6.808847e-005, 6.850171e-005, 7.009119e-005, 7.285684e-005, 
    7.616289e-005, 7.943719e-005, 8.236177e-005, 8.387174e-005, 
    8.409427e-005, 8.360157e-005, 8.314062e-005, 8.178959e-005, 
    7.937363e-005, 7.721194e-005, 7.535229e-005, 7.417609e-005, 
    7.352442e-005, 7.390586e-005, 7.60676e-005, 7.948495e-005, 8.396723e-005, 
    8.892635e-005, 9.468017e-005, 0.0001010697, 0.0001077614, 0.0001146595, 
    0.0001208902, 0.0001257064, 0.0001299184, 0.0001344961, 0.0001385491, 
    0.0001426815, 0.0001496434, 0.0001580199, 0.0001674773, 0.0001788738, 
    0.000192098, 0.0002062124, 0.0002198339, 0.0002358395, 0.0002466321, 
    0.0002570112, 0.0002551357, 0.0002580285, 0.0002602378, 0.0002594114, 
    0.0002551198, 0.0002470138, 0.0002336941, 0.0002183875, 0.0002023499, 
    0.0001864552, 0.0001699409, 0.0001563193, 0.0001474501, 0.0001422049, 
    0.0001383902, 0.0001389784, 0.000144001, 0.0001536173, 0.0001658082, 
    0.0001810511, 0.0001983285, 0.0002158126, 0.0002321999, 0.0002462507, 
    0.0002591888, 0.0002664049, 0.0002672315, 0.0002667069, 0.0002585055, 
    0.0002506216, 0.0002370636, 0.0002214551, 0.0002032718, 0.0001854221, 
    0.0001684626, 0.0001533946, 0.0001400114, 0.0001291554, 0.0001216055, 
    0.000116265, 0.0001118304,
  0.0001047892, 9.836775e-005, 9.180326e-005, 8.641498e-005, 8.290226e-005, 
    8.080417e-005, 7.997765e-005, 8.020023e-005, 8.116971e-005, 
    8.199623e-005, 8.218692e-005, 8.145577e-005, 7.997756e-005, 
    7.857886e-005, 7.722783e-005, 7.810199e-005, 8.201206e-005, 
    8.670092e-005, 9.069056e-005, 9.351986e-005, 9.393311e-005, 
    9.266144e-005, 8.921229e-005, 8.450754e-005, 7.951664e-005, 
    7.516154e-005, 7.257075e-005, 7.228463e-005, 7.425557e-005, 
    7.776823e-005, 8.215514e-005, 8.829052e-005, 9.464839e-005, 0.000102246, 
    0.0001111469, 0.0001216375, 0.0001350364, 0.0001507721, 0.0001686693, 
    0.0001862964, 0.0002029697, 0.0002172112, 0.0002321046, 0.0002431989, 
    0.0002516867, 0.0002579013, 0.0002597295, 0.0002618118, 0.0002601745, 
    0.0002563123, 0.0002520049, 0.0002453291, 0.0002387485, 0.0002346796, 
    0.0002328993, 0.0002301655, 0.0002270185, 0.00022411, 0.000222902, 
    0.0002226792, 0.0002189757, 0.0002121567, 0.0002066097, 0.0002041302, 
    0.0002020795, 0.0001978993, 0.0001960238, 0.0001924158, 0.0001957378, 
    0.0002056243, 0.0002159715, 0.0002264301, 0.0002377311, 0.0002499541, 
    0.0002608738, 0.0002702674, 0.0002802809, 0.0002862255, 0.0002891183, 
    0.0002871474, 0.0002831101, 0.000276832, 0.0002692026, 0.0002566458, 
    0.0002402742, 0.000222965, 0.0002093276, 0.0002015075, 0.0001895073, 
    0.0001739146, 0.0001602451, 0.0001466712, 0.000134957, 0.0001253884, 
    0.0001178385, 0.000111894,
  0.0001531881, 0.0001358631, 0.0001185538, 0.0001019122, 8.835411e-005, 
    8.015253e-005, 7.935776e-005, 8.447585e-005, 9.49027e-005, 0.0001074753, 
    0.0001168214, 0.0001212242, 0.0001225275, 0.000122909, 0.0001258335, 
    0.0001320959, 0.0001396618, 0.0001450977, 0.0001447639, 0.0001375477, 
    0.0001276137, 0.0001151842, 0.0001021029, 9.440997e-005, 9.205757e-005, 
    9.404437e-005, 9.882863e-005, 0.0001054567, 0.0001109404, 0.0001149776, 
    0.000117028, 0.0001187605, 0.0001225434, 0.0001262786, 0.0001265965, 
    0.0001251978, 0.0001248004, 0.0001257859, 0.0001309833, 0.0001426499, 
    0.0001571298, 0.0001730722, 0.0001924634, 0.0002099794, 0.0002327085, 
    0.000257997, 0.0002443434, 0.0002800904, 0.0002887528, 0.0002763553, 
    0.0002613983, 0.0002467118, 0.000230992, 0.0002209786, 0.0002177835, 
    0.0002071024, 0.0001929246, 0.0002112356, 0.0001999342, 0.0001941164, 
    0.0001939737, 0.0001950227, 0.0002025249, 0.000205831, 0.0002031926, 
    0.0002047661, 0.0002035104, 0.0002096775, 0.0002186259, 0.000229466, 
    0.0002455354, 0.000266087, 0.0002833644, 0.0003007852, 0.0003131829, 
    0.000312102, 0.0003110372, 0.0003139938, 0.0003207646, 0.000334593, 
    0.0003400289, 0.000343319, 0.000343208, 0.000343764, 0.0003431283, 
    0.0003357532, 0.0003213845, 0.0003030582, 0.0002926469, 0.0002817276, 
    0.0002672317, 0.0002483964, 0.0002286077, 0.0002044003, 0.0001846115, 
    0.0001680654,
  0.000234457, 0.0002359987, 0.0002341073, 0.0002175928, 0.0001943867, 
    0.0001684151, 0.0001543643, 0.0001537445, 0.00016255, 0.0001707674, 
    0.0001658083, 0.0001518529, 0.0001322548, 0.0001183472, 0.0001148185, 
    0.0001267553, 0.0001455268, 0.0001594664, 0.0001659513, 0.0001629313, 
    0.0001544436, 0.0001445095, 0.0001345438, 0.0001240691, 0.0001147709, 
    0.0001110357, 0.0001159313, 0.0001245301, 0.0001275183, 0.0001253884, 
    0.0001199366, 0.0001199843, 0.00012817, 0.0001385491, 0.0001508674, 
    0.0001577816, 0.0001609128, 0.0001642031, 0.0001727702, 0.0001918596, 
    0.0002152405, 0.0002361735, 0.0002476175, 0.0002504946, 0.0002600314, 
    0.0002771501, 0.0002707762, 0.0002835873, 0.000272302, 0.0002455357, 
    0.0002103292, 0.0001916371, 0.000188347, 0.0001953405, 0.0002027156, 
    0.0002073091, 0.0002076272, 0.0002087557, 0.0002037648, 0.0002073885, 
    0.0002155586, 0.0002244434, 0.0002361261, 0.0002475067, 0.0002484601, 
    0.0002507016, 0.0002416095, 0.0002232196, 0.0001947049, 0.0001637102, 
    0.000232518, 0.0002252383, 0.000251337, 0.0002705536, 0.0002734782, 
    0.0002484922, 0.0002691073, 0.0002684556, 0.0002787234, 0.0002918364, 
    0.00029945, 0.0003058079, 0.0003083828, 0.0003073975, 0.0003146136, 
    0.0003248812, 0.0003305874, 0.0003239275, 0.0003096543, 0.0002862418, 
    0.0002753378, 0.0002431832, 0.0002353948, 0.0002386692, 0.0002329787, 
    0.0002304038,
  0.0002307855, 0.0001913828, 0.0002465846, 0.0002520685, 0.0002489053, 
    0.0002460602, 0.0002421978, 0.0002561692, 0.0002780402, 0.0002976381, 
    0.0003056014, 0.0002894205, 0.0002580443, 0.0002294024, 0.000216512, 
    0.0002118549, 0.0002097569, 0.0002014278, 0.0001920183, 0.0001879338, 
    0.0001975499, 0.0002243799, 0.0002272092, 0.0002053698, 0.0001796841, 
    0.0001646321, 0.0001710694, 0.0001997113, 0.0002280832, 0.0002364595, 
    0.0002214392, 0.0001943707, 0.0001836262, 0.0001904608, 0.0002002042, 
    0.0002006649, 0.0001929561, 0.0001837373, 0.0001814961, 0.0001978198, 
    0.0002243322, 0.0002503995, 0.0002437235, 0.000215193, 0.0001798752, 
    0.0001909379, 0.0002228857, 0.0002400677, 0.0002214077, 0.0001857404, 
    0.0001487695, 0.0001408539, 0.0001489602, 0.0001517578, 0.000142507, 
    0.0001292033, 0.0001285991, 0.0001421573, 0.0001593712, 0.000169639, 
    0.0001783173, 0.0001892212, 0.000197232, 0.0002048931, 0.0002021592, 
    0.0001914306, 0.0001821162, 0.0001760765, 0.0001731517, 0.0001745187, 
    0.0001899842, 0.0002036693, 0.0002156699, 0.0002317552, 0.0002413078, 
    0.0002331377, 0.0002057038, 0.0001758379, 0.0002427222, 0.0002742095, 
    0.0002947771, 0.0003061893, 0.0002952698, 0.0002848906, 0.0002912963, 
    0.0003123882, 0.0003320021, 0.0003399176, 0.000333528, 0.000321782, 
    0.0003188255, 0.0003260099, 0.0003274721, 0.0003123246, 0.0002904537, 
    0.0002639734,
  0.0002561533, 0.0002735418, 0.0002966048, 0.0003139775, 0.0003231172, 
    0.0003201924, 0.0003174904, 0.0003204467, 0.0003255489, 0.0003268365, 
    0.0003264071, 0.0003226879, 0.0003244681, 0.0003267727, 0.0003215913, 
    0.0003049655, 0.0002726042, 0.0002367778, 0.0002076908, 0.0001981859, 
    0.0002107583, 0.000230531, 0.000252879, 0.000265531, 0.0002558671, 
    0.000246664, 0.0002381445, 0.0002199295, 0.0001965645, 0.0001586082, 
    0.0001277728, 0.0001030089, 9.611086e-005, 0.0002013964, 0.0002374134, 
    0.0002551994, 0.0002277812, 0.0002129199, 0.0001881721, 0.0001596892, 
    0.0001515828, 0.0001383268, 0.0001219399, 0.0001152323, 0.0001069985, 
    9.620609e-005, 0.0001017856, 0.0001009752, 8.741673e-005, 7.857941e-005, 
    8.523883e-005, 8.686003e-005, 8.488959e-005, 7.753051e-005, 
    5.632709e-005, 4.098821e-005, 7.675122e-005, 0.0001203341, 0.0001442241, 
    0.0001391533, 0.0001311107, 0.0001502952, 0.0001784605, 0.0002015394, 
    0.0002235058, 0.0002433264, 0.0002409269, 0.0002528636, 0.0002685038, 
    0.0002912807, 0.0003124205, 0.0003169028, 0.0003200977, 0.0003112282, 
    0.0002996414, 0.0002772775, 0.0002524662, 0.0002285603, 0.0002346162, 
    0.0002606513, 0.0002249521, 0.0002034947, 0.000194387, 0.0001949591, 
    0.0002158764, 0.0002279563, 0.0002231086, 0.0002152564, 0.0002249205, 
    0.0002514962, 0.0002734785, 0.0002831263, 0.000279089, 0.0002685192, 
    0.000257377, 0.0002556923,
  0.0001700681, 0.0001487059, 0.0001444144, 0.0001504226, 0.000160754, 
    0.0001672073, 0.0001790961, 0.0002080405, 0.0002349338, 0.0002572341, 
    0.0002696477, 0.0002855104, 0.0003031853, 0.0003075087, 0.0003023746, 
    0.0002803924, 0.0002745432, 0.0002783102, 0.0002548182, 0.0002106628, 
    0.0001714192, 0.000158211, 0.0001664599, 0.0001807811, 0.0002020639, 
    0.0002144617, 0.0002043846, 0.0001800975, 0.0001584019, 0.0001457499, 
    0.0001405207, 0.0001701799, 0.0001997282, 0.0002275752, 0.000236969, 
    0.0002596506, 0.000249621, 0.0002544688, 0.0002670414, 0.0002719688, 
    0.0002558834, 0.0002441534, 0.0002689487, 0.000300166, 0.0002997848, 
    0.0002608746, 0.0001852801, 0.0001280596, 6.783474e-005, -1.578592e-005, 
    -8.8186e-005, -0.000126397, -0.0001405748, -0.0001443101, -0.000109501, 
    -5.31387e-005, 1.646345e-005, 6.815279e-005, 9.612716e-005, 0.0001192377, 
    0.0001562086, 0.0001983768, 0.0002383839, 0.000274067, 0.0003157589, 
    0.0003712308, 0.0004188349, 0.000452738, 0.0004789005, 0.0005262501, 
    0.000591927, 0.0006406754, 0.0006603687, 0.0006556797, 0.0006619107, 
    0.0006803484, 0.000669969, 0.0006279438, 0.0005679578, 0.0004988005, 
    0.0004360965, 0.0003672244, 0.0002958898, 0.0002794552, 0.0002848275, 
    0.0002559465, 0.0002189919, 0.0001924001, 0.0001866145, 0.000186678, 
    0.000187139, 0.0001923842, 0.0002081199, 0.000221662, 0.0002159716, 
    0.0001956744,
  0.0002500978, 0.0002309449, 0.0002211856, 0.0002287356, 0.0002568848, 
    0.0002790738, 0.000290486, 0.0003095276, 0.000318571, 0.0003417779, 
    0.0003722317, 0.0003891913, 0.0003814029, 0.0003883648, 0.0004214416, 
    0.0004466346, 0.0004532784, 0.0004559648, 0.000451816, 0.0004282126, 
    0.0004063894, 0.0003847571, 0.0003751088, 0.0003690054, 0.000362711, 
    0.0003701178, 0.0003606288, 0.0003417458, 0.0003295552, 0.0003264556, 
    0.0003046962, 0.0002505588, 0.0002117287, 0.0002069445, 0.0002051955, 
    0.0001997747, 0.000234155, 0.0003070161, 0.00037398, 0.000410283, 
    0.0004039411, 0.0004360643, 0.0005234205, 0.0005839942, 0.0006094095, 
    0.0006027026, 0.000504347, 0.0003235145, 0.0001581949, 6.671995e-006, 
    -0.0001149382, -0.0001592357, -0.0001703142, -0.0001876396, 
    -0.0001974301, -0.0001784363, -0.0001450572, -0.0001323577, 
    -0.0001107254, 1.843367e-005, 0.0001812894, 0.0002827449, 0.0003441134, 
    0.0004162272, 0.0004932843, 0.0005442579, 0.0005919258, 0.0006412943, 
    0.0006862762, 0.0007269657, 0.0007652561, 0.0007960438, 0.0008120975, 
    0.0008147042, 0.0008044681, 0.0007546856, 0.0006552967, 0.0006373045, 
    0.0006505447, 0.000674244, 0.0006684582, 0.0005853144, 0.00047054, 
    0.0003718345, 0.0003333539, 0.000317205, 0.0003180155, 0.000326074, 
    0.0003111488, 0.0002869572, 0.0002971459, 0.0003150904, 0.0003232602, 
    0.0002949683, 0.000270443, 0.0002638784,
  0.0004181513, 0.0004284829, 0.0004682827, 0.0005057622, 0.0005063666, 
    0.0005081622, 0.0005165229, 0.0005214503, 0.0005299696, 0.0005430509, 
    0.0005607414, 0.0005703897, 0.0005629989, 0.0005710884, 0.0006237472, 
    0.0006768666, 0.000705509, 0.0007432899, 0.0007187012, 0.0005725985, 
    0.0004776604, 0.0004592547, 0.0004531667, 0.0004519746, 0.000480664, 
    0.0005304939, 0.000558516, 0.0005707708, 0.0005876506, 0.0006124144, 
    0.0006028772, 0.0005515218, 0.0005187625, 0.0004940308, 0.0004501459, 
    0.0004234426, 0.0004633539, 0.0005310331, 0.0005706423, 0.0005675587, 
    0.0005682902, 0.0006416752, 0.0007184143, 0.0007178262, 0.0007178257, 
    0.0007303027, 0.0006848923, 0.0005364213, 0.0004229024, 0.0003619147, 
    0.0002894993, 0.0002486347, 0.000195038, 0.0001363391, 7.752934e-005, 
    3.960496e-005, 2.771569e-005, 2.733432e-005, 3.532926e-005, 0.0001211124, 
    0.0002545947, 0.0003446853, 0.0004161154, 0.0005196366, 0.0006031943, 
    0.0006133192, 0.0006321706, 0.0006854804, 0.0007270291, 0.0007419223, 
    0.0007535252, 0.0007474222, 0.0007433686, 0.0007378692, 0.0006948109, 
    0.0005785897, 0.0005781925, 0.0006279103, 0.0007154574, 0.0007754122, 
    0.0007800055, 0.0006980849, 0.0005378048, 0.0004364611, 0.0004179762, 
    0.0004147179, 0.0004499876, 0.0004686327, 0.0004520705, 0.0004480332, 
    0.0004499725, 0.0004634988, 0.0004515299, 0.0004101088, 0.0004021931, 
    0.0004173566,
  0.0005890485, 0.0006399597, 0.0007176842, 0.0007731873, 0.0008085854, 
    0.0008416777, 0.000861085, 0.0008693342, 0.000863723, 0.0008762958, 
    0.0009074653, 0.0009105015, 0.0009124405, 0.0009254259, 0.0009370614, 
    0.000953496, 0.0009809458, 0.001043777, 0.00104338, 0.0009305598, 
    0.0008561728, 0.000864327, 0.0008545835, 0.0008351761, 0.0008459683, 
    0.0009251391, 0.0009933906, 0.0009861905, 0.000967768, 0.0009803567, 
    0.0009961878, 0.0009739669, 0.0009056842, 0.0008078841, 0.0007345309, 
    0.0006998964, 0.0006922833, 0.0006758799, 0.000645394, 0.0006748941, 
    0.0007544947, 0.0008158158, 0.0008015265, 0.0007751891, 0.0008131294, 
    0.0008649454, 0.0008446961, 0.0007868716, 0.000740984, 0.0007272828, 
    0.0007391721, 0.0007258365, 0.0006481917, 0.0005736779, 0.0005347519, 
    0.0004786919, 0.0004419596, 0.0004093279, 0.0003721504, 0.0004025567, 
    0.0005026129, 0.000586187, 0.0006394815, 0.0006698873, 0.0006860681, 
    0.0006959229, 0.0007105777, 0.0007196693, 0.000713137, 0.0007228963, 
    0.0007451964, 0.0007406501, 0.0007088454, 0.0006675352, 0.000625208, 
    0.0006464436, 0.0006289911, 0.0006788042, 0.0008152276, 0.0008709221, 
    0.0008193124, 0.0007354217, 0.0006291028, 0.0005580536, 0.0005566869, 
    0.0006222995, 0.0007161736, 0.0007671793, 0.000754416, 0.0007349928, 
    0.0007049046, 0.0006557745, 0.0006179293, 0.0005937861, 0.000585394, 
    0.0005812924,
  0.0007884302, 0.0008868491, 0.0009362651, 0.0009514447, 0.001003181, 
    0.0010824, 0.001170027, 0.001236545, 0.001269082, 0.001282147, 
    0.001318434, 0.001334091, 0.001303303, 0.001255174, 0.001213959, 
    0.001175749, 0.001184506, 0.001200576, 0.001217504, 0.001250565, 
    0.001350319, 0.001409557, 0.001422925, 0.001362366, 0.00132929, 
    0.001322789, 0.001281686, 0.001214801, 0.001175128, 0.001178943, 
    0.001169962, 0.001125188, 0.001029693, 0.0009656218, 0.0009383629, 
    0.00091975, 0.0008850847, 0.0008215061, 0.0007440196, 0.0007477393, 
    0.0008697775, 0.0009475346, 0.0009810235, 0.001002561, 0.001110008, 
    0.001157677, 0.001152686, 0.001133198, 0.001111089, 0.001115254, 
    0.001179548, 0.001204501, 0.001112456, 0.0009993184, 0.0009369645, 
    0.0008830498, 0.0008558538, 0.0008537406, 0.0008397056, 0.0008109994, 
    0.0007871576, 0.0007727575, 0.0007982044, 0.0007842812, 0.0007744418, 
    0.000809506, 0.0008111112, 0.0007874593, 0.000772757, 0.0007483908, 
    0.0007217671, 0.000709306, 0.0007160613, 0.0006929035, 0.0006770398, 
    0.0006786617, 0.0007190178, 0.0007516178, 0.0005713576, 0.0008613542, 
    0.0008349526, 0.0007856959, 0.0008008587, 0.0008357633, 0.0008702385, 
    0.0009032357, 0.0009206561, 0.0009174929, 0.000926204, 0.0009248848, 
    0.0009005498, 0.000841279, 0.0007722331, 0.0007428443, 0.000735342, 
    0.0007302873,
  0.001009888, 0.00107237, 0.001140812, 0.001227119, 0.001328082, 0.00146967, 
    0.001697154, 0.001912064, 0.002053573, 0.00214802, 0.002204048, 
    0.002166966, 0.001989074, 0.00180449, 0.001678319, 0.001589325, 0.001572, 
    0.001564498, 0.00154339, 0.001556646, 0.001525047, 0.001474662, 
    0.001401007, 0.001280191, 0.001199209, 0.001189847, 0.00116254, 
    0.00115774, 0.001182155, 0.001169614, 0.001141082, 0.001129781, 
    0.001126825, 0.001119053, 0.001073102, 0.001017169, 0.0009804834, 
    0.0009256164, 0.0009132493, 0.0009675296, 0.001128224, 0.001192659, 
    0.001239294, 0.001313807, 0.001408269, 0.001460498, 0.001418887, 
    0.001415851, 0.001582664, 0.001658147, 0.001707723, 0.00171238, 
    0.001581727, 0.001401323, 0.001274198, 0.001192023, 0.001155529, 
    0.00114728, 0.001111518, 0.001080127, 0.001051755, 0.001021603, 
    0.001050498, 0.00104643, 0.001021841, 0.001029185, 0.0009972854, 
    0.0009635873, 0.000941447, 0.0009060334, 0.0008830028, 0.0008796807, 
    0.0008694604, 0.0008319337, 0.0007665111, 0.0006781053, 0.0007483596, 
    0.0007468811, 0.0004668823, 0.0009352323, 0.0008978955, 0.0009052539, 
    0.001027421, 0.001170487, 0.001191278, 0.001115301, 0.001033555, 
    0.0009972835, 0.001029503, 0.001053344, 0.001042154, 0.001005994, 
    0.0009805788, 0.0009720121, 0.0009642229, 0.0009578657,
  0.001140525, 0.001196967, 0.001263946, 0.001298374, 0.001364639, 
    0.00163766, 0.00183957, 0.002074508, 0.002307902, 0.002414444, 
    0.002302164, 0.002095344, 0.001866257, 0.001675443, 0.001572367, 
    0.001472453, 0.001387496, 0.001347234, 0.001266014, 0.001201561, 
    0.001153814, 0.001145136, 0.001141734, 0.001056411, 0.0009938981, 
    0.00102049, 0.001041598, 0.001057016, 0.001091968, 0.001153433, 
    0.001239009, 0.001259163, 0.001246337, 0.001155054, 0.001092493, 
    0.001116445, 0.001136536, 0.001132913, 0.001048957, 0.001500283, 
    0.001345773, 0.001705149, 0.001825423, 0.001799896, 0.001791473, 
    0.001781126, 0.001745569, 0.001738337, 0.001758507, 0.001725765, 
    0.001612707, 0.001565244, 0.001520645, 0.001427726, 0.001331452, 
    0.001281925, 0.001272022, 0.001290047, 0.001249006, 0.001241743, 
    0.001247877, 0.001212973, 0.001200957, 0.00118894, 0.001195887, 
    0.001194727, 0.00116858, 0.001182265, 0.001179086, 0.001141782, 
    0.001125824, 0.001071114, 0.0009273635, 0.0008307574, 0.0007790988, 
    0.000718113, 0.0007927688, 0.0009823591, 0.001252105, 0.001617904, 
    0.0011654, 0.001138252, 0.00134733, 0.001483674, 0.001418792, 
    0.001286835, 0.001238261, 0.001228263, 0.001240645, 0.001202784, 
    0.001137727, 0.001117764, 0.00107496, 0.001025385, 0.001014593, 
    0.001064835,
  0.001293671, 0.001262327, 0.001233955, 0.001283389, 0.001550321, 
    0.001781031, 0.002056864, 0.002315772, 0.002463814, 0.002401983, 
    0.001988025, 0.001753659, 0.001637661, 0.001565533, 0.001544503, 
    0.001447816, 0.00130359, 0.001227947, 0.001178801, 0.001175289, 
    0.00118039, 0.001171489, 0.001145137, 0.001102109, 0.001097548, 
    0.001157375, 0.001205027, 0.001262233, 0.0013051, 0.001482944, 
    0.001559333, 0.001550814, 0.001530342, 0.001403041, 0.00133239, 
    0.001335092, 0.001143673, 0.001675299, 0.001785909, 0.002026442, 
    0.002072298, 0.002344556, 0.002498829, 0.002192843, 0.002052558, 
    0.002000009, 0.001863395, 0.001743041, 0.001591915, 0.001488077, 
    0.001403423, 0.001357885, 0.00134021, 0.001282704, 0.001263201, 
    0.001295722, 0.001325318, 0.001327209, 0.001325969, 0.001339098, 
    0.001357329, 0.00135825, 0.001385367, 0.001401849, 0.001407429, 
    0.001399959, 0.001342945, 0.001280717, 0.001241998, 0.001183219, 
    0.001110089, 0.0009923903, 0.000915492, 0.0008411687, 0.0007245811, 
    0.000784169, 0.0009160312, 0.002077575, 0.002155266, 0.001658784, 
    0.001492099, 0.001776484, 0.00170383, 0.001908202, 0.001884616, 
    0.001689207, 0.001646451, 0.001592839, 0.001507613, 0.001426916, 
    0.001350462, 0.001329418, 0.001275027, 0.001242697, 0.001248674, 
    0.001272801,
  0.001283322, 0.001253347, 0.00121973, 0.001422608, 0.001694723, 
    0.001599942, 0.00223431, 0.003559443, 0.003179912, 0.002604117, 
    0.002328042, 0.002251511, 0.002235393, 0.002166505, 0.002063365, 
    0.001977345, 0.001911096, 0.001910143, 0.001871264, 0.001869039, 
    0.001858452, 0.001771653, 0.001746841, 0.001692371, 0.001689191, 
    0.001663441, 0.001672137, 0.001765547, 0.001732694, 0.001734601, 
    0.001832306, 0.002439241, 0.001863858, 0.001532471, 0.001414405, 
    0.001435132, 0.0016736, 0.001665937, 0.001709138, 0.002292549, 
    0.002722148, 0.002085459, 0.001709346, 0.001600325, 0.001747429, 
    0.00181355, 0.001754645, 0.001602678, 0.001586148, 0.001607143, 
    0.001579392, 0.00159872, 0.001608209, 0.001552355, 0.001485836, 
    0.001496756, 0.001488411, 0.001398909, 0.001371585, 0.001415438, 
    0.001458927, 0.001489588, 0.001491114, 0.001464681, 0.001446735, 
    0.001417284, 0.001375862, 0.001198795, 0.001111757, 0.001070558, 
    0.0009265859, 0.0008801743, 0.0008761203, 0.0008032126, 0.0006517535, 
    0.0007889243, 0.0009815022, 0.001593745, 0.001995162, 0.002104389, 
    0.00222139, 0.002696336, 0.002652913, 0.002391478, 0.00242775, 
    0.002244261, 0.002187042, 0.00206904, 0.001915467, 0.001820736, 
    0.001687475, 0.00157324, 0.001482817, 0.001450518, 0.001434227, 
    0.001360825,
  0.001312729, 0.00126808, 0.001333692, 0.001544788, 0.002055594, 
    0.002320301, 0.003324742, 0.003673295, 0.003108721, 0.002624207, 
    0.002652245, 0.002721943, 0.002746292, 0.002753939, 0.002691377, 
    0.00261324, 0.002605515, 0.002573916, 0.002461192, 0.002345703, 
    0.002228001, 0.002129725, 0.002103881, 0.002011262, 0.001914719, 
    0.001858898, 0.00180039, 0.001793762, 0.00177658, 0.001990329, 
    0.002443246, 0.003153862, 0.00267672, 0.001318354, 0.0007586442, 
    0.001156754, 0.001468335, 0.001647101, 0.002077352, 0.00260103, 
    0.002789368, 0.001765072, 0.00141444, 0.001577405, 0.001804475, 
    0.001974356, 0.002086715, 0.002141074, 0.002158526, 0.002154283, 
    0.002140708, 0.002084823, 0.001993493, 0.001897649, 0.001751244, 
    0.001574195, 0.001489651, 0.00143542, 0.001441189, 0.001489604, 
    0.00151203, 0.001526447, 0.001489222, 0.001480942, 0.001473105, 
    0.001368439, 0.001263424, 0.001108532, 0.001020078, 0.0009266008, 
    0.0008346038, 0.0008990243, 0.0007925155, 0.0008123359, 0.0007854262, 
    0.0008692071, 0.001162779, 0.0009225802, 0.002530299, 0.00263004, 
    0.002753317, 0.003310472, 0.003526096, 0.003364114, 0.003110868, 
    0.002856172, 0.002668712, 0.0023701, 0.002141981, 0.001965854, 
    0.001809498, 0.001711937, 0.00162938, 0.00154738, 0.00149275, 0.001388753,
  0.001457321, 0.001471451, 0.001717739, 0.00203485, 0.002425841, 
    0.003789596, 0.003869403, 0.003686059, 0.003129859, 0.00288286, 
    0.002966335, 0.003061544, 0.003293812, 0.002874514, 0.002717968, 
    0.00278274, 0.002671413, 0.002542778, 0.00242794, 0.002326087, 
    0.002241846, 0.0021845, 0.00214098, 0.002068994, 0.001970176, 
    0.001965185, 0.001903149, 0.001937703, 0.002022945, 0.002321416, 
    0.002720989, 0.002917953, 0.002063443, 0.0004582852, 0.0005431941, 
    0.001305496, 0.001346106, 0.001811053, 0.002380827, 0.002836431, 
    0.002314119, 0.001731314, 0.001875445, 0.002177935, 0.002343716, 
    0.002445757, 0.002594722, 0.002645633, 0.002622347, 0.002564841, 
    0.002539743, 0.002477102, 0.002321463, 0.002125245, 0.001931951, 
    0.001743743, 0.001662252, 0.001684742, 0.001708202, 0.001696965, 
    0.001728659, 0.001755807, 0.001715706, 0.001599562, 0.001491115, 
    0.001359634, 0.001215232, 0.00109316, 0.001016263, 0.0009588357, 
    0.0009977147, 0.001005804, 0.0008564582, 0.0009270934, 0.0008525336, 
    0.00117578, 0.001964422, 0.0008909665, 0.002385707, 0.003196792, 
    0.003356088, 0.003516415, 0.003794763, 0.003612451, 0.003408873, 
    0.002991196, 0.002645615, 0.002328791, 0.002094584, 0.00192723, 
    0.001799566, 0.001695439, 0.001662521, 0.001613517, 0.001575943, 
    0.001489746,
  0.001822356, 0.001846961, 0.002032816, 0.0022493, 0.002932131, 0.003883406, 
    0.0039501, 0.003693848, 0.003366341, 0.003029392, 0.002993912, 
    0.003342113, 0.003106004, 0.002855966, 0.002728697, 0.00273747, 
    0.002631215, 0.002598885, 0.002514059, 0.002454231, 0.002459761, 
    0.002434457, 0.002335688, 0.002290579, 0.002240209, 0.002239923, 
    0.002215335, 0.00226499, 0.002424777, 0.002646476, 0.002976285, 
    0.002873864, 0.002235964, 0.0001784291, 0.0006851628, 0.001281733, 
    0.001535904, 0.002421153, 0.002707288, 0.002507398, 0.002021883, 
    0.002229799, 0.002468774, 0.002596581, 0.002804119, 0.002870765, 
    0.002977367, 0.003018597, 0.003008172, 0.002996234, 0.002969865, 
    0.00283961, 0.002632629, 0.00240138, 0.00225294, 0.002231261, 
    0.002223598, 0.00220214, 0.002187835, 0.002207624, 0.002263637, 
    0.002234327, 0.00218275, 0.002019307, 0.001817096, 0.001670468, 
    0.001511269, 0.00143596, 0.001393314, 0.00139368, 0.001327082, 
    0.001284356, 0.001268303, 0.001265219, 0.001235083, 0.001725541, 
    0.002395753, 0.001354054, 0.002907764, 0.003476268, 0.003763516, 
    0.003595542, 0.003486803, 0.003290365, 0.00312611, 0.003196759, 
    0.002395038, 0.002348896, 0.002209025, 0.002080326, 0.002003016, 
    0.001877051, 0.001823947, 0.001775309, 0.001775007, 0.001790566,
  0.002205831, 0.00229263, 0.002412125, 0.002648588, 0.003147616, 
    0.003755821, 0.00371292, 0.003515082, 0.003446259, 0.002890631, 
    0.002652563, 0.003212288, 0.003101965, 0.002997873, 0.002902491, 
    0.002888663, 0.002819965, 0.00281572, 0.002796931, 0.00279423, 
    0.002752047, 0.002737438, 0.002705492, 0.002706159, 0.002645362, 
    0.002630072, 0.002733449, 0.002831042, 0.002950361, 0.002971012, 
    0.00310945, 0.003341781, 0.003440676, 0.003246067, 0.003115207, 
    0.002492249, 0.002213633, 0.002846032, 0.003034778, 0.002384596, 
    0.00252164, 0.002748452, 0.0028481, 0.002892286, 0.003045158, 
    0.003133772, 0.003278714, 0.003324777, 0.00335359, 0.003323739, 
    0.00331635, 0.00318196, 0.003086021, 0.003046904, 0.002997074, 0.0029801, 
    0.002916584, 0.002890343, 0.002878167, 0.002892541, 0.002873927, 
    0.002782244, 0.002671588, 0.002521336, 0.002318634, 0.002203333, 
    0.002070344, 0.001993813, 0.00196312, 0.001919678, 0.001884536, 
    0.001904818, 0.001837282, 0.001796624, 0.001776738, 0.002128422, 
    0.002142965, 0.002396038, 0.002703995, 0.003728736, 0.003835725, 
    0.003597064, 0.003407124, 0.003146121, 0.003066552, 0.002798427, 
    0.002516536, 0.002462685, 0.002368655, 0.002290279, 0.002281106, 
    0.002208882, 0.002200744, 0.002167366, 0.002208724, 0.002194656,
  0.002630771, 0.002686244, 0.002908386, 0.002944561, 0.002896941, 
    0.003121245, 0.003150381, 0.003138443, 0.003216455, 0.002803179, 
    0.002633536, 0.00302365, 0.00312876, 0.003037335, 0.003078168, 
    0.003104204, 0.003084973, 0.003038418, 0.003078105, 0.003113585, 
    0.003057636, 0.003035225, 0.003027596, 0.002999589, 0.003018565, 
    0.003072688, 0.003166912, 0.003209718, 0.003285244, 0.003306573, 
    0.003305683, 0.003331337, 0.003569201, 0.003488917, 0.003478251, 
    0.003511744, 0.003324062, 0.003216324, 0.002927905, 0.002621278, 
    0.002815733, 0.00294343, 0.002920574, 0.00302268, 0.003168434, 
    0.003313884, 0.003387541, 0.003257919, 0.003249496, 0.003209809, 
    0.003226068, 0.003257174, 0.003272781, 0.003317669, 0.003353573, 
    0.003330734, 0.003370898, 0.003451563, 0.003449896, 0.003328094, 
    0.003187479, 0.003060417, 0.002964476, 0.002919225, 0.002781944, 
    0.002659412, 0.002533544, 0.002445488, 0.002476736, 0.002465563, 
    0.002445171, 0.002385455, 0.002340393, 0.002376966, 0.002327105, 
    0.002922244, 0.00340064, 0.002905888, 0.002921627, 0.003760222, 
    0.00358942, 0.003101345, 0.003209524, 0.003199223, 0.002744179, 
    0.002334513, 0.002658347, 0.002707096, 0.002753332, 0.002695858, 
    0.002671858, 0.002632074, 0.002620392, 0.002603767, 0.00260817, 0.00262249,
  0.003075087, 0.003000304, 0.003143562, 0.003023066, 0.002749377, 
    0.002814783, 0.002788557, 0.002712135, 0.002978878, 0.0029846, 
    0.002952477, 0.003150599, 0.003108099, 0.003153827, 0.003163379, 
    0.00320817, 0.003203005, 0.003187746, 0.003179511, 0.003118971, 
    0.0031489, 0.003189383, 0.003285928, 0.003248796, 0.003229247, 
    0.003228515, 0.003215879, 0.003285116, 0.00334294, 0.003299564, 
    0.003361568, 0.003209123, 0.003215991, 0.003307987, 0.003300408, 
    0.003272973, 0.003150966, 0.003104156, 0.002902219, 0.002771864, 
    0.003027068, 0.003149265, 0.002935467, 0.003026066, 0.003112406, 
    0.003125917, 0.003127791, 0.003067663, 0.003079392, 0.00310743, 
    0.003175665, 0.003388733, 0.003416963, 0.00346552, 0.003565639, 
    0.00360962, 0.003662277, 0.003677743, 0.003646161, 0.003541671, 
    0.003435956, 0.003317624, 0.003268398, 0.003232047, 0.003153941, 
    0.003027627, 0.002978355, 0.002951508, 0.002935374, 0.002960345, 
    0.002940874, 0.002912804, 0.0029767, 0.002996903, 0.002962237, 
    0.003068428, 0.00265741, 0.002732655, 0.002950108, 0.003472358, 
    0.003241343, 0.002934404, 0.002695223, 0.003115125, 0.003018646, 
    0.002898404, 0.002648684, 0.00302526, 0.003084594, 0.002999095, 
    0.00302971, 0.003038451, 0.003033603, 0.003050055, 0.00302672, 0.003019568,
  0.003484992, 0.003387367, 0.003338143, 0.003179945, 0.003024828, 
    0.002973378, 0.002922785, 0.002762315, 0.002814448, 0.002970024, 
    0.003246686, 0.003244489, 0.003157292, 0.003104428, 0.00316675, 
    0.003350664, 0.003295273, 0.003213432, 0.003227182, 0.003193595, 
    0.003217278, 0.003225129, 0.003352571, 0.003388669, 0.00340604, 
    0.0033678, 0.003343973, 0.003346486, 0.003147982, 0.003436847, 
    0.003329206, 0.003286213, 0.003281048, 0.003309624, 0.003250515, 
    0.003178542, 0.003062941, 0.002632964, 0.00253631, 0.002793087, 
    0.003073813, 0.003195122, 0.003090566, 0.003159294, 0.003108941, 
    0.003152221, 0.003272209, 0.003488677, 0.003653917, 0.003811417, 
    0.00390467, 0.004130295, 0.004158951, 0.004290288, 0.004395733, 
    0.004408274, 0.004404729, 0.004328929, 0.00430407, 0.004230781, 
    0.004155999, 0.004028415, 0.003932744, 0.003785986, 0.003656145, 
    0.003550446, 0.003476171, 0.003424147, 0.003339734, 0.003375813, 
    0.003348252, 0.003378898, 0.003300281, 0.003183169, 0.003358329, 
    0.003352687, 0.002390826, 0.003712986, 0.003849883, 0.003242301, 
    0.002819519, 0.002342299, 0.00217161, 0.002312672, 0.003236689, 
    0.003064105, 0.003114982, 0.003198966, 0.003272908, 0.003295245, 
    0.003327496, 0.003331689, 0.003341336, 0.003421558, 0.003421001, 
    0.003392026,
  0.003357742, 0.003301647, 0.003316527, 0.003004229, 0.002799317, 
    0.002568847, 0.002395818, 0.00227249, 0.002556337, 0.002974617, 
    0.003179326, 0.003682023, 0.003299484, 0.003147025, 0.003058413, 
    0.003126249, 0.003190972, 0.003152175, 0.003225876, 0.003258731, 
    0.00317147, 0.003216721, 0.003305208, 0.003371695, 0.003452104, 
    0.003369087, 0.003287213, 0.002843853, 0.002696525, 0.003256505, 
    0.003033681, 0.002735054, 0.002587173, 0.002993276, 0.003192419, 
    0.002998589, 0.002823507, 0.002868712, 0.002957484, 0.003058983, 
    0.003135627, 0.003188301, 0.003283605, 0.003323199, 0.003324851, 
    0.003626611, 0.003875569, 0.004194811, 0.004230207, 0.004297489, 
    0.004393397, 0.004448932, 0.004392253, 0.004416322, 0.004388187, 
    0.004394321, 0.004379937, 0.004284028, 0.004223535, 0.004147066, 
    0.004076891, 0.003991775, 0.00392694, 0.003865922, 0.003789134, 
    0.003749257, 0.003688633, 0.003636595, 0.00357502, 0.003540734, 
    0.00346452, 0.003469398, 0.003409827, 0.003339652, 0.003167279, 
    0.003389817, 0.0034533, 0.004468773, 0.004072806, 0.002722532, 
    0.002030417, 0.001553563, 0.001610227, 0.001988885, 0.002586966, 
    0.003181133, 0.003184296, 0.00321928, 0.003272258, 0.003261214, 
    0.00330211, 0.003342737, 0.003350288, 0.003375402, 0.003341451, 
    0.003352974,
  0.003178272, 0.003356451, 0.00327442, 0.002596693, 0.002093631, 
    0.002307142, 0.002221183, 0.002234805, 0.002694223, 0.003307291, 
    0.003230648, 0.003557362, 0.003601896, 0.00338568, 0.003389066, 
    0.003162203, 0.003181119, 0.003094969, 0.003073178, 0.003067726, 
    0.003012571, 0.003035858, 0.003069172, 0.003170675, 0.003306318, 
    0.003323041, 0.00316551, 0.002614273, 0.002847252, 0.002971627, 
    0.002901947, 0.002463497, 0.002454389, 0.002852131, 0.002849923, 
    0.002882699, 0.002917126, 0.003047206, 0.003121609, 0.003071159, 
    0.002992401, 0.003008805, 0.002997058, 0.002986234, 0.003079806, 
    0.003321227, 0.003543753, 0.003866477, 0.003953228, 0.004079623, 
    0.004167853, 0.004179949, 0.004214155, 0.004243547, 0.004248427, 
    0.004315391, 0.004377456, 0.004409563, 0.004390966, 0.004332079, 
    0.004175436, 0.004059708, 0.003884202, 0.003760271, 0.003670434, 
    0.003609637, 0.003550032, 0.003503112, 0.003484771, 0.003537126, 
    0.003550114, 0.00353023, 0.003295911, 0.00315389, 0.002849212, 
    0.003231984, 0.003302682, 0.003218552, 0.003430618, 0.002139771, 
    0.00193203, 0.001488522, 0.002134304, 0.003002701, 0.002860921, 
    0.002846712, 0.002822075, 0.002940729, 0.002963027, 0.002986271, 
    0.003090678, 0.003079126, 0.003088932, 0.003190227, 0.003231678, 
    0.003225114,
  0.002864151, 0.002989622, 0.001684233, 0.00189296, 0.001842272, 
    0.002297619, 0.002452306, 0.002251351, 0.002640371, 0.003152924, 
    0.003188114, 0.003136854, 0.003252408, 0.003193136, 0.003376355, 
    0.003477918, 0.003527714, 0.003415389, 0.003334103, 0.003248256, 
    0.0032453, 0.00327073, 0.003197188, 0.003159678, 0.00320245, 0.003422827, 
    0.003222685, 0.002753588, 0.003132544, 0.002937136, 0.002792321, 
    0.002707047, 0.002915312, 0.00308691, 0.002924994, 0.002976364, 
    0.003011793, 0.003029117, 0.003065597, 0.003070109, 0.003038146, 
    0.003048526, 0.00296344, 0.0029334, 0.002933733, 0.002992036, 
    0.003063865, 0.003130795, 0.003230708, 0.0033901, 0.003456555, 
    0.003515951, 0.003569152, 0.003639471, 0.003667347, 0.003681924, 
    0.003682829, 0.00368976, 0.003598016, 0.003589768, 0.00349912, 
    0.003532674, 0.003533613, 0.003541242, 0.003572935, 0.003565671, 
    0.003560411, 0.003579807, 0.003566947, 0.003610101, 0.003499839, 
    0.003504751, 0.003433635, 0.003410334, 0.003384363, 0.003569648, 
    0.003234287, 0.002966607, 0.003282862, 0.00137459, 0.002022883, 
    0.002666995, 0.002870221, 0.002899995, 0.002772389, 0.002746847, 
    0.002731778, 0.002776457, 0.002769325, 0.002878536, 0.002930066, 
    0.002994105, 0.003132723, 0.003022365, 0.002234931, 0.002607469,
  0.00174393, 0.001678113, 0.00158473, 0.00175253, 0.001821115, 0.001896187, 
    0.001728149, 0.001747985, 0.002342109, 0.002882302, 0.00331371, 
    0.003159327, 0.002996266, 0.002969499, 0.003289664, 0.003515033, 
    0.003529642, 0.003597444, 0.003679015, 0.003690844, 0.003388163, 
    0.003081352, 0.003166273, 0.003119722, 0.00303923, 0.00316661, 
    0.003180293, 0.00337691, 0.003020536, 0.002850974, 0.002860429, 
    0.002913246, 0.002842087, 0.002717428, 0.002817927, 0.002972852, 
    0.003020804, 0.003017992, 0.002985995, 0.003014734, 0.002979672, 
    0.002950249, 0.002933957, 0.002961423, 0.002952188, 0.00297638, 
    0.002986217, 0.002951473, 0.002969021, 0.002991481, 0.002995484, 
    0.003076309, 0.00307712, 0.003086513, 0.003062846, 0.003038384, 
    0.002966447, 0.002921702, 0.002837254, 0.002805816, 0.002800617, 
    0.002882062, 0.003005913, 0.003138632, 0.003237622, 0.003307352, 
    0.003328048, 0.003482495, 0.003510358, 0.003561253, 0.003626404, 
    0.003614631, 0.003376558, 0.003319247, 0.003272132, 0.003376577, 
    0.003079523, 0.003013353, 0.003051247, 0.002872463, 0.002888899, 
    0.002678296, 0.002850974, 0.002777349, 0.002657996, 0.002687387, 
    0.002769498, 0.002879394, 0.003003674, 0.003056632, 0.003079442, 
    0.003245605, 0.003053186, 0.002456263, 0.001847231, 0.001675664,
  0.002030812, 0.001799419, 0.00162051, 0.001630667, 0.001657386, 
    0.001724301, 0.001578199, 0.001714082, 0.00203563, 0.00326509, 
    0.003339539, 0.002539932, 0.002278958, 0.002356063, 0.002949123, 
    0.003200846, 0.003321756, 0.003434272, 0.00348644, 0.003667828, 
    0.003037497, 0.002714233, 0.003173253, 0.003120385, 0.002936821, 
    0.002864772, 0.002799588, 0.003024399, 0.002538041, 0.00236255, 
    0.002605483, 0.002825368, 0.002725789, 0.00267313, 0.002824714, 
    0.002954811, 0.002952507, 0.002996026, 0.002942905, 0.003013413, 
    0.002967542, 0.002922544, 0.002913723, 0.00294343, 0.002957338, 
    0.002967145, 0.002967482, 0.00301178, 0.003062008, 0.003105208, 
    0.003066154, 0.003075102, 0.003104048, 0.003106717, 0.003065787, 
    0.003045268, 0.002992578, 0.00297457, 0.002925217, 0.002842963, 
    0.00283527, 0.002810586, 0.002827244, 0.002914552, 0.002999587, 
    0.003087614, 0.00306347, 0.003237719, 0.003263071, 0.003132278, 
    0.003318671, 0.003283959, 0.002893222, 0.002609011, 0.003084194, 
    0.003205167, 0.003059272, 0.002910482, 0.002853787, 0.002778383, 
    0.002842646, 0.002710275, 0.00271444, 0.002485098, 0.002509354, 
    0.002480758, 0.00256899, 0.002686594, 0.002833458, 0.0028827, 
    0.003047765, 0.002938713, 0.002194288, 0.002042447, 0.00202455, 
    0.001690828,
  0.001173413, 0.001062485, 0.0009979848, 0.0009114069, 0.0008133692, 
    0.0009311964, 0.000933151, 0.0008531378, 0.0007699132, 0.001787529, 
    0.003393487, 0.002916616, 0.001894756, 0.001262995, 0.001631001, 
    0.002730827, 0.003095003, 0.003084132, 0.003090935, 0.003177036, 
    0.002551646, 0.002446298, 0.002995456, 0.002940541, 0.002797648, 
    0.002656075, 0.002718825, 0.002432006, 0.002189855, 0.002273079, 
    0.002538536, 0.002628639, 0.002651036, 0.002555098, 0.002689693, 
    0.002737759, 0.002765251, 0.002875164, 0.00290565, 0.002920548, 
    0.00291921, 0.002939573, 0.002901537, 0.002890823, 0.002839593, 
    0.002836542, 0.00282702, 0.002869746, 0.002861766, 0.002909593, 
    0.002911899, 0.002894271, 0.002870429, 0.002790956, 0.00277468, 
    0.002726169, 0.002670952, 0.002556622, 0.002461939, 0.002403812, 
    0.002345081, 0.002328075, 0.00233386, 0.002382911, 0.002453357, 
    0.002535483, 0.002523959, 0.002522275, 0.002512166, 0.001686092, 
    0.001708185, 0.00173918, 0.001867275, 0.002869252, 0.003261292, 
    0.003158215, 0.003072083, 0.002983505, 0.002971502, 0.002841851, 
    0.002740333, 0.002583945, 0.002445122, 0.002342364, 0.002296, 
    0.002166713, 0.002341442, 0.002361278, 0.002497416, 0.002599299, 
    0.002803545, 0.002696224, 0.001667637, 0.001390151, 0.001150414, 
    0.0009805802,
  0.0008451112, 0.0008424409, 0.0007167461, 0.0009639552, 0.0006659946, 
    0.0008279763, 0.0008437913, 0.0008316957, 0.0006398798, 0.001113156, 
    0.002731924, 0.002108426, 0.001563625, 0.00100164, 0.001040153, 
    0.001925893, 0.002921212, 0.002822809, 0.002706571, 0.002502263, 
    0.002037011, 0.001717261, 0.001652759, 0.001947829, 0.002396468, 
    0.002098333, 0.001899602, 0.001962735, 0.001882007, 0.001941388, 
    0.002249332, 0.002317457, 0.00242357, 0.002444964, 0.002440004, 
    0.002529267, 0.002522735, 0.002534576, 0.00264563, 0.00268955, 
    0.002703996, 0.002683317, 0.00264816, 0.00271328, 0.002614222, 
    0.002557082, 0.002522703, 0.002538519, 0.002551585, 0.002569973, 
    0.002639083, 0.002658127, 0.002661798, 0.00267092, 0.002672702, 
    0.002565302, 0.00249473, 0.002402556, 0.002325294, 0.002288704, 
    0.002164328, 0.002064081, 0.001936877, 0.001883265, 0.001901177, 
    0.00197531, 0.001996594, 0.001794956, 0.0011476, 0.0009561181, 
    0.001023447, 0.001157057, 0.001545966, 0.002570864, 0.003024431, 
    0.003202625, 0.003261356, 0.003172966, 0.00303904, 0.002883717, 
    0.002727156, 0.00249899, 0.002368049, 0.002165411, 0.001986247, 
    0.001920251, 0.00197396, 0.001958255, 0.002132078, 0.002202603, 
    0.002374296, 0.002379078, 0.001167628, 0.0008435689, 0.0006245896, 
    0.0004640226,
  0.0007660361, 0.0006614807, 0.0006166261, 0.0005616627, 0.0006893917, 
    0.0009381101, 0.0008245432, 0.0009199744, 0.0007247091, 0.0008382597, 
    0.002033452, 0.001088059, 0.001068159, 0.001166944, 0.001036863, 
    0.001543216, 0.002625222, 0.002478294, 0.001738098, 0.001411196, 
    0.001272675, 0.001337142, 0.001138777, 0.001245908, 0.00166511, 
    0.001593871, 0.00132263, 0.001503415, 0.001403168, 0.001319071, 
    0.001495245, 0.001644431, 0.001956856, 0.0020901, 0.002134082, 
    0.002201108, 0.002211473, 0.0022092, 0.00227618, 0.002259219, 
    0.002212711, 0.002187995, 0.002159338, 0.002229322, 0.002212665, 
    0.00215929, 0.002067674, 0.002028018, 0.002023852, 0.002074811, 
    0.002213173, 0.002257027, 0.00228125, 0.002303501, 0.002329967, 
    0.002304805, 0.002277005, 0.002206147, 0.002105074, 0.002047662, 
    0.001987994, 0.001896711, 0.001772719, 0.001646593, 0.001569043, 
    0.001549684, 0.001492226, 0.0004371433, 0.0003589736, 0.0006990223, 
    0.0008873092, 0.001616362, 0.00172939, 0.002113832, 0.002594072, 
    0.002941845, 0.003072482, 0.003161683, 0.003119482, 0.002867315, 
    0.002716824, 0.00260507, 0.002402605, 0.002119126, 0.00207017, 
    0.001951325, 0.001860344, 0.001935112, 0.001950816, 0.001923111, 
    0.002080405, 0.002068658, 0.001064774, 0.0007883043, 0.0008962762, 
    0.0007169533,
  0.0005321624, 0.0007369167, 0.0006790287, 0.0006269903, 0.0009920239, 
    0.001162699, 0.0008135922, 0.0009381103, 0.001078761, 0.0006996912, 
    0.0006156089, 0.0004982275, 0.0007290004, 0.001063772, 0.00105759, 
    0.001024354, 0.001254093, 0.001291859, 0.001248865, 0.001048005, 
    0.0009358684, 0.0009211348, 0.0009773227, 0.0007173978, 0.0009838231, 
    0.001268081, 0.0009988281, 0.001041567, 0.001001068, 0.000815595, 
    0.0007804681, 0.000780134, 0.00117365, 0.001798879, 0.001879005, 
    0.001912892, 0.002018559, 0.002072727, 0.002072267, 0.00201813, 
    0.001931616, 0.00192041, 0.001887413, 0.001860361, 0.001833753, 
    0.001769793, 0.001662504, 0.001608226, 0.001589342, 0.001587196, 
    0.001703131, 0.001843575, 0.001941725, 0.001998468, 0.002061888, 
    0.002119951, 0.00209169, 0.002017796, 0.001978807, 0.001944267, 
    0.001894978, 0.001791934, 0.001678018, 0.001526797, 0.001411466, 
    0.001318498, 0.0005445755, 0.0002988768, 0.0002783095, 0.0005806559, 
    0.0007820241, 0.001488857, 0.001750068, 0.001938927, 0.001624564, 
    0.002328885, 0.002578352, 0.00273868, 0.002858635, 0.002785123, 
    0.002623968, 0.002412667, 0.002243705, 0.00211461, 0.001968745, 
    0.001743916, 0.001809211, 0.001922174, 0.001860805, 0.001836678, 
    0.001850219, 0.001885442, 0.001851887, 0.0009358204, 0.0005325768, 
    0.0003150268,
  0.0004151785, 0.0004201543, 0.0003876653, 0.0008267355, 0.001135598, 
    0.001539861, 0.001090172, 0.001166529, 0.001566263, 0.0008878824, 
    0.0003948978, 0.0003335285, 0.0006270371, 0.0008365435, 0.001035814, 
    0.001042299, 0.000989815, 0.001136649, 0.001275949, 0.0009302103, 
    0.0003118797, 0.0006199961, 0.0005563539, 0.0004340927, 0.0004556298, 
    0.0005675438, 0.0006016854, 0.0006844008, 0.0007611713, 0.0007952813, 
    0.0007589939, 0.0006903133, 0.0008613393, 0.001202975, 0.001404327, 
    0.001719233, 0.001881499, 0.001899604, 0.001928357, 0.001911636, 
    0.001802314, 0.00173999, 0.001698792, 0.001659437, 0.001628157, 
    0.001565627, 0.001509838, 0.001435038, 0.00138462, 0.001334234, 
    0.001337095, 0.001382394, 0.001504352, 0.001671595, 0.001806572, 
    0.001898125, 0.001877351, 0.001824692, 0.001801344, 0.001797434, 
    0.001735921, 0.001611467, 0.001478397, 0.001356136, 0.001269891, 
    0.0009581838, 0.000572233, 0.0003672568, 0.0004132395, 0.0005412698, 
    0.0005960581, 0.0007139319, 0.0006733686, 0.000805039, 0.001138094, 
    0.001912478, 0.002125593, 0.002178983, 0.002246217, 0.002272729, 
    0.002251399, 0.002187788, 0.002132046, 0.001990441, 0.001774164, 
    0.001646037, 0.001666176, 0.001696725, 0.001804999, 0.00185219, 
    0.001752658, 0.00172985, 0.001762577, 0.00161285, 0.0006161486, 
    0.0004179119,
  0.0005457201, 0.0007253443, 0.0009017899, 0.001606044, 0.001710044, 
    0.001611116, 0.001353434, 0.001271194, 0.001449261, 0.001469336, 
    0.0005823565, 0.0003714692, 0.0005309384, 0.000688422, 0.0008512307, 
    0.001044333, 0.0009791339, 0.001088902, 0.001099949, 0.0006542649, 
    0.0004426122, 0.0004952073, 0.0004853366, 0.0003707688, 0.0003675421, 
    0.0003954371, 0.0004820625, 0.0005706593, 0.0007117393, 0.0007391575, 
    0.0007699453, 0.0008404218, 0.0009234711, 0.001044841, 0.001066983, 
    0.001410447, 0.001211354, 0.001276108, 0.001625088, 0.001660262, 
    0.001570854, 0.001492399, 0.001418235, 0.001373016, 0.001313761, 
    0.001256652, 0.001256605, 0.001262613, 0.001280145, 0.001277093, 
    0.001259004, 0.001253217, 0.001291475, 0.001403136, 0.001549715, 
    0.001730374, 0.001784893, 0.001717404, 0.001681721, 0.001666208, 
    0.001590231, 0.00147981, 0.001320023, 0.001164066, 0.0008373219, 
    0.0005960432, 0.0004998331, 0.0005182864, 0.0004997216, 0.0003385511, 
    0.0005409531, 0.0006793467, 0.0007468662, 0.0007998268, 0.0008813818, 
    0.001152813, 0.001742708, 0.001930264, 0.001920759, 0.001896376, 
    0.001876476, 0.001753214, 0.001708758, 0.001688254, 0.001528434, 
    0.001349891, 0.001218172, 0.001308087, 0.001571667, 0.001659389, 
    0.001656719, 0.00159438, 0.00153735, 0.001751974, 0.001634958, 
    0.0008075191,
  0.001127286, 0.001597971, 0.001610687, 0.001625929, 0.001627773, 
    0.001480957, 0.0009961086, 0.0007496323, 0.0006360337, 0.0005823895, 
    0.0005214817, 0.0005813721, 0.0006691418, 0.0007673232, 0.00107903, 
    0.0009025065, 0.0009238683, 0.001020364, 0.001069431, 0.0006915855, 
    0.0004902323, 0.0003699899, 0.0002412918, 0.0002465051, 0.0003587683, 
    0.000384883, 0.0004771193, 0.0005490422, 0.0006903133, 0.0006595096, 
    0.000579258, 0.0006394027, 0.0007153476, 0.0006439646, 0.0007297482, 
    0.001129591, 0.001158535, 0.000953655, 0.001234496, 0.001311933, 
    0.001333677, 0.001300203, 0.001233891, 0.001219458, 0.001188972, 
    0.001119132, 0.001088773, 0.001080667, 0.001091666, 0.00108925, 
    0.001103364, 0.001140907, 0.001162651, 0.001207617, 0.001277267, 
    0.001375051, 0.001496405, 0.001552656, 0.001553182, 0.001491716, 
    0.001391946, 0.001276807, 0.001125267, 0.0008418988, 0.0006755958, 
    0.0006433448, 0.0006683788, 0.0005860131, 0.0005595966, 0.0005689743, 
    0.0005248508, 0.0005848052, 0.0006857049, 0.0006711297, 0.00065293, 
    0.000829821, 0.001186765, 0.001781395, 0.001900238, 0.001910538, 
    0.001830939, 0.001536046, 0.001340734, 0.00134644, 0.001243698, 
    0.001017661, 0.000787762, 0.0007626964, 0.0009532245, 0.001192564, 
    0.001437104, 0.001500984, 0.001424706, 0.001451407, 0.001141019, 
    0.0008929055,
  0.001053154, 0.001432811, 0.00145829, 0.001221191, 0.001396301, 
    0.001085611, 0.0008917302, 0.0007369169, 0.0005643019, 0.0005046653, 
    0.0006026071, 0.0006974658, 0.0006238902, 0.0007635392, 0.000749012, 
    0.0009261251, 0.001070464, 0.001359793, 0.001295594, 0.0009553077, 
    0.0006953522, 0.0006147819, 0.0005600094, 0.0004685203, 0.0003308895, 
    0.0002793116, 0.0002964935, 0.0002994022, 0.0003587685, 0.0004064203, 
    0.0003976147, 0.0004222671, 0.0004084071, 0.0003095429, 0.0003369611, 
    0.0004662474, 0.0008742297, 0.0009697396, 0.0007554812, 0.001055619, 
    0.001005439, 0.0009113434, 0.0008420912, 0.0007982058, 0.0007907194, 
    0.0008076634, 0.0008144658, 0.0008157692, 0.0008265772, 0.0008380529, 
    0.000875643, 0.0009592487, 0.001012352, 0.001041217, 0.001086994, 
    0.001110486, 0.001184617, 0.001292907, 0.001333677, 0.001280255, 
    0.00121833, 0.001194981, 0.001107942, 0.0008606869, 0.0007308128, 
    0.0006948274, 0.0005903207, 0.0004689337, 0.0005591197, 0.0006036563, 
    0.0007578973, 0.0005653822, 0.0005599142, 0.0006485265, 0.0009055897, 
    0.0007955194, 0.0008104607, 0.000952224, 0.001282672, 0.001353323, 
    0.00127377, 0.001112551, 0.001051373, 0.0008806656, 0.000759962, 
    0.0007248987, 0.0006177863, 0.0004251273, 0.000530174, 0.0008255588, 
    0.001097038, 0.001266585, 0.001312918, 0.001245526, 0.0008782027, 
    0.0007639057,
  0.0007904014, 0.0007752385, 0.0008290899, 0.000854155, 0.0008250682, 
    0.0007524611, 0.0006459041, 0.0005691014, 0.0005958837, 0.0005529206, 
    0.0005574825, 0.0004691724, 0.0003659211, 0.0004305963, 0.0006856564, 
    0.0008555218, 0.0008541548, 0.0009467885, 0.0009473446, 0.0009471378, 
    0.0009753826, 0.0007206881, 0.0004721125, 0.0003240865, 0.0002515755, 
    0.0002205016, 0.0002075476, 0.0002130471, 0.0002488098, 0.0002708556, 
    0.0002871952, 0.0003378514, 0.0003377877, 0.0002798837, 0.0002918205, 
    0.0002724768, 0.0002952538, 0.0006907743, 0.0008079971, 0.000712232, 
    0.0006484312, 0.0006507519, 0.0006681404, 0.0006650102, 0.0006574441, 
    0.0006711613, 0.0006838446, 0.0006998824, 0.0007514441, 0.0007797205, 
    0.0007779882, 0.0008129082, 0.000881223, 0.0009356141, 0.0009995899, 
    0.001043172, 0.001069239, 0.00111349, 0.001159584, 0.001168882, 
    0.001172379, 0.001144881, 0.001048814, 0.0008735303, 0.0008328084, 
    0.0007129631, 0.0006166424, 0.0005787334, 0.0006304386, 0.0006875, 
    0.0007053021, 0.0004949691, 0.0005385999, 0.0007566574, 0.0007139167, 
    0.0007253136, 0.0007044754, 0.0007638417, 0.0008084895, 0.0008086483, 
    0.0008992795, 0.0008050082, 0.0006169127, 0.0005189856, 0.0004951432, 
    0.0005164896, 0.0004191031, 0.0002345508, 0.0002301643, 0.0004533716, 
    0.000657951, 0.0008585406, 0.0009944709, 0.001042138, 0.001024972, 
    0.0008199965,
  0.0007327516, 0.0007036333, 0.0007527322, 0.0007483766, 0.0007336421, 
    0.0007011057, 0.0005900345, 0.0005094809, 0.000456234, 0.0004603507, 
    0.0005488994, 0.0005647307, 0.0005078756, 0.0005228641, 0.0005595647, 
    0.0005439086, 0.0005339744, 0.0005781455, 0.0005300802, 0.0005187632, 
    0.0005529206, 0.0005565287, 0.0004796147, 0.0003506144, 0.0002803765, 
    0.0002165438, 0.000202048, 0.0002004427, 0.0002345524, 0.0002326292, 
    0.0002523066, 0.0002508284, 0.0002492866, 0.0002529742, 0.0002424043, 
    0.0002267481, 0.0002047341, 0.0002378744, 0.0004341407, 0.0004840177, 
    0.0005402369, 0.0005559726, 0.0005939128, 0.0005830091, 0.000576254, 
    0.0006031962, 0.0006484163, 0.0007100075, 0.0007669893, 0.0007861739, 
    0.0007831855, 0.0008174544, 0.000874023, 0.0009305123, 0.001018409, 
    0.001083052, 0.001095879, 0.001096626, 0.001094242, 0.001085404, 
    0.001078649, 0.001019998, 0.0008672997, 0.0007489643, 0.0006244308, 
    0.0006217125, 0.0006379092, 0.0007110559, 0.0007391894, 0.0005574984, 
    0.0005639676, 0.0005599464, 0.0005317336, 0.0005445606, 0.0006225868, 
    0.0006836378, 0.0006781701, 0.0006139082, 0.0005593261, 0.0005952324, 
    0.0007906882, 0.0005821032, 0.0004651991, 0.0004636892, 0.0004546768, 
    0.0003625513, 0.0002135392, -2.856692e-005, -0.0001875451, -7.26115e-005, 
    0.0002765288, 0.0006035119, 0.0007698806, 0.0008427096, 0.0009092758, 
    0.0009084176,
  0.0007283972, 0.0008136225, 0.0008055177, 0.0007290174, 0.0006056111, 
    0.0005810382, 0.0005498691, 0.0004833024, 0.0004270677, 0.0004145745, 
    0.0004268135, 0.0004073106, 0.0003981076, 0.000410267, 0.0004118405, 
    0.000398791, 0.0003794155, 0.0003647127, 0.0003815928, 0.0003989975, 
    0.0004075487, 0.000431645, 0.0004040678, 0.0003169497, 0.0002780401, 
    0.0002813302, 0.0002904219, 0.0002623681, 0.0002331219, 0.0002040666, 
    0.0001889032, 0.0001798273, 0.0001894435, 0.0001859944, 0.0001724522, 
    0.0001499614, 0.0001494528, 0.0002159239, 0.0005202892, 0.0005027098, 
    0.000571708, 0.0005923393, 0.0005176349, 0.0005497895, 0.000551363, 
    0.0006000164, 0.00065409, 0.000708672, 0.0007479799, 0.0007737924, 
    0.0007885904, 0.0008248771, 0.0008878987, 0.0009568497, 0.001010939, 
    0.001040757, 0.001051661, 0.001079253, 0.001083656, 0.001057399, 
    0.0009539085, 0.0008446339, 0.0007185421, 0.0005136612, 0.0004442973, 
    0.0004658344, 0.00049907, 0.0005621874, 0.0005598669, 0.0005361842, 
    0.0005062065, 0.0004997053, 0.0005209564, 0.0006242236, 0.000751619, 
    0.00102038, 0.0006913946, 0.0005501547, 0.0004420399, 0.0004461884, 
    0.0005320355, 0.00049214, 0.0004283073, 0.0003968049, 0.0003704678, 
    0.0003432082, 0.0002560737, 5.750265e-005, -0.0001641954, -0.0001936001, 
    5.551474e-005, 0.0004023979, 0.000607104, 0.0007156646, 0.0007687691, 
    0.0007595504,
  0.0006543272, 0.0007555918, 0.0007803403, 0.0007558784, 0.000683272, 
    0.0006774548, 0.0006401669, 0.0005294601, 0.0004687589, 0.0004402759, 
    0.0004484934, 0.000405308, 0.0003805282, 0.00040437, 0.0004244609, 
    0.0003867109, 0.0003629485, 0.0003653805, 0.0004076761, 0.0004168471, 
    0.0004098216, 0.0004067381, 0.0003956595, 0.0003626625, 0.0003369611, 
    0.0003077629, 0.0002802652, 0.0002304993, 0.0002067687, 0.0001953245, 
    0.0001733105, 0.000160563, 0.0001717529, 0.0001720708, 0.000155747, 
    0.0001388193, 0.0001513283, 0.0002015234, 0.0005621875, 0.0004322969, 
    0.0004856072, 0.0005488518, 0.000371786, 0.0003988863, 0.0005402847, 
    0.0006411993, 0.0007118825, 0.0007744434, 0.0008434101, 0.0008895362, 
    0.0009075133, 0.0009174629, 0.0009487276, 0.001029711, 0.001070798, 
    0.001080764, 0.001038627, 0.001000703, 0.0009998921, 0.0009738728, 
    0.0008603695, 0.0006719555, 0.0005192243, 0.0004695538, 0.0005028213, 
    0.000560423, 0.0005376779, 0.0004546922, 0.0003820857, 0.0004001736, 
    0.0004968761, 0.0006457129, 0.001167786, 0.001215502, 0.001219301, 
    0.001246147, 0.0007343888, 0.0006188989, 0.0005655726, 0.0005736945, 
    0.0006793784, 0.0005001668, 0.0004425331, 0.0004248265, 0.0004141612, 
    0.0003828174, 0.0003432403, 0.0002827132, 0.0002109171, 0.0002170997, 
    0.000332335, 0.0004941896, 0.0006307559, 0.0006960351, 0.000677343, 
    0.0006598281,
  0.0006368277, 0.0007175249, 0.000725202, 0.0006562674, 0.0006449982, 
    0.0006240015, 0.0006339513, 0.0005541926, 0.0004735909, 0.0004347448, 
    0.0004161003, 0.0003855985, 0.0003655235, 0.0003744243, 0.0003895878, 
    0.0004032095, 0.0003937841, 0.0003721197, 0.0003567974, 0.0003399969, 
    0.0003475308, 0.0003487072, 0.0003323201, 0.0003116092, 0.0002877515, 
    0.0002575996, 0.0002386691, 0.0002263509, 0.0002209943, 0.0002144139, 
    0.0001930198, 0.0001696865, 0.0001571616, 0.0001484356, 0.0001365623, 
    0.0001139443, 9.599935e-005, 9.646025e-005, 0.0001136582, 0.00014265, 
    0.0001652203, 0.0001801929, 0.0001862487, 0.0002023658, 0.0002573452, 
    0.0003650788, 0.0005072077, 0.0007156653, 0.0009669904, 0.00110602, 
    0.001168613, 0.001184667, 0.0009598059, 0.0008689526, 0.0008278334, 
    0.0008330945, 0.0008328561, 0.000750411, 0.0006414537, 0.0005560998, 
    0.0004971788, 0.0004587135, 0.0004356981, 0.0004126984, 0.0004116334, 
    0.0004312155, 0.0004378279, 0.0004137954, 0.0003885548, 0.0004215044, 
    0.0005222759, 0.001105638, 0.001228202, 0.001347681, 0.001438026, 
    0.001420081, 0.0007864436, 0.0007321159, 0.001320501, 0.001245288, 
    0.0009923422, 0.000684337, 0.0005423666, 0.0005514268, 0.0003795903, 
    0.000393705, 0.0004428199, 0.0004557893, 0.0004377491, 0.0004492239, 
    0.0004632277, 0.0004491764, 0.0003968515, 0.0003737886, 0.0004966855, 
    0.0005842648,
  0.0005169357, 0.0005665747, 0.0004880712, 0.0006480021, 0.0006118896, 
    0.000604324, 0.0006377818, 0.0006001119, 0.000576842, 0.0005397123, 
    0.000511102, 0.000466645, 0.0004390039, 0.0004178326, 0.0003991246, 
    0.0003872673, 0.0003685276, 0.0003539047, 0.000353857, 0.0003699741, 
    0.0003840408, 0.0003694337, 0.000328537, 0.0002798519, 0.0002450269, 
    0.0002200565, 0.000210329, 0.000199934, 0.0001885375, 0.000176092, 
    0.0001662534, 0.0001637102, 0.0001580676, 0.0001476249, 0.000129823, 
    0.0001163921, 0.0001166623, 0.0001021505, 0.0001057268, 0.0001058381, 
    0.0001054089, 0.0001386763, 0.0001621367, 0.0001840871, 0.0002035102, 
    0.0002201836, 0.0002422294, 0.0003067137, 0.0004535002, 0.0006738146, 
    0.0009063204, 0.001639378, 0.0009083705, 0.0006798387, 0.0005084156, 
    0.0004499714, 0.0004574259, 0.0004532615, 0.0004086454, 0.0003631552, 
    0.0003411412, 0.0003485004, 0.0003633936, 0.0003407915, 0.000300038, 
    0.0002814414, 0.0002945702, 0.0003287595, 0.0003522041, 0.0003295385, 
    0.0002974471, 0.0003007214, 0.0003509325, 0.0004410387, 0.0007195436, 
    0.0007139964, 0.0006882313, 0.0004224262, 0.0004630528, 0.000600668, 
    0.001148824, 0.001065489, 0.0005116423, 0.0002821407, 0.0001783493, 
    0.0001872343, 0.0002930124, 0.0004146856, 0.0005575302, 0.0006265133, 
    0.0006472557, 0.0008584461, 0.0005969487, 0.0004609078, 0.0004099496, 
    0.0004238412,
  0.0004943819, 0.0004502265, 0.0004389894, 0.0004194388, 0.000444409, 
    0.000635064, 0.0005881273, 0.0005379004, 0.0005157434, 0.000515187, 
    0.000544481, 0.0005413336, 0.0005903048, 0.0007326088, 0.00054758, 
    0.0004984976, 0.0004292607, 0.0003791295, 0.0003595157, 0.000351775, 
    0.0003371043, 0.0003209394, 0.0002923768, 0.0002612075, 0.0002313257, 
    0.0002064507, 0.0001849612, 0.0001624387, 0.0001501839, 0.0001473865, 
    0.0001485309, 0.0001426182, 0.000130125, 0.0001156768, 0.0001246732, 
    0.0001313012, 0.0001360378, 0.0001547775, 0.0001447957, 0.0001405996, 
    0.0001368802, 0.0001433652, 0.0001648228, 0.0001832924, 0.0002001565, 
    0.0001858673, 0.0001776816, 0.0001986942, 0.0002790412, 0.0005214176, 
    0.0009177169, 0.001183252, 0.001113459, 0.0005313518, 0.0004034482, 
    0.0003345133, 0.0003156623, 0.0003258667, 0.0003221633, 0.0003136756, 
    0.0003056171, 0.0002850494, 0.0002700767, 0.0002396546, 0.0002241255, 
    0.0002415459, 0.0002925835, 0.0003645858, 0.0004235707, 0.0009235027, 
    0.0004281642, 0.0003932119, 0.0003648243, 0.0005816262, 0.0003275675, 
    0.0003895244, 0.0003144543, 0.0003665567, 0.0004774055, 0.0009077034, 
    0.001102809, 0.001059735, 0.0003854873, 0.0001815439, 7.775237e-005, 
    5.673978e-005, 0.0001032949, 0.0002087077, 0.0003604375, 0.0005248985, 
    0.001112505, 0.001207618, 0.001076265, 0.0009035072, 0.0007546546, 
    0.0006121446,
  0.0007344687, 0.0006162606, 0.0005081145, 0.0004478581, 0.0003805764, 
    0.0003962326, 0.0005069538, 0.000624923, 0.0006934446, 0.0007162215, 
    0.0007097526, 0.0007379495, 0.0008922699, 0.001084785, 0.001106036, 
    0.0006594936, 0.0007638892, 0.0007064464, 0.0006247004, 0.0004277987, 
    0.000373598, 0.0003243566, 0.0002864957, 0.0002537688, 0.000227066, 
    0.0002062759, 0.0001930993, 0.0001818777, 0.0001770935, 0.000180177, 
    0.0001761239, 0.0001778564, 0.0001755358, 0.0001721184, 0.0001719913, 
    0.0002270184, 0.0002164961, 0.0002094548, 0.0001693687, 0.0001555881, 
    0.0001760126, 0.0001755358, 0.0001864872, 0.0002004744, 0.000209121, 
    0.0002086124, 0.0002020162, 0.0002010148, 0.0002180061, 0.0002535782, 
    0.0003017069, 0.000342254, 0.0003603738, 0.0003530941, 0.0003450355, 
    0.0003342272, 0.0003296973, 0.0003326219, 0.0003381532, 0.0003438911, 
    0.00034707, 0.0003385982, 0.0003147405, 0.0002453447, 0.0002318661, 
    0.0002294502, 0.0002428016, 0.0002738278, 0.0003111006, 0.0005640945, 
    0.0003395996, 0.0003113072, 0.0004335047, 0.0002325496, 0.0002150815, 
    0.0002158921, 0.0002490164, 0.0004038137, 0.0005285701, 0.0006298982, 
    0.0006367168, 0.0003577353, 0.000238065, 0.0001397094, 7.234825e-005, 
    3.971666e-005, 3.858816e-005, 6.524338e-005, 0.0001194756, 0.0001984717, 
    0.0003068885, 0.0005338472, 0.0007477241, 0.001047337, 0.001134233, 
    0.0008746905,
  0.0008941772, 0.0008084259, 0.000679235, 0.0006316146, 0.0005926571, 
    0.0007553226, 0.001054983, 0.001211735, 0.001219412, 0.0011795, 
    0.001113888, 0.001040487, 0.0009708682, 0.0008842747, 0.000791514, 
    0.0007099272, 0.0006535015, 0.0005922916, 0.0005297306, 0.0004748784, 
    0.0004383844, 0.0004018905, 0.0003725649, 0.0003428739, 0.0003166795, 
    0.0002804876, 0.0002632897, 0.0002314847, 0.0002124907, 0.0001986783, 
    0.000187107, 0.0002154312, 0.0002095184, 0.0002120297, 0.0002162577, 
    0.0002184194, 0.0002186737, 0.0002159557, 0.0002105992, 0.0002068163, 
    0.000202636, 0.0002030016, 0.0002075793, 0.0002132854, 0.00021621, 
    0.0002132377, 0.00020626, 0.0001992664, 0.0001965166, 0.0002004903, 
    0.0002133649, 0.0002325655, 0.0002524655, 0.0002671839, 0.0002739074, 
    0.0002716821, 0.0002639096, 0.0002549451, 0.0002506536, 0.0002538325, 
    0.0002632898, 0.0002744159, 0.000285272, 0.0002883237, 0.000283142, 
    0.0002382717, 0.0002262872, 0.0002173704, 0.0002100111, 0.0002058786, 
    0.0002004426, 0.0001910807, 0.0001833718, 0.0001747888, 0.000165856, 
    0.0001887442, 0.0001866461, 0.0002194207, 0.0001593551, 0.0001538715, 
    0.00014354, 0.0001301091, 0.000117314, 0.0001017214, 8.705072e-005, 
    7.416024e-005, 6.816798e-005, 7.576559e-005, 9.85584e-005, 0.0001393121, 
    0.0001927496, 0.0002646884, 0.0003836435, 0.0004989269, 0.0006287536, 
    0.0007729013,
  0.0004515452, 0.0004795989, 0.0005053162, 0.0005069375, 0.0004804414, 
    0.0004904073, 0.0004974169, 0.0005723916, 0.0005712154, 0.0005702458, 
    0.0005672894, 0.000561027, 0.0005496147, 0.0005337995, 0.0005114836, 
    0.0004834615, 0.0004526895, 0.0004213454, 0.0003920834, 0.0003652852, 
    0.0003444633, 0.0003259461, 0.0003124834, 0.000304266, 0.0003012937, 
    0.0002543888, 0.0002486667, 0.0002814889, 0.0002668501, 0.0002559464, 
    0.0002453607, 0.0002321364, 0.0002216301, 0.0002139689, 0.000207468, 
    0.0001999816, 0.00019329, 0.0001855494, 0.0001775226, 0.000170974, 
    0.0001658083, 0.0001621844, 0.0001611671, 0.0001627248, 0.0001671594, 
    0.0001727542, 0.000178524, 0.0001854858, 0.0001927178, 0.0002000293, 
    0.0002073408, 0.0002135715, 0.0002165915, 0.0002155424, 0.0002118231, 
    0.0002065143, 0.0002006492, 0.0001966915, 0.0001960398, 0.0002000135, 
    0.0002086601, 0.0002200088, 0.0002300065, 0.0002384942, 0.0002428493, 
    0.0002389869, 0.0002327722, 0.0002237918, 0.0002120616, 0.0001996638, 
    0.0001916847, 0.0001401545, 0.0001327635, 0.0001181405, 0.0001085561, 
    9.952794e-005, 8.957794e-005, 8.026375e-005, 7.309527e-005, 
    6.812029e-005, 6.490956e-005, 6.409893e-005, 6.524335e-005, 
    6.757984e-005, 7.190317e-005, 7.749803e-005, 8.655793e-005, 0.0001012605, 
    0.0001210333, 0.0001476885, 0.0001810512, 0.0002188644, 0.0002855262, 
    0.0003287913, 0.00037363, 0.0004153691,
  0.0003245157, 0.0003395042, 0.0003529192, 0.0003629646, 0.0003691317, 
    0.0003781916, 0.000387633, 0.000391384, 0.0003926556, 0.0003954531, 
    0.0003976625, 0.000398187, 0.0003962002, 0.0003920358, 0.000384613, 
    0.0003744563, 0.0003617884, 0.0003468475, 0.0003308098, 0.0003144544, 
    0.0002981623, 0.0002824586, 0.0002675813, 0.0002548497, 0.0002441845, 
    0.0002359193, 0.0002308489, 0.000225556, 0.0002181809, 0.0002140007, 
    0.0002107582, 0.000207627, 0.0002053699, 0.0002037646, 0.0002025407, 
    0.0002009035, 0.0001994571, 0.0001982174, 0.0001972955, 0.0001962941, 
    0.0001955788, 0.000195404, 0.0001955153, 0.000194959, 0.0001947047, 
    0.0001945616, 0.0001940053, 0.0001933854, 0.0001925589, 0.0001910012, 
    0.0001890303, 0.000186662, 0.0001841983, 0.0001816393, 0.0001793028, 
    0.0001776816, 0.0001769981, 0.00017792, 0.0001800499, 0.0001831652, 
    0.0001871706, 0.0001924635, 0.000197375, 0.0002019367, 0.000205513, 
    0.000207627, 0.0002075475, 0.0002063236, 0.0002035103, 0.0001998545, 
    0.0001953404, 0.0001870117, 0.0001811307, 0.0001760603, 0.0001708628, 
    0.0001663328, 0.0001606426, 0.0001536489, 0.0001475295, 0.0001431426, 
    0.0001394392, 0.0001358788, 0.0001342576, 0.0001361173, 0.0001392167, 
    0.0001452248, 0.0001546822, 0.0001666825, 0.000179732, 0.0001954358, 
    0.0002124589, 0.0002321841, 0.0002521635, 0.0002717138, 0.0002904217, 
    0.0003078264,
  0.0002526562, 0.0002569637, 0.000261589, 0.0002650381, 0.0002679945, 
    0.0002707284, 0.0002735258, 0.0002752424, 0.0002770226, 0.0002782942, 
    0.0002785485, 0.000278326, 0.0002772929, 0.00027591, 0.0002740504, 
    0.0002718251, 0.0002689164, 0.0002654196, 0.0002614459, 0.00025752, 
    0.0002537212, 0.0002496045, 0.0002453448, 0.0002411645, 0.0002370478, 
    0.0002332172, 0.0002294661, 0.0002263508, 0.0002234421, 0.0002209784, 
    0.0002190074, 0.0002172432, 0.000215463, 0.0002142391, 0.0002126179, 
    0.0002111397, 0.0002099316, 0.000208819, 0.0002077382, 0.0002065779, 
    0.0002054653, 0.0002043527, 0.0002033036, 0.0002020003, 0.0002005857, 
    0.0001993141, 0.0001978677, 0.0001964531, 0.0001947205, 0.0001928927, 
    0.0001915734, 0.0001899999, 0.0001885217, 0.0001875521, 0.0001865984, 
    0.0001857878, 0.000185613, 0.0001858514, 0.0001865349, 0.0001873614, 
    0.0001882991, 0.000189221, 0.0001907946, 0.0001924, 0.0001937828, 
    0.0001947524, 0.0001959127, 0.0001971842, 0.0001986624, 0.0001994254, 
    0.0002004903, 0.0002009353, 0.0002017142, 0.0002023341, 0.0002030017, 
    0.000203701, 0.0002038123, 0.0002036851, 0.000204003, 0.0002043209, 
    0.0002045752, 0.0002049408, 0.0002057037, 0.0002069912, 0.0002089621, 
    0.0002110761, 0.000213349, 0.0002162418, 0.0002192777, 0.0002221705, 
    0.0002260965, 0.0002299906, 0.0002344729, 0.0002388598, 0.0002434216, 
    0.0002472998 ;
}
