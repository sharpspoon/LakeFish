netcdf CGMR_SRA1B_1_tas-change_2070-2099
dimensions:
	time = 12 ;
	latitude = 160 ;
	longitude = 320 ;
	bounds = 2 ;
 latitude = 
    -89.14201, -88.02072, -86.89944, -85.77816, -84.65688, -83.53559, 
    -82.41431, -81.29302, -80.17174, -79.05046, -77.92918, -76.80789, 
    -75.68661, -74.56532, -73.44405, -72.32276, -71.20148, -70.08019, 
    -68.95891, -67.83763, -66.71635, -65.59506, -64.47378, -63.35249, 
    -62.23121, -61.10993, -59.98865, -58.86736, -57.74608, -56.6248, 
    -55.50351, -54.38223, -53.26095, -52.13966, -51.01838, -49.8971, 
    -48.77582, -47.65453, -46.53325, -45.41197, -44.29068, -43.1694, 
    -42.04812, -40.92683, -39.80555, -38.68427, -37.56298, -36.4417, 
    -35.32042, -34.19913, -33.07785, -31.95657, -30.83529, -29.714, 
    -28.59272, -27.47144, -26.35015, -25.22887, -24.10759, -22.98631, 
    -21.86502, -20.74374, -19.62246, -18.50117, -17.37989, -16.25861, 
    -15.13732, -14.01604, -12.89476, -11.77348, -10.65219, -9.530907, 
    -8.40963, -7.288345, -6.167061, -5.045776, -3.924492, -2.803207, 
    -1.681931, -0.5606461, 0.5606384, 1.681923, 2.803207, 3.924484, 5.045769, 
    6.167053, 7.288338, 8.409622, 9.530907, 10.65218, 11.77347, 12.89475, 
    14.01604, 15.13732, 16.2586, 17.37988, 18.50117, 19.62245, 20.74374, 
    21.86501, 22.9863, 24.10758, 25.22887, 26.35015, 27.47143, 28.59271, 
    29.714, 30.83528, 31.95657, 33.07785, 34.19913, 35.32041, 36.4417, 
    37.56298, 38.68427, 39.80555, 40.92683, 42.04812, 43.1694, 44.29067, 
    45.41196, 46.53324, 47.65453, 48.77581, 49.89709, 51.01838, 52.13966, 
    53.26095, 54.38223, 55.5035, 56.62479, 57.74607, 58.86736, 59.98864, 
    61.10992, 62.23121, 63.35249, 64.47378, 65.59505, 66.71633, 67.83762, 
    68.9589, 70.08019, 71.20147, 72.32275, 73.44404, 74.56532, 75.68661, 
    76.80788, 77.92918, 79.05045, 80.17173, 81.29302, 82.4143, 83.53559, 
    84.65687, 85.77814, 86.89944, 88.02071, 89.14201 ;
 longitude 
     0, 1.125, 2.25, 3.375, 4.5, 5.625, 6.750001, 7.875001, 9.000001, 
    10.125, 11.25, 12.375, 13.5, 14.625, 15.75, 16.875, 18, 19.125, 20.25, 
    21.375, 22.5, 23.625, 24.75, 25.875, 27, 28.125, 29.25, 30.375, 31.5, 
    32.625, 33.75, 34.875, 36, 37.125, 38.25, 39.375, 40.5, 41.625, 42.75, 
    43.875, 45, 46.125, 47.25, 48.375, 49.5, 50.625, 51.75, 52.875, 54.00001, 
    55.12501, 56.25001, 57.37501, 58.50001, 59.62501, 60.75001, 61.87501, 
    63.00001, 64.12501, 65.25001, 66.37501, 67.50001, 68.62501, 69.75001, 
    70.87501, 72.00001, 73.12501, 74.25001, 75.37501, 76.50001, 77.62501, 
    78.75001, 79.87501, 81.00001, 82.12501, 83.25001, 84.37501, 85.50001, 
    86.62501, 87.75001, 88.87501, 90.00001, 91.12501, 92.25001, 93.37501, 
    94.50001, 95.62501, 96.75001, 97.87501, 99.00001, 100.125, 101.25, 
    102.375, 103.5, 104.625, 105.75, 106.875, 108, 109.125, 110.25, 111.375, 
    112.5, 113.625, 114.75, 115.875, 117, 118.125, 119.25, 120.375, 121.5, 
    122.625, 123.75, 124.875, 126, 127.125, 128.25, 129.375, 130.5, 131.625, 
    132.75, 133.875, 135, 136.125, 137.25, 138.375, 139.5, 140.625, 141.75, 
    142.875, 144, 145.125, 146.25, 147.375, 148.5, 149.625, 150.75, 151.875, 
    153, 154.125, 155.25, 156.375, 157.5, 158.625, 159.75, 160.875, 162, 
    163.125, 164.25, 165.375, 166.5, 167.625, 168.75, 169.875, 171, 172.125, 
    173.25, 174.375, 175.5, 176.625, 177.75, 178.875, 180, 181.125, 182.25, 
    183.375, 184.5, 185.625, 186.75, 187.875, 189, 190.125, 191.25, 192.375, 
    193.5, 194.625, 195.75, 196.875, 198, 199.125, 200.25, 201.375, 202.5, 
    203.625, 204.75, 205.875, 207, 208.125, 209.25, 210.375, 211.5, 212.625, 
    213.75, 214.875, 216, 217.125, 218.25, 219.375, 220.5, 221.625, 222.75, 
    223.875, 225, 226.125, 227.25, 228.375, 229.5, 230.625, 231.75, 232.875, 
    234, 235.125, 236.25, 237.375, 238.5, 239.625, 240.75, 241.875, 243, 
    244.125, 245.25, 246.375, 247.5, 248.625, 249.75, 250.875, 252, 253.125, 
    254.25, 255.375, 256.5, 257.625, 258.75, 259.875, 261, 262.125, 263.25, 
    264.375, 265.5, 266.625, 267.75, 268.875, 270, 271.125, 272.25, 273.375, 
    274.5, 275.625, 276.75, 277.875, 279, 280.125, 281.25, 282.375, 283.5, 
    284.625, 285.75, 286.875, 288, 289.125, 290.25, 291.375, 292.5, 293.625, 
    294.75, 295.875, 297, 298.125, 299.25, 300.375, 301.5, 302.625, 303.75, 
    304.875, 306, 307.125, 308.25, 309.375, 310.5, 311.625, 312.75, 313.875, 
    315, 316.125, 317.25, 318.375, 319.5, 320.625, 321.75, 322.875, 324, 
    325.125, 326.25, 327.375, 328.5, 329.625, 330.75, 331.875, 333, 334.125, 
    335.25, 336.375, 337.5, 338.625, 339.75, 340.875, 342, 343.125, 344.25, 
    345.375, 346.5, 347.625, 348.75, 349.875, 351, 352.125, 353.25, 354.375, 
    355.5, 356.625, 357.75, 358.875 ;
