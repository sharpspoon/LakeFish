netcdf CGMR_SRA1B_1_tas-change_2070-2099
dimensions:
	time = 12 ;
	latitude = 48 ;
	longitude = 96 ;
	bounds = 2 ;
data: latitude 
    -87.16, -83.45, -79.74, -76.03, -72.32, -68.61, -64.91, -61.2, 
    -57.49, -53.78, -50.07, -46.36, -42.65, -38.94, -35.23, -31.53, -27.82, 
    -24.11, -20.4, -16.69, -12.98, -9.272, -5.563, -1.854, 1.854, 5.563, 
    9.272, 12.98, 16.69, 20.4, 24.11, 27.82, 31.53, 35.23, 38.94, 42.65, 
    46.36, 50.07, 53.78, 57.49, 61.2, 64.91, 68.61, 72.32, 76.03, 79.74, 
    83.45, 87.16 ;
 longitude 
    0, 3.75, 7.5, 11.25, 15, 18.75, 22.5, 26.25, 30, 33.75, 37.5, 
    41.25, 45, 48.75, 52.5, 56.25, 60, 63.75, 67.5, 71.25, 75, 78.75, 82.5, 
    86.25, 90, 93.75, 97.5, 101.3, 105, 108.8, 112.5, 116.3, 120, 123.8, 
    127.5, 131.3, 135, 138.8, 142.5, 146.3, 150, 153.8, 157.5, 161.3, 165, 
    168.8, 172.5, 176.3, 180, 183.8, 187.5, 191.3, 195, 198.8, 202.5, 206.3, 
    210, 213.8, 217.5, 221.3, 225, 228.8, 232.5, 236.3, 240, 243.8, 247.5, 
    251.3, 255, 258.8, 262.5, 266.3, 270, 273.8, 277.5, 281.3, 285, 288.8, 
    292.5, 296.3, 300, 303.8, 307.5, 311.3, 315, 318.8, 322.5, 326.3, 330, 
    333.8, 337.5, 341.3, 345, 348.8, 352.5, 356.3 ;
